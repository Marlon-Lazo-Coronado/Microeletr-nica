magic
tech scmos
timestamp 1626400951
<< metal1 >>
rect 576 1803 578 1807
rect 582 1803 585 1807
rect 589 1803 592 1807
rect 1600 1803 1602 1807
rect 1606 1803 1609 1807
rect 1613 1803 1616 1807
rect 1094 1788 1102 1791
rect 2374 1768 2382 1771
rect 10 1758 17 1761
rect 102 1761 105 1768
rect 894 1761 897 1768
rect 102 1758 113 1761
rect 142 1758 153 1761
rect 270 1758 281 1761
rect 342 1758 353 1761
rect 382 1758 393 1761
rect 422 1758 433 1761
rect 470 1758 481 1761
rect 886 1758 897 1761
rect 2662 1758 2670 1761
rect 886 1756 890 1758
rect 214 1748 241 1751
rect 14 1738 25 1741
rect 174 1738 193 1741
rect 206 1738 214 1741
rect 246 1738 254 1741
rect 446 1738 449 1748
rect 662 1748 678 1751
rect 718 1751 722 1753
rect 718 1748 729 1751
rect 910 1748 921 1751
rect 910 1742 913 1748
rect 1298 1748 1305 1751
rect 1874 1748 1881 1751
rect 2014 1748 2033 1751
rect 2182 1748 2190 1751
rect 606 1738 634 1741
rect 1270 1738 1278 1741
rect 1630 1738 1646 1741
rect 2222 1738 2225 1748
rect 2278 1742 2281 1751
rect 2422 1748 2430 1751
rect 2438 1748 2449 1751
rect 2534 1748 2553 1751
rect 2234 1738 2241 1741
rect 2550 1742 2553 1748
rect 2674 1748 2681 1751
rect 230 1728 241 1731
rect 258 1728 265 1731
rect 69 1718 70 1722
rect 238 1718 241 1728
rect 414 1718 417 1731
rect 886 1731 890 1733
rect 886 1728 897 1731
rect 902 1728 913 1731
rect 1278 1728 1289 1731
rect 1838 1731 1841 1738
rect 1838 1728 1849 1731
rect 1854 1728 1865 1731
rect 2422 1731 2425 1738
rect 2414 1728 2425 1731
rect 437 1718 438 1722
rect 1080 1703 1082 1707
rect 1086 1703 1089 1707
rect 1093 1703 1096 1707
rect 2104 1703 2106 1707
rect 2110 1703 2113 1707
rect 2117 1703 2120 1707
rect 2642 1688 2644 1692
rect 270 1678 281 1681
rect 54 1668 70 1671
rect 238 1671 241 1678
rect 134 1668 153 1671
rect 190 1668 209 1671
rect 222 1668 241 1671
rect 418 1668 420 1672
rect 462 1671 465 1681
rect 662 1678 670 1681
rect 758 1678 770 1681
rect 766 1677 770 1678
rect 950 1678 958 1681
rect 966 1678 977 1681
rect 1046 1678 1062 1681
rect 1318 1678 1329 1681
rect 1390 1678 1398 1681
rect 1414 1678 1425 1681
rect 1430 1678 1442 1681
rect 1702 1678 1713 1681
rect 1838 1678 1849 1681
rect 1858 1678 1866 1681
rect 2106 1678 2134 1681
rect 2242 1678 2257 1681
rect 950 1677 954 1678
rect 1438 1677 1442 1678
rect 1862 1677 1866 1678
rect 774 1672 778 1674
rect 1446 1672 1450 1674
rect 462 1668 473 1671
rect 486 1668 494 1671
rect 522 1668 529 1671
rect 534 1668 542 1671
rect 586 1668 593 1671
rect 854 1668 866 1671
rect 974 1668 985 1671
rect 1526 1668 1537 1671
rect 46 1658 54 1661
rect 254 1661 257 1668
rect 254 1658 265 1661
rect 326 1661 329 1668
rect 974 1662 977 1668
rect 326 1658 337 1661
rect 346 1658 361 1661
rect 454 1658 465 1661
rect 494 1658 510 1661
rect 630 1658 641 1661
rect 694 1658 705 1661
rect 742 1658 753 1661
rect 818 1658 825 1661
rect 1030 1658 1041 1661
rect 1174 1658 1185 1661
rect 1326 1661 1329 1668
rect 1326 1658 1337 1661
rect 1374 1658 1385 1661
rect 1414 1661 1417 1668
rect 1534 1662 1537 1668
rect 1950 1668 1962 1671
rect 2070 1668 2086 1671
rect 2262 1668 2273 1671
rect 1406 1658 1417 1661
rect 1490 1658 1497 1661
rect 1702 1661 1705 1668
rect 1682 1658 1689 1661
rect 1694 1658 1705 1661
rect 1838 1661 1841 1668
rect 1830 1658 1841 1661
rect 2270 1662 2273 1668
rect 2154 1658 2161 1661
rect 2166 1658 2182 1661
rect 2286 1658 2294 1661
rect 2318 1658 2334 1661
rect 2422 1661 2425 1671
rect 2494 1668 2505 1671
rect 2494 1662 2497 1668
rect 2422 1658 2433 1661
rect 2466 1658 2473 1661
rect 2478 1658 2486 1661
rect 2582 1658 2593 1661
rect 318 1648 329 1651
rect 2118 1648 2129 1651
rect 2318 1648 2321 1658
rect 2370 1648 2374 1652
rect 274 1638 297 1641
rect 2027 1638 2030 1642
rect 2118 1641 2121 1648
rect 2206 1641 2210 1644
rect 2102 1638 2121 1641
rect 2198 1638 2210 1641
rect 45 1618 46 1622
rect 250 1618 251 1622
rect 362 1618 363 1622
rect 576 1603 578 1607
rect 582 1603 585 1607
rect 589 1603 592 1607
rect 1600 1603 1602 1607
rect 1606 1603 1609 1607
rect 1613 1603 1616 1607
rect 885 1588 886 1592
rect 914 1588 915 1592
rect 2338 1588 2339 1592
rect 2413 1588 2414 1592
rect 2437 1588 2438 1592
rect 2554 1588 2555 1592
rect 1917 1568 1918 1572
rect 86 1558 97 1561
rect 998 1561 1001 1568
rect 990 1558 1001 1561
rect 54 1548 65 1551
rect 126 1548 137 1551
rect 166 1548 177 1551
rect 222 1548 241 1551
rect 382 1548 393 1551
rect 462 1548 470 1551
rect 134 1542 137 1548
rect 14 1538 33 1541
rect 86 1538 94 1541
rect 278 1538 292 1541
rect 310 1538 329 1541
rect 342 1538 369 1541
rect 410 1538 417 1541
rect 598 1538 626 1541
rect 806 1541 809 1551
rect 842 1548 857 1551
rect 806 1538 825 1541
rect 878 1541 881 1551
rect 1014 1551 1017 1558
rect 942 1548 961 1551
rect 1014 1548 1025 1551
rect 1062 1548 1078 1551
rect 1390 1548 1401 1551
rect 1686 1542 1689 1551
rect 1710 1548 1729 1551
rect 1774 1551 1777 1561
rect 2246 1558 2257 1561
rect 1758 1548 1777 1551
rect 1870 1548 1889 1551
rect 1902 1548 1913 1551
rect 1930 1548 1945 1551
rect 1950 1548 1969 1551
rect 1990 1548 1998 1551
rect 1902 1542 1905 1548
rect 2226 1548 2233 1551
rect 2370 1548 2372 1552
rect 2438 1548 2457 1551
rect 2614 1548 2625 1551
rect 874 1538 881 1541
rect 1098 1538 1110 1541
rect 1742 1538 1750 1541
rect 1778 1538 1785 1541
rect 1862 1538 1870 1541
rect 2002 1538 2009 1541
rect 2582 1538 2601 1541
rect 278 1532 281 1538
rect 350 1528 353 1538
rect 390 1531 393 1538
rect 390 1528 401 1531
rect 478 1528 489 1531
rect 774 1528 777 1538
rect 782 1528 793 1531
rect 962 1528 969 1531
rect 974 1528 982 1531
rect 1010 1528 1022 1531
rect 1038 1528 1049 1531
rect 1830 1528 1838 1531
rect 2598 1528 2601 1538
rect 2606 1528 2614 1531
rect 2630 1528 2646 1531
rect 101 1518 102 1522
rect 1810 1518 1811 1522
rect 1080 1503 1082 1507
rect 1086 1503 1089 1507
rect 1093 1503 1096 1507
rect 2104 1503 2106 1507
rect 2110 1503 2113 1507
rect 2117 1503 2120 1507
rect 845 1488 846 1492
rect 390 1478 401 1481
rect 1052 1478 1054 1482
rect 1122 1478 1129 1481
rect 1470 1478 1482 1481
rect 390 1477 394 1478
rect 1478 1477 1482 1478
rect 1726 1478 1737 1481
rect 2198 1478 2209 1481
rect 2254 1478 2262 1481
rect 1494 1474 1498 1478
rect 22 1468 33 1471
rect 126 1468 145 1471
rect 22 1462 25 1468
rect 230 1462 233 1471
rect 406 1468 417 1471
rect 446 1468 457 1471
rect 510 1468 537 1471
rect 558 1468 569 1471
rect 618 1468 625 1471
rect 1006 1468 1017 1471
rect 1078 1468 1094 1471
rect 1110 1468 1126 1471
rect 1386 1468 1393 1471
rect 58 1458 73 1461
rect 78 1458 86 1461
rect 174 1458 193 1461
rect 598 1458 617 1461
rect 958 1461 961 1468
rect 958 1458 969 1461
rect 974 1458 993 1461
rect 1070 1458 1078 1461
rect 1142 1458 1161 1461
rect 1326 1458 1337 1461
rect 1374 1458 1385 1461
rect 1414 1458 1422 1461
rect 1454 1458 1465 1461
rect 1510 1458 1518 1461
rect 1734 1461 1737 1468
rect 1846 1468 1854 1471
rect 1910 1462 1913 1471
rect 1938 1468 1945 1471
rect 2086 1468 2113 1471
rect 2138 1468 2153 1471
rect 2258 1468 2273 1471
rect 2290 1468 2297 1471
rect 1674 1458 1681 1461
rect 1734 1458 1745 1461
rect 1750 1458 1769 1461
rect 1830 1458 1841 1461
rect 1946 1458 1953 1461
rect 1958 1458 1966 1461
rect 2166 1458 2177 1461
rect 2234 1458 2241 1461
rect 2334 1461 2337 1468
rect 2334 1458 2345 1461
rect 2422 1458 2430 1461
rect 2550 1461 2553 1471
rect 2590 1468 2601 1471
rect 2646 1471 2649 1478
rect 2662 1472 2665 1481
rect 2682 1478 2689 1482
rect 2686 1472 2689 1478
rect 2646 1468 2657 1471
rect 2666 1468 2673 1471
rect 2590 1462 2593 1468
rect 2550 1458 2561 1461
rect 2606 1458 2614 1461
rect 174 1456 178 1458
rect 106 1448 111 1452
rect 138 1448 145 1451
rect 1974 1451 1978 1454
rect 1966 1448 1978 1451
rect 2402 1448 2409 1451
rect 838 1442 842 1444
rect 1166 1441 1170 1444
rect 1026 1438 1049 1441
rect 1166 1438 1182 1441
rect 2509 1438 2510 1442
rect 18 1418 19 1422
rect 1138 1418 1139 1422
rect 576 1403 578 1407
rect 582 1403 585 1407
rect 589 1403 592 1407
rect 1600 1403 1602 1407
rect 1606 1403 1609 1407
rect 1613 1403 1616 1407
rect 562 1388 563 1392
rect 2554 1388 2555 1392
rect 770 1368 773 1372
rect 1522 1368 1525 1372
rect 1998 1368 2006 1371
rect 2346 1368 2353 1371
rect 2589 1368 2590 1372
rect 30 1358 41 1361
rect 150 1361 153 1368
rect 142 1358 153 1361
rect 198 1358 209 1361
rect 118 1348 126 1351
rect 158 1348 169 1351
rect 230 1348 241 1351
rect 350 1351 353 1361
rect 2262 1358 2270 1361
rect 2322 1358 2329 1361
rect 302 1348 329 1351
rect 334 1348 353 1351
rect 366 1348 385 1351
rect 166 1342 169 1348
rect 542 1348 554 1351
rect 574 1348 617 1351
rect 674 1348 681 1351
rect 794 1348 809 1351
rect 1106 1348 1113 1351
rect 1130 1348 1138 1351
rect 550 1346 554 1348
rect 1134 1346 1138 1348
rect 1926 1348 1942 1351
rect 2046 1348 2057 1351
rect 2210 1348 2217 1351
rect 2438 1351 2441 1361
rect 2450 1358 2454 1362
rect 2422 1348 2441 1351
rect 2486 1348 2494 1351
rect 2626 1348 2633 1351
rect 130 1338 137 1341
rect 1806 1338 1814 1341
rect 2202 1338 2209 1341
rect 2290 1338 2297 1341
rect 2338 1338 2345 1341
rect 2678 1338 2686 1341
rect 70 1332 73 1338
rect 70 1328 78 1332
rect 98 1328 105 1331
rect 390 1328 393 1338
rect 486 1331 490 1333
rect 486 1328 497 1331
rect 1018 1328 1030 1331
rect 1114 1328 1121 1331
rect 1182 1328 1185 1338
rect 2046 1328 2054 1331
rect 2606 1331 2609 1338
rect 2606 1328 2617 1331
rect 306 1318 307 1322
rect 2282 1318 2283 1322
rect 2306 1318 2307 1322
rect 1080 1303 1082 1307
rect 1086 1303 1089 1307
rect 1093 1303 1096 1307
rect 2104 1303 2106 1307
rect 2110 1303 2113 1307
rect 2117 1303 2120 1307
rect 36 1288 38 1292
rect 330 1288 331 1292
rect 566 1288 574 1291
rect 1086 1288 1102 1291
rect 1757 1288 1758 1292
rect 1909 1288 1910 1292
rect 86 1271 89 1281
rect 262 1278 273 1281
rect 262 1272 265 1278
rect 438 1272 441 1281
rect 614 1278 622 1281
rect 1262 1278 1273 1281
rect 1414 1278 1425 1281
rect 1522 1278 1529 1282
rect 1574 1278 1585 1281
rect 2114 1278 2129 1281
rect 2462 1278 2473 1281
rect 86 1268 105 1271
rect 182 1268 190 1271
rect 218 1268 225 1271
rect 606 1268 614 1271
rect 798 1268 817 1271
rect 934 1271 937 1278
rect 934 1268 953 1271
rect 110 1258 121 1261
rect 198 1258 217 1261
rect 254 1258 265 1261
rect 282 1258 297 1261
rect 414 1258 433 1261
rect 586 1258 593 1261
rect 830 1258 846 1261
rect 934 1258 937 1268
rect 1026 1268 1033 1271
rect 1054 1268 1073 1271
rect 1406 1268 1414 1271
rect 1502 1271 1505 1278
rect 1526 1272 1529 1278
rect 1582 1272 1585 1278
rect 1502 1268 1513 1271
rect 1198 1258 1217 1261
rect 1326 1258 1334 1261
rect 1454 1261 1457 1268
rect 1438 1258 1457 1261
rect 1546 1258 1561 1261
rect 1602 1258 1625 1261
rect 1878 1261 1881 1271
rect 2134 1268 2150 1271
rect 2158 1268 2174 1271
rect 2190 1268 2217 1271
rect 2226 1268 2241 1271
rect 2262 1268 2281 1271
rect 2390 1268 2401 1271
rect 2630 1271 2633 1281
rect 2630 1268 2649 1271
rect 2654 1268 2670 1271
rect 2686 1268 2694 1271
rect 1878 1258 1897 1261
rect 2102 1258 2118 1261
rect 2494 1258 2521 1261
rect 2598 1258 2609 1261
rect 2662 1258 2681 1261
rect 164 1248 166 1252
rect 366 1248 377 1251
rect 410 1248 414 1252
rect 1510 1251 1513 1258
rect 1502 1248 1513 1251
rect 1894 1248 1905 1251
rect 2422 1248 2430 1251
rect 2534 1248 2545 1251
rect 1902 1242 1906 1244
rect 706 1238 709 1242
rect 2374 1238 2382 1241
rect 2410 1228 2411 1232
rect 2341 1218 2342 1222
rect 576 1203 578 1207
rect 582 1203 585 1207
rect 589 1203 592 1207
rect 1600 1203 1602 1207
rect 1606 1203 1609 1207
rect 1613 1203 1616 1207
rect 186 1188 187 1192
rect 274 1188 275 1192
rect 2138 1188 2139 1192
rect 2237 1188 2238 1192
rect 2650 1188 2651 1192
rect 306 1168 307 1172
rect 454 1168 462 1171
rect 734 1168 745 1171
rect 1310 1168 1318 1171
rect 1675 1168 1678 1172
rect 1979 1168 1982 1172
rect 478 1158 489 1161
rect 742 1158 745 1168
rect 1098 1158 1105 1161
rect 1150 1158 1161 1161
rect 1190 1158 1201 1161
rect 1270 1158 1281 1161
rect 1338 1158 1342 1162
rect 14 1148 25 1151
rect 30 1148 49 1151
rect 94 1148 105 1151
rect 114 1148 140 1151
rect 322 1148 329 1151
rect 610 1148 617 1151
rect 878 1148 889 1151
rect 886 1142 889 1148
rect 1054 1148 1062 1151
rect 1502 1151 1505 1158
rect 1550 1151 1553 1161
rect 1502 1148 1537 1151
rect 1550 1148 1561 1151
rect 1582 1148 1590 1151
rect 70 1138 89 1141
rect 226 1138 233 1141
rect 470 1138 478 1141
rect 1014 1138 1033 1141
rect 1442 1138 1457 1141
rect 1558 1141 1561 1148
rect 2070 1151 2073 1161
rect 2434 1158 2441 1161
rect 2482 1158 2489 1161
rect 2054 1148 2073 1151
rect 2130 1148 2137 1151
rect 2166 1148 2177 1151
rect 2294 1148 2310 1151
rect 2470 1148 2478 1151
rect 2590 1148 2617 1151
rect 2634 1148 2649 1151
rect 1558 1138 1569 1141
rect 1694 1138 1705 1141
rect 1710 1138 1737 1141
rect 2086 1138 2094 1141
rect 2102 1138 2129 1141
rect 2378 1138 2385 1141
rect 2566 1138 2574 1141
rect 2686 1138 2702 1141
rect 70 1128 73 1138
rect 1470 1128 1473 1138
rect 1694 1136 1698 1138
rect 2194 1128 2201 1131
rect 2206 1128 2214 1131
rect 2330 1128 2337 1131
rect 1034 1118 1035 1122
rect 1146 1118 1147 1122
rect 1186 1118 1187 1122
rect 1778 1118 1785 1121
rect 2370 1118 2371 1122
rect 2493 1118 2494 1122
rect 2677 1118 2678 1122
rect 1080 1103 1082 1107
rect 1086 1103 1089 1107
rect 1093 1103 1096 1107
rect 2104 1103 2106 1107
rect 2110 1103 2113 1107
rect 2117 1103 2120 1107
rect 1510 1088 1521 1091
rect 2434 1088 2436 1092
rect 342 1078 353 1081
rect 454 1072 457 1081
rect 514 1078 521 1081
rect 1174 1078 1182 1081
rect 1198 1078 1209 1081
rect 1510 1081 1513 1088
rect 1502 1078 1513 1081
rect 1606 1078 1622 1081
rect 2186 1078 2187 1082
rect 46 1068 54 1071
rect 138 1068 145 1071
rect 190 1068 198 1071
rect 414 1068 441 1071
rect 462 1068 481 1071
rect 602 1068 625 1071
rect 790 1068 809 1071
rect 854 1068 873 1071
rect 950 1071 954 1072
rect 958 1071 961 1078
rect 950 1068 961 1071
rect 1066 1068 1068 1072
rect 1114 1068 1121 1071
rect 1134 1068 1158 1071
rect 1494 1068 1502 1071
rect 46 1058 65 1061
rect 70 1058 86 1061
rect 214 1061 217 1068
rect 206 1058 217 1061
rect 350 1061 353 1068
rect 350 1058 361 1061
rect 470 1058 478 1061
rect 494 1058 513 1061
rect 606 1058 614 1061
rect 774 1058 777 1068
rect 1542 1068 1550 1071
rect 1574 1068 1593 1071
rect 2398 1071 2401 1081
rect 2382 1068 2401 1071
rect 2494 1071 2497 1081
rect 2478 1068 2497 1071
rect 2670 1068 2681 1071
rect 886 1058 894 1061
rect 1022 1058 1041 1061
rect 1142 1058 1150 1061
rect 1174 1058 1185 1061
rect 1438 1058 1446 1061
rect 1854 1061 1857 1068
rect 1846 1058 1857 1061
rect 1974 1061 1977 1068
rect 1966 1058 1977 1061
rect 2046 1058 2065 1061
rect 2246 1058 2254 1061
rect 2370 1058 2377 1061
rect 2522 1058 2537 1061
rect 2542 1058 2550 1061
rect 162 1048 164 1052
rect 678 1051 682 1054
rect 670 1048 682 1051
rect 906 1048 913 1051
rect 918 1048 929 1051
rect 1638 1051 1641 1058
rect 1638 1048 1649 1051
rect 1834 1048 1838 1052
rect 1846 1048 1849 1058
rect 1954 1048 1958 1052
rect 1966 1048 1969 1058
rect 2046 1052 2049 1058
rect 2122 1048 2137 1051
rect 1884 1038 1886 1042
rect 2004 1038 2006 1042
rect 578 1018 585 1021
rect 981 1018 982 1022
rect 1042 1018 1043 1022
rect 2362 1018 2363 1022
rect 2578 1018 2580 1022
rect 576 1003 578 1007
rect 582 1003 585 1007
rect 589 1003 592 1007
rect 1600 1003 1602 1007
rect 1606 1003 1609 1007
rect 1613 1003 1616 1007
rect 242 988 243 992
rect 1450 988 1451 992
rect 2221 988 2222 992
rect 404 968 406 972
rect 710 968 721 971
rect 1298 968 1301 972
rect 1611 968 1614 972
rect 2642 968 2644 972
rect 10 958 17 961
rect 718 958 721 968
rect 1874 958 1878 962
rect 1886 958 1897 961
rect 822 952 826 954
rect 70 948 81 951
rect 334 948 345 951
rect 506 948 513 951
rect 518 948 537 951
rect 766 948 785 951
rect 854 951 858 954
rect 1222 953 1226 958
rect 854 948 862 951
rect 1014 948 1025 951
rect 1014 942 1017 948
rect 1434 948 1449 951
rect 1650 948 1657 951
rect 1942 948 1950 951
rect 2030 948 2049 951
rect 2134 951 2137 961
rect 2282 958 2289 961
rect 2102 948 2137 951
rect 2330 948 2337 951
rect 2442 948 2449 951
rect 2526 948 2534 951
rect 2670 948 2681 951
rect 14 938 25 941
rect 54 938 73 941
rect 78 938 89 941
rect 138 938 145 941
rect 278 938 294 941
rect 310 938 329 941
rect 550 938 569 941
rect 898 938 905 941
rect 994 938 1001 941
rect 1146 938 1154 941
rect 1254 938 1265 941
rect 1670 938 1697 941
rect 2350 938 2358 941
rect 2622 941 2625 948
rect 2550 938 2569 941
rect 2614 938 2625 941
rect 2670 942 2673 948
rect 78 928 81 938
rect 310 928 313 938
rect 1262 932 1265 938
rect 434 928 441 931
rect 1398 928 1409 931
rect 2130 928 2142 931
rect 2278 928 2294 931
rect 2694 928 2702 931
rect 204 918 206 922
rect 269 918 270 922
rect 566 918 574 921
rect 1126 918 1134 921
rect 1630 918 1646 921
rect 2178 918 2180 922
rect 2317 918 2318 922
rect 2405 918 2406 922
rect 2586 918 2588 922
rect 1080 903 1082 907
rect 1086 903 1089 907
rect 1093 903 1096 907
rect 2104 903 2106 907
rect 2110 903 2113 907
rect 2117 903 2120 907
rect 77 888 78 892
rect 140 888 142 892
rect 244 888 246 892
rect 2602 888 2604 892
rect 2658 888 2660 892
rect 54 881 58 882
rect 46 878 58 881
rect 1090 878 1105 881
rect 1322 878 1329 881
rect 1334 878 1345 881
rect 30 868 41 871
rect 78 868 97 871
rect 106 868 113 871
rect 182 868 201 871
rect 326 862 329 871
rect 550 868 558 871
rect 1018 868 1025 871
rect 1206 871 1210 874
rect 1974 872 1977 881
rect 2090 878 2097 881
rect 1198 868 1210 871
rect 1346 868 1353 871
rect 1362 868 1370 871
rect 1670 868 1681 871
rect 1910 868 1929 871
rect 2102 868 2129 871
rect 2182 868 2201 871
rect 2206 868 2214 871
rect 2454 868 2465 871
rect 2502 868 2521 871
rect 2630 868 2638 871
rect 22 858 30 861
rect 38 858 57 861
rect 766 861 769 868
rect 766 858 777 861
rect 986 858 993 861
rect 998 858 1014 861
rect 1038 858 1046 861
rect 1238 858 1246 861
rect 1302 861 1305 868
rect 1302 858 1313 861
rect 1418 858 1425 861
rect 1618 858 1633 861
rect 1694 858 1713 861
rect 1910 858 1913 868
rect 2010 858 2022 861
rect 2074 858 2081 861
rect 2086 858 2094 861
rect 2142 858 2161 861
rect 2214 858 2222 861
rect 2254 861 2257 868
rect 2246 858 2257 861
rect 2342 858 2350 861
rect 2390 861 2393 868
rect 2382 858 2393 861
rect 2422 858 2441 861
rect 2458 858 2473 861
rect 2478 858 2497 861
rect 2566 858 2574 861
rect 1134 856 1138 858
rect 18 848 22 852
rect 526 848 537 851
rect 594 848 609 851
rect 662 841 665 851
rect 1174 848 1185 851
rect 1574 848 1582 851
rect 1694 848 1697 858
rect 2158 848 2161 858
rect 2246 848 2249 858
rect 2278 848 2289 851
rect 662 838 673 841
rect 1862 841 1866 844
rect 1854 838 1866 841
rect 2298 838 2305 841
rect 2173 818 2174 822
rect 576 803 578 807
rect 582 803 585 807
rect 589 803 592 807
rect 1600 803 1602 807
rect 1606 803 1609 807
rect 1613 803 1616 807
rect 574 788 582 791
rect 773 788 774 792
rect 1426 788 1427 792
rect 2322 788 2323 792
rect 2621 788 2622 792
rect 85 778 86 782
rect 2230 768 2238 771
rect 2286 771 2289 781
rect 2270 768 2289 771
rect 206 758 214 761
rect 442 758 446 762
rect 1654 758 1665 761
rect 14 748 22 751
rect 22 738 33 741
rect 46 738 54 741
rect 94 738 105 741
rect 126 738 145 741
rect 198 738 209 741
rect 326 738 345 741
rect 418 738 425 741
rect 462 741 465 751
rect 514 748 529 751
rect 458 738 465 741
rect 486 738 505 741
rect 542 738 545 748
rect 694 742 697 751
rect 894 751 897 758
rect 886 748 897 751
rect 918 748 934 751
rect 966 748 977 751
rect 710 738 729 741
rect 918 738 921 748
rect 974 742 977 748
rect 1410 748 1425 751
rect 2334 751 2337 761
rect 2334 748 2353 751
rect 2358 748 2385 751
rect 1186 738 1194 741
rect 1398 738 1417 741
rect 1790 738 1798 741
rect 1838 738 1849 741
rect 1966 738 1977 741
rect 2242 738 2249 741
rect 2270 738 2273 748
rect 2390 742 2393 751
rect 2454 748 2462 751
rect 2542 751 2546 754
rect 2542 748 2561 751
rect 2570 748 2585 751
rect 2622 748 2649 751
rect 2406 741 2409 748
rect 2406 738 2417 741
rect 2446 738 2465 741
rect 22 728 25 738
rect 958 731 961 738
rect 1846 732 1849 738
rect 894 728 910 731
rect 950 728 961 731
rect 1882 728 1894 731
rect 2210 728 2217 731
rect 234 718 235 722
rect 378 718 380 722
rect 1650 718 1651 722
rect 2426 718 2427 722
rect 2482 718 2484 722
rect 1080 703 1082 707
rect 1086 703 1089 707
rect 1093 703 1096 707
rect 2104 703 2106 707
rect 2110 703 2113 707
rect 2117 703 2120 707
rect 314 688 315 692
rect 1962 688 1964 692
rect 2282 688 2283 692
rect 2594 688 2596 692
rect 30 668 46 671
rect 70 671 73 681
rect 1766 678 1774 682
rect 54 668 73 671
rect 194 668 201 671
rect 206 668 214 671
rect 294 668 305 671
rect 326 668 345 671
rect 414 671 418 672
rect 422 671 425 678
rect 1766 672 1769 678
rect 414 668 425 671
rect 610 668 625 671
rect 906 668 908 672
rect 986 668 993 671
rect 1014 668 1025 671
rect 1110 668 1121 671
rect 1334 668 1342 671
rect 1426 668 1433 671
rect 1478 668 1497 671
rect 1606 668 1614 671
rect 1626 668 1633 671
rect 1754 668 1761 671
rect 1846 668 1854 671
rect 2066 668 2073 671
rect 2078 668 2097 671
rect 2318 668 2326 671
rect 2478 671 2481 678
rect 2478 668 2492 671
rect 2630 668 2641 671
rect 294 662 297 668
rect 342 662 345 668
rect 42 658 49 661
rect 130 658 137 661
rect 210 658 217 661
rect 250 658 257 661
rect 430 658 449 661
rect 686 658 705 661
rect 1014 662 1017 668
rect 1118 662 1121 668
rect 1038 658 1046 661
rect 1082 658 1097 661
rect 1154 658 1162 661
rect 1282 658 1289 661
rect 1510 658 1513 668
rect 2630 662 2633 668
rect 1562 658 1577 661
rect 1698 658 1705 661
rect 1730 658 1737 661
rect 1786 658 1793 661
rect 1822 658 1849 661
rect 1886 658 1894 661
rect 2134 658 2142 661
rect 2230 658 2238 661
rect 2390 658 2409 661
rect 2522 658 2537 661
rect 2654 658 2662 661
rect 22 651 25 658
rect 430 656 434 658
rect 14 648 25 651
rect 326 648 345 651
rect 350 648 361 651
rect 454 651 457 658
rect 1158 656 1162 658
rect 454 648 465 651
rect 834 648 838 652
rect 1646 648 1657 651
rect 2038 648 2049 651
rect 2174 648 2182 651
rect 2250 648 2254 652
rect 2262 648 2270 651
rect 2334 648 2345 651
rect 2462 648 2473 651
rect 2550 648 2561 651
rect 358 642 361 648
rect 414 638 430 641
rect 2102 638 2110 641
rect 709 628 710 632
rect 1237 618 1238 622
rect 1810 618 1811 622
rect 576 603 578 607
rect 582 603 585 607
rect 589 603 592 607
rect 1600 603 1602 607
rect 1606 603 1609 607
rect 1613 603 1616 607
rect 85 588 86 592
rect 266 588 268 592
rect 717 588 718 592
rect 2293 588 2294 592
rect 850 568 853 572
rect 1234 568 1241 571
rect 1274 568 1281 571
rect 1458 568 1497 571
rect 36 558 38 562
rect 342 558 353 561
rect 70 548 81 551
rect 110 548 118 551
rect 158 548 169 551
rect 214 548 233 551
rect 166 542 169 548
rect 734 551 737 561
rect 2446 558 2454 561
rect 2618 558 2622 562
rect 822 552 826 554
rect 1222 552 1226 554
rect 722 548 737 551
rect 1070 548 1086 551
rect 1278 548 1297 551
rect 770 538 777 541
rect 1270 541 1273 548
rect 1342 542 1345 551
rect 2286 542 2289 551
rect 2478 548 2513 551
rect 2670 551 2673 561
rect 2670 548 2689 551
rect 1262 538 1273 541
rect 1310 538 1318 541
rect 1718 538 1726 541
rect 1790 538 1798 541
rect 1834 538 1842 541
rect 2038 538 2046 541
rect 2302 538 2313 541
rect 2498 538 2505 541
rect 2646 538 2657 541
rect 2662 538 2670 541
rect 1102 536 1106 538
rect 174 528 193 531
rect 398 528 417 531
rect 1950 531 1954 533
rect 2302 532 2305 538
rect 1942 528 1954 531
rect 1080 503 1082 507
rect 1086 503 1089 507
rect 1093 503 1096 507
rect 2104 503 2106 507
rect 2110 503 2113 507
rect 2117 503 2120 507
rect 36 488 38 492
rect 212 488 214 492
rect 402 488 403 492
rect 2685 488 2686 492
rect 126 478 145 481
rect 414 471 417 481
rect 670 478 686 481
rect 702 478 713 481
rect 734 478 745 481
rect 702 472 705 478
rect 410 468 417 471
rect 614 468 622 471
rect 930 468 937 471
rect 986 468 993 471
rect 1018 468 1025 471
rect 1046 468 1065 471
rect 1173 468 1174 472
rect 1270 471 1273 481
rect 1474 478 1490 481
rect 1486 474 1490 478
rect 1598 478 1625 481
rect 1598 477 1602 478
rect 1270 468 1289 471
rect 66 458 73 461
rect 110 458 121 461
rect 274 458 289 461
rect 294 458 305 461
rect 746 458 753 461
rect 850 458 857 461
rect 1006 458 1030 461
rect 1406 462 1409 471
rect 2022 468 2033 471
rect 2078 468 2094 471
rect 2702 471 2705 478
rect 2694 468 2705 471
rect 1238 458 1257 461
rect 1262 458 1270 461
rect 1542 458 1550 461
rect 1562 458 1569 461
rect 1638 458 1649 461
rect 1818 458 1833 461
rect 2022 462 2026 464
rect 2054 458 2062 461
rect 1582 452 1586 457
rect 246 448 257 451
rect 406 448 425 451
rect 1098 448 1105 451
rect 1126 441 1129 451
rect 2054 448 2057 458
rect 1126 438 1137 441
rect 338 418 340 422
rect 1078 418 1094 421
rect 576 403 578 407
rect 582 403 585 407
rect 589 403 592 407
rect 1600 403 1602 407
rect 1606 403 1609 407
rect 1613 403 1616 407
rect 197 388 198 392
rect 317 388 318 392
rect 698 388 699 392
rect 36 368 38 372
rect 1242 368 1257 371
rect 942 358 961 361
rect 1046 358 1062 361
rect 122 348 129 351
rect 154 348 161 351
rect 246 348 265 351
rect 270 348 278 351
rect 350 348 377 351
rect 62 338 65 348
rect 110 338 118 341
rect 142 338 150 341
rect 162 338 169 341
rect 238 341 241 348
rect 222 338 241 341
rect 350 338 353 348
rect 638 351 642 354
rect 814 352 818 354
rect 846 352 850 354
rect 638 348 649 351
rect 474 338 481 341
rect 646 338 649 348
rect 1718 348 1729 351
rect 1718 342 1721 348
rect 1922 348 1929 351
rect 2070 348 2078 351
rect 2470 348 2481 351
rect 2670 348 2689 351
rect 2470 342 2473 348
rect 678 338 689 341
rect 918 338 945 341
rect 1190 338 1198 341
rect 1534 338 1553 341
rect 1914 338 1921 341
rect 2006 332 2009 342
rect 2526 338 2537 341
rect 2594 338 2601 341
rect 2630 338 2638 341
rect 326 328 342 331
rect 422 328 433 331
rect 658 328 673 331
rect 1710 328 1721 331
rect 2374 328 2385 331
rect 2502 328 2521 331
rect 92 318 94 322
rect 1046 318 1062 321
rect 1562 318 1563 322
rect 1080 303 1082 307
rect 1086 303 1089 307
rect 1093 303 1096 307
rect 2104 303 2106 307
rect 2110 303 2113 307
rect 2117 303 2120 307
rect 2157 288 2158 292
rect 94 278 113 281
rect 30 268 41 271
rect 134 271 137 281
rect 542 278 553 281
rect 1086 281 1089 288
rect 1070 278 1089 281
rect 1270 278 1278 281
rect 134 268 142 271
rect 286 271 289 278
rect 230 268 241 271
rect 262 268 281 271
rect 286 268 297 271
rect 1302 268 1310 271
rect 1453 268 1454 272
rect 1538 268 1546 271
rect 1982 271 1986 274
rect 1982 268 1993 271
rect 2010 268 2017 271
rect 2194 268 2201 271
rect 2310 268 2326 271
rect 2550 268 2553 278
rect 38 262 41 268
rect 14 258 25 261
rect 54 258 73 261
rect 118 261 121 268
rect 118 258 129 261
rect 190 258 201 261
rect 310 261 313 268
rect 310 258 321 261
rect 542 261 545 268
rect 534 258 545 261
rect 694 258 713 261
rect 786 258 793 261
rect 942 258 961 261
rect 1046 261 1049 268
rect 1030 258 1049 261
rect 1082 258 1097 261
rect 1266 258 1273 261
rect 1334 258 1342 261
rect 1350 258 1358 261
rect 1382 258 1401 261
rect 1594 258 1601 261
rect 1798 258 1809 261
rect 1998 258 2014 261
rect 2182 258 2190 261
rect 2230 258 2249 261
rect 2290 258 2297 261
rect 2470 258 2486 261
rect 210 248 217 251
rect 294 251 297 258
rect 294 248 305 251
rect 310 248 321 251
rect 1230 248 1241 251
rect 1378 248 1382 252
rect 2130 248 2137 251
rect 2190 248 2201 251
rect 2230 248 2233 258
rect 2362 248 2366 252
rect 1342 241 1346 244
rect 1334 238 1346 241
rect 576 203 578 207
rect 582 203 585 207
rect 589 203 592 207
rect 1600 203 1602 207
rect 1606 203 1609 207
rect 1613 203 1616 207
rect 437 188 438 192
rect 653 188 654 192
rect 853 188 854 192
rect 917 188 918 192
rect 941 188 942 192
rect 2149 188 2150 192
rect 2466 188 2467 192
rect 540 168 542 172
rect 2182 166 2186 168
rect 698 158 702 162
rect 1046 158 1057 161
rect 1198 158 1209 161
rect 26 148 33 151
rect 150 148 161 151
rect 478 148 489 151
rect 606 148 614 151
rect 674 148 681 151
rect 690 148 697 151
rect 714 148 721 151
rect 950 148 969 151
rect 974 148 993 151
rect 1014 148 1025 151
rect 1070 148 1105 151
rect 1110 148 1137 151
rect 1142 148 1153 151
rect 1170 148 1177 151
rect 1222 151 1225 158
rect 1222 148 1233 151
rect 158 142 161 148
rect 6 138 25 141
rect 506 138 513 141
rect 630 141 633 148
rect 602 138 617 141
rect 622 138 633 141
rect 678 138 689 141
rect 742 138 761 141
rect 934 141 937 148
rect 926 138 937 141
rect 950 142 953 148
rect 1070 138 1073 148
rect 1878 148 1889 151
rect 1918 148 1929 151
rect 2058 148 2065 151
rect 2106 148 2113 151
rect 2174 148 2185 151
rect 2250 148 2257 151
rect 2326 148 2337 151
rect 2446 148 2462 151
rect 1554 138 1561 141
rect 1846 141 1849 148
rect 1886 142 1889 148
rect 1846 138 1857 141
rect 1926 138 1929 148
rect 2182 142 2185 148
rect 2358 138 2377 141
rect 2398 138 2406 141
rect 2446 138 2449 148
rect 22 128 25 138
rect 182 131 186 133
rect 158 128 169 131
rect 174 128 186 131
rect 198 132 202 136
rect 1054 132 1057 138
rect 422 128 430 131
rect 446 128 457 131
rect 490 128 497 131
rect 578 128 585 131
rect 1054 128 1062 132
rect 1350 128 1361 131
rect 1446 128 1457 131
rect 1462 128 1470 131
rect 1590 128 1617 131
rect 1622 128 1630 131
rect 1838 128 1849 131
rect 2306 128 2321 131
rect 2422 128 2425 138
rect 2534 128 2545 131
rect 741 118 742 122
rect 1213 118 1214 122
rect 2437 118 2438 122
rect 1080 103 1082 107
rect 1086 103 1089 107
rect 1093 103 1096 107
rect 2104 103 2106 107
rect 2110 103 2113 107
rect 2117 103 2120 107
rect 676 88 678 92
rect 930 88 931 92
rect 1173 88 1174 92
rect 1413 88 1414 92
rect 1586 88 1601 91
rect 2146 88 2161 91
rect 2618 88 2619 92
rect 62 78 73 81
rect 230 78 241 81
rect 246 72 249 81
rect 390 78 401 81
rect 406 72 409 81
rect 1006 78 1017 81
rect 1086 78 1102 81
rect 1198 78 1206 81
rect 1214 78 1222 81
rect 1006 72 1009 78
rect 46 58 54 61
rect 342 58 353 61
rect 390 61 393 68
rect 382 58 393 61
rect 694 62 697 71
rect 766 68 785 71
rect 790 68 798 71
rect 1034 68 1041 71
rect 1054 68 1065 71
rect 1334 71 1337 81
rect 1334 68 1353 71
rect 1374 68 1382 71
rect 1598 71 1602 74
rect 1942 72 1945 81
rect 1950 78 1961 81
rect 2022 78 2033 81
rect 2366 78 2377 81
rect 2382 78 2401 81
rect 2590 78 2598 81
rect 1574 68 1602 71
rect 2278 68 2286 71
rect 2422 68 2433 71
rect 2462 68 2481 71
rect 782 62 785 68
rect 1054 62 1057 68
rect 502 58 513 61
rect 566 58 598 61
rect 622 58 633 61
rect 726 58 761 61
rect 874 58 881 61
rect 1070 58 1081 61
rect 1474 58 1489 61
rect 1642 58 1657 61
rect 1838 58 1850 61
rect 1958 61 1961 68
rect 1958 58 1969 61
rect 2022 61 2025 68
rect 2014 58 2025 61
rect 2158 58 2166 61
rect 2430 62 2434 64
rect 2342 58 2353 61
rect 2358 58 2366 61
rect 2478 58 2494 61
rect 2502 58 2513 61
rect 2558 61 2561 68
rect 2558 58 2569 61
rect 2598 58 2606 61
rect 342 57 346 58
rect 502 57 506 58
rect 1270 52 1273 58
rect 1130 48 1132 52
rect 1186 48 1193 51
rect 1270 48 1279 52
rect 1382 51 1385 58
rect 1846 57 1850 58
rect 1382 48 1393 51
rect 1546 48 1548 52
rect 576 3 578 7
rect 582 3 585 7
rect 589 3 592 7
rect 1600 3 1602 7
rect 1606 3 1609 7
rect 1613 3 1616 7
<< m2contact >>
rect 578 1803 582 1807
rect 585 1803 589 1807
rect 1602 1803 1606 1807
rect 1609 1803 1613 1807
rect 510 1788 514 1792
rect 766 1788 770 1792
rect 790 1788 794 1792
rect 950 1788 954 1792
rect 974 1788 978 1792
rect 1102 1788 1106 1792
rect 1134 1788 1138 1792
rect 1238 1788 1242 1792
rect 1318 1788 1322 1792
rect 1438 1788 1442 1792
rect 1462 1788 1466 1792
rect 1486 1788 1490 1792
rect 1510 1788 1514 1792
rect 1518 1788 1522 1792
rect 1686 1788 1690 1792
rect 1694 1788 1698 1792
rect 1734 1788 1738 1792
rect 1894 1788 1898 1792
rect 2694 1788 2698 1792
rect 742 1778 746 1782
rect 2150 1778 2154 1782
rect 102 1768 106 1772
rect 894 1768 898 1772
rect 1142 1768 1146 1772
rect 1542 1768 1546 1772
rect 1830 1768 1834 1772
rect 2382 1768 2386 1772
rect 6 1758 10 1762
rect 62 1758 66 1762
rect 86 1758 90 1762
rect 2022 1758 2026 1762
rect 2054 1758 2058 1762
rect 2222 1758 2226 1762
rect 2230 1758 2234 1762
rect 2398 1758 2402 1762
rect 2670 1758 2674 1762
rect 30 1748 34 1752
rect 46 1748 50 1752
rect 182 1748 186 1752
rect 446 1748 450 1752
rect 494 1748 498 1752
rect 38 1738 42 1742
rect 54 1738 58 1742
rect 78 1738 82 1742
rect 102 1738 106 1742
rect 126 1738 130 1742
rect 214 1738 218 1742
rect 254 1738 258 1742
rect 294 1738 298 1742
rect 310 1738 314 1742
rect 366 1738 370 1742
rect 406 1738 410 1742
rect 582 1747 586 1751
rect 678 1748 682 1752
rect 750 1748 754 1752
rect 774 1748 778 1752
rect 830 1748 834 1752
rect 926 1748 930 1752
rect 934 1748 938 1752
rect 958 1748 962 1752
rect 1014 1748 1018 1752
rect 1078 1748 1082 1752
rect 1118 1748 1122 1752
rect 1206 1747 1210 1751
rect 1254 1748 1258 1752
rect 1262 1748 1266 1752
rect 1294 1748 1298 1752
rect 1358 1748 1362 1752
rect 1422 1748 1426 1752
rect 1446 1748 1450 1752
rect 1470 1748 1474 1752
rect 1494 1748 1498 1752
rect 1534 1748 1538 1752
rect 1606 1747 1610 1751
rect 1670 1748 1674 1752
rect 1710 1748 1714 1752
rect 1718 1748 1722 1752
rect 1774 1748 1778 1752
rect 1838 1748 1842 1752
rect 1870 1748 1874 1752
rect 1934 1748 1938 1752
rect 2006 1748 2010 1752
rect 2086 1747 2090 1751
rect 2174 1748 2178 1752
rect 2190 1748 2194 1752
rect 2206 1748 2210 1752
rect 2222 1748 2226 1752
rect 2254 1748 2258 1752
rect 454 1738 458 1742
rect 662 1738 666 1742
rect 910 1738 914 1742
rect 990 1738 994 1742
rect 1038 1738 1042 1742
rect 1278 1738 1282 1742
rect 1334 1738 1338 1742
rect 1646 1738 1650 1742
rect 1750 1738 1754 1742
rect 1838 1738 1842 1742
rect 1910 1738 1914 1742
rect 1998 1738 2002 1742
rect 2038 1738 2042 1742
rect 2070 1738 2074 1742
rect 2198 1738 2202 1742
rect 2310 1747 2314 1751
rect 2430 1748 2434 1752
rect 2470 1748 2474 1752
rect 2526 1748 2530 1752
rect 2230 1738 2234 1742
rect 2246 1738 2250 1742
rect 2262 1738 2266 1742
rect 2278 1738 2282 1742
rect 2294 1738 2298 1742
rect 2382 1738 2386 1742
rect 2422 1738 2426 1742
rect 2494 1738 2498 1742
rect 2502 1740 2506 1744
rect 2590 1747 2594 1751
rect 2670 1748 2674 1752
rect 2550 1738 2554 1742
rect 2574 1738 2578 1742
rect 6 1728 10 1732
rect 118 1728 122 1732
rect 158 1728 162 1732
rect 166 1728 170 1732
rect 254 1728 258 1732
rect 302 1728 306 1732
rect 334 1728 338 1732
rect 374 1728 378 1732
rect 30 1718 34 1722
rect 70 1718 74 1722
rect 78 1718 82 1722
rect 86 1718 90 1722
rect 102 1718 106 1722
rect 126 1718 130 1722
rect 142 1718 146 1722
rect 198 1718 202 1722
rect 278 1718 282 1722
rect 294 1718 298 1722
rect 326 1718 330 1722
rect 350 1718 354 1722
rect 390 1718 394 1722
rect 486 1728 490 1732
rect 822 1728 826 1732
rect 1206 1728 1210 1732
rect 1294 1728 1298 1732
rect 1654 1728 1658 1732
rect 1870 1728 1874 1732
rect 2054 1728 2058 1732
rect 2190 1728 2194 1732
rect 2278 1728 2282 1732
rect 2406 1728 2410 1732
rect 2430 1728 2434 1732
rect 2462 1728 2466 1732
rect 2486 1728 2490 1732
rect 2542 1728 2546 1732
rect 2550 1728 2554 1732
rect 2670 1728 2674 1732
rect 438 1718 442 1722
rect 470 1718 474 1722
rect 518 1718 522 1722
rect 718 1718 722 1722
rect 1070 1718 1074 1722
rect 1414 1718 1418 1722
rect 1662 1718 1666 1722
rect 1990 1718 1994 1722
rect 2398 1718 2402 1722
rect 2454 1718 2458 1722
rect 2478 1718 2482 1722
rect 2518 1718 2522 1722
rect 2558 1718 2562 1722
rect 2654 1718 2658 1722
rect 6 1708 10 1712
rect 166 1708 170 1712
rect 334 1708 338 1712
rect 374 1708 378 1712
rect 486 1708 490 1712
rect 1082 1703 1086 1707
rect 1089 1703 1093 1707
rect 2106 1703 2110 1707
rect 2113 1703 2117 1707
rect 46 1698 50 1702
rect 62 1698 66 1702
rect 158 1698 162 1702
rect 182 1698 186 1702
rect 342 1688 346 1692
rect 494 1688 498 1692
rect 542 1688 546 1692
rect 598 1688 602 1692
rect 654 1688 658 1692
rect 678 1688 682 1692
rect 1158 1688 1162 1692
rect 1198 1688 1202 1692
rect 1214 1688 1218 1692
rect 1358 1688 1362 1692
rect 1550 1688 1554 1692
rect 1670 1688 1674 1692
rect 1814 1688 1818 1692
rect 2062 1688 2066 1692
rect 2206 1688 2210 1692
rect 2350 1688 2354 1692
rect 2398 1688 2402 1692
rect 2638 1688 2642 1692
rect 62 1678 66 1682
rect 158 1678 162 1682
rect 174 1678 178 1682
rect 182 1678 186 1682
rect 238 1678 242 1682
rect 310 1678 314 1682
rect 382 1678 386 1682
rect 446 1678 450 1682
rect 70 1668 74 1672
rect 118 1668 122 1672
rect 254 1668 258 1672
rect 326 1668 330 1672
rect 342 1668 346 1672
rect 350 1668 354 1672
rect 398 1668 402 1672
rect 414 1668 418 1672
rect 518 1678 522 1682
rect 566 1678 570 1682
rect 622 1678 626 1682
rect 670 1678 674 1682
rect 710 1678 714 1682
rect 718 1678 722 1682
rect 958 1678 962 1682
rect 1062 1678 1066 1682
rect 1166 1678 1170 1682
rect 1206 1678 1210 1682
rect 1310 1678 1314 1682
rect 1350 1678 1354 1682
rect 1398 1678 1402 1682
rect 1534 1678 1538 1682
rect 1662 1678 1666 1682
rect 1718 1678 1722 1682
rect 1854 1678 1858 1682
rect 2054 1678 2058 1682
rect 2086 1678 2090 1682
rect 2102 1678 2106 1682
rect 2182 1678 2186 1682
rect 2270 1678 2274 1682
rect 2558 1678 2562 1682
rect 2590 1678 2594 1682
rect 494 1668 498 1672
rect 502 1668 506 1672
rect 518 1668 522 1672
rect 542 1668 546 1672
rect 582 1668 586 1672
rect 606 1668 610 1672
rect 646 1668 650 1672
rect 686 1668 690 1672
rect 734 1668 738 1672
rect 774 1668 778 1672
rect 822 1668 826 1672
rect 1006 1668 1010 1672
rect 1022 1668 1026 1672
rect 1078 1668 1082 1672
rect 1190 1668 1194 1672
rect 1294 1668 1298 1672
rect 1326 1668 1330 1672
rect 1366 1668 1370 1672
rect 1414 1668 1418 1672
rect 1446 1668 1450 1672
rect 6 1658 10 1662
rect 54 1658 58 1662
rect 86 1658 90 1662
rect 110 1658 114 1662
rect 142 1658 146 1662
rect 198 1658 202 1662
rect 230 1658 234 1662
rect 286 1658 290 1662
rect 342 1658 346 1662
rect 430 1658 434 1662
rect 510 1658 514 1662
rect 542 1658 546 1662
rect 550 1658 554 1662
rect 598 1658 602 1662
rect 726 1658 730 1662
rect 814 1658 818 1662
rect 894 1658 898 1662
rect 918 1658 922 1662
rect 974 1658 978 1662
rect 990 1658 994 1662
rect 998 1658 1002 1662
rect 1014 1658 1018 1662
rect 1094 1659 1098 1663
rect 1278 1659 1282 1663
rect 1342 1658 1346 1662
rect 1398 1658 1402 1662
rect 1702 1668 1706 1672
rect 1734 1668 1738 1672
rect 1838 1668 1842 1672
rect 1910 1668 1914 1672
rect 2086 1668 2090 1672
rect 2142 1668 2146 1672
rect 2174 1668 2178 1672
rect 2222 1668 2226 1672
rect 2230 1668 2234 1672
rect 2294 1668 2298 1672
rect 2326 1668 2330 1672
rect 2358 1668 2362 1672
rect 2390 1668 2394 1672
rect 1470 1658 1474 1662
rect 1486 1658 1490 1662
rect 1534 1658 1538 1662
rect 1582 1658 1586 1662
rect 1606 1658 1610 1662
rect 1678 1658 1682 1662
rect 1750 1659 1754 1663
rect 1822 1658 1826 1662
rect 1918 1658 1922 1662
rect 1982 1659 1986 1663
rect 2078 1658 2082 1662
rect 2102 1658 2106 1662
rect 2150 1658 2154 1662
rect 2182 1658 2186 1662
rect 2198 1658 2202 1662
rect 2270 1658 2274 1662
rect 2278 1658 2282 1662
rect 2294 1658 2298 1662
rect 2302 1658 2306 1662
rect 2310 1658 2314 1662
rect 2334 1658 2338 1662
rect 2366 1658 2370 1662
rect 2398 1658 2402 1662
rect 2414 1658 2418 1662
rect 2454 1668 2458 1672
rect 2462 1668 2466 1672
rect 2526 1668 2530 1672
rect 2574 1668 2578 1672
rect 2606 1668 2610 1672
rect 2622 1668 2626 1672
rect 2670 1668 2674 1672
rect 2446 1658 2450 1662
rect 2462 1658 2466 1662
rect 2486 1658 2490 1662
rect 2494 1658 2498 1662
rect 2518 1658 2522 1662
rect 2534 1658 2538 1662
rect 2542 1658 2546 1662
rect 2614 1658 2618 1662
rect 2678 1658 2682 1662
rect 30 1648 34 1652
rect 78 1648 82 1652
rect 278 1648 282 1652
rect 374 1648 378 1652
rect 438 1648 442 1652
rect 614 1648 618 1652
rect 2150 1648 2154 1652
rect 2246 1648 2250 1652
rect 2350 1648 2354 1652
rect 2366 1648 2370 1652
rect 2382 1648 2386 1652
rect 2486 1648 2490 1652
rect 2550 1648 2554 1652
rect 94 1638 98 1642
rect 134 1638 138 1642
rect 270 1638 274 1642
rect 422 1638 426 1642
rect 470 1638 474 1642
rect 550 1638 554 1642
rect 2030 1638 2034 1642
rect 2046 1638 2050 1642
rect 46 1618 50 1622
rect 86 1618 90 1622
rect 166 1618 170 1622
rect 206 1618 210 1622
rect 246 1618 250 1622
rect 286 1618 290 1622
rect 358 1618 362 1622
rect 390 1618 394 1622
rect 406 1618 410 1622
rect 1542 1618 1546 1622
rect 2558 1618 2562 1622
rect 2694 1618 2698 1622
rect 578 1603 582 1607
rect 585 1603 589 1607
rect 1602 1603 1606 1607
rect 1609 1603 1613 1607
rect 446 1588 450 1592
rect 710 1588 714 1592
rect 726 1588 730 1592
rect 766 1588 770 1592
rect 822 1588 826 1592
rect 886 1588 890 1592
rect 910 1588 914 1592
rect 1214 1588 1218 1592
rect 1326 1588 1330 1592
rect 1518 1588 1522 1592
rect 1566 1588 1570 1592
rect 1846 1588 1850 1592
rect 2310 1588 2314 1592
rect 2334 1588 2338 1592
rect 2414 1588 2418 1592
rect 2438 1588 2442 1592
rect 2478 1588 2482 1592
rect 2550 1588 2554 1592
rect 510 1578 514 1582
rect 2110 1578 2114 1582
rect 158 1568 162 1572
rect 294 1568 298 1572
rect 998 1568 1002 1572
rect 1358 1568 1362 1572
rect 1502 1568 1506 1572
rect 1590 1568 1594 1572
rect 1918 1568 1922 1572
rect 2182 1568 2186 1572
rect 134 1558 138 1562
rect 142 1558 146 1562
rect 254 1558 258 1562
rect 310 1558 314 1562
rect 438 1558 442 1562
rect 494 1558 498 1562
rect 846 1558 850 1562
rect 926 1558 930 1562
rect 950 1558 954 1562
rect 1014 1558 1018 1562
rect 1030 1558 1034 1562
rect 1046 1558 1050 1562
rect 1078 1558 1082 1562
rect 1718 1558 1722 1562
rect 22 1548 26 1552
rect 150 1548 154 1552
rect 278 1548 282 1552
rect 302 1548 306 1552
rect 318 1548 322 1552
rect 334 1548 338 1552
rect 350 1548 354 1552
rect 358 1548 362 1552
rect 422 1548 426 1552
rect 470 1548 474 1552
rect 502 1548 506 1552
rect 566 1548 570 1552
rect 646 1547 650 1551
rect 742 1548 746 1552
rect 750 1548 754 1552
rect 46 1538 50 1542
rect 94 1538 98 1542
rect 110 1538 114 1542
rect 118 1538 122 1542
rect 134 1538 138 1542
rect 206 1538 210 1542
rect 230 1538 234 1542
rect 390 1538 394 1542
rect 406 1538 410 1542
rect 430 1538 434 1542
rect 654 1538 658 1542
rect 662 1538 666 1542
rect 774 1538 778 1542
rect 838 1548 842 1552
rect 862 1548 866 1552
rect 870 1538 874 1542
rect 910 1548 914 1552
rect 1078 1548 1082 1552
rect 1174 1548 1178 1552
rect 1230 1548 1234 1552
rect 1270 1548 1274 1552
rect 1294 1548 1298 1552
rect 1374 1548 1378 1552
rect 1438 1547 1442 1551
rect 1470 1548 1474 1552
rect 1510 1548 1514 1552
rect 1542 1548 1546 1552
rect 1550 1548 1554 1552
rect 1654 1547 1658 1551
rect 1734 1548 1738 1552
rect 1750 1548 1754 1552
rect 1814 1558 1818 1562
rect 1878 1558 1882 1562
rect 1958 1558 1962 1562
rect 1998 1558 2002 1562
rect 2214 1558 2218 1562
rect 2278 1558 2282 1562
rect 2494 1558 2498 1562
rect 2566 1558 2570 1562
rect 2638 1558 2642 1562
rect 1838 1548 1842 1552
rect 1894 1548 1898 1552
rect 1926 1548 1930 1552
rect 1998 1548 2002 1552
rect 2046 1547 2050 1551
rect 2150 1548 2154 1552
rect 2182 1548 2186 1552
rect 2198 1548 2202 1552
rect 2222 1548 2226 1552
rect 2270 1548 2274 1552
rect 2294 1548 2298 1552
rect 2342 1548 2346 1552
rect 2366 1548 2370 1552
rect 2406 1548 2410 1552
rect 2430 1548 2434 1552
rect 2502 1548 2506 1552
rect 2534 1548 2538 1552
rect 2550 1548 2554 1552
rect 2574 1548 2578 1552
rect 902 1538 906 1542
rect 934 1538 938 1542
rect 998 1538 1002 1542
rect 1070 1538 1074 1542
rect 1094 1538 1098 1542
rect 1110 1538 1114 1542
rect 1198 1538 1202 1542
rect 1342 1538 1346 1542
rect 1382 1538 1386 1542
rect 1518 1538 1522 1542
rect 1534 1538 1538 1542
rect 1646 1538 1650 1542
rect 1670 1538 1674 1542
rect 1686 1538 1690 1542
rect 1702 1538 1706 1542
rect 1750 1538 1754 1542
rect 1774 1538 1778 1542
rect 1790 1538 1794 1542
rect 1798 1538 1802 1542
rect 1870 1538 1874 1542
rect 1902 1538 1906 1542
rect 1934 1538 1938 1542
rect 1974 1538 1978 1542
rect 1998 1538 2002 1542
rect 2014 1538 2018 1542
rect 2030 1538 2034 1542
rect 2158 1538 2162 1542
rect 2190 1538 2194 1542
rect 2206 1538 2210 1542
rect 2222 1538 2226 1542
rect 2350 1538 2354 1542
rect 2398 1538 2402 1542
rect 2462 1538 2466 1542
rect 2526 1538 2530 1542
rect 2542 1538 2546 1542
rect 2654 1538 2658 1542
rect 2678 1538 2682 1542
rect 6 1528 10 1532
rect 70 1528 74 1532
rect 78 1528 82 1532
rect 190 1528 194 1532
rect 198 1528 202 1532
rect 262 1528 266 1532
rect 278 1528 282 1532
rect 382 1528 386 1532
rect 406 1528 410 1532
rect 470 1528 474 1532
rect 894 1528 898 1532
rect 958 1528 962 1532
rect 982 1528 986 1532
rect 1022 1528 1026 1532
rect 1334 1528 1338 1532
rect 1366 1528 1370 1532
rect 1406 1528 1410 1532
rect 1686 1528 1690 1532
rect 1766 1528 1770 1532
rect 1822 1528 1826 1532
rect 1838 1528 1842 1532
rect 1846 1528 1850 1532
rect 1926 1528 1930 1532
rect 1990 1528 1994 1532
rect 2166 1528 2170 1532
rect 2262 1528 2266 1532
rect 2286 1528 2290 1532
rect 2326 1528 2330 1532
rect 2422 1528 2426 1532
rect 2446 1528 2450 1532
rect 2478 1528 2482 1532
rect 2486 1528 2490 1532
rect 2510 1528 2514 1532
rect 2590 1528 2594 1532
rect 2614 1528 2618 1532
rect 2686 1528 2690 1532
rect 38 1518 42 1522
rect 62 1518 66 1522
rect 102 1518 106 1522
rect 110 1518 114 1522
rect 118 1518 122 1522
rect 182 1518 186 1522
rect 254 1518 258 1522
rect 270 1518 274 1522
rect 422 1518 426 1522
rect 710 1518 714 1522
rect 726 1518 730 1522
rect 798 1518 802 1522
rect 966 1518 970 1522
rect 1078 1518 1082 1522
rect 1118 1518 1122 1522
rect 1326 1518 1330 1522
rect 1806 1518 1810 1522
rect 2134 1518 2138 1522
rect 2246 1518 2250 1522
rect 2518 1518 2522 1522
rect 2662 1518 2666 1522
rect 6 1508 10 1512
rect 70 1508 74 1512
rect 1082 1503 1086 1507
rect 1089 1503 1093 1507
rect 2106 1503 2110 1507
rect 2113 1503 2117 1507
rect 38 1488 42 1492
rect 54 1488 58 1492
rect 118 1488 122 1492
rect 198 1488 202 1492
rect 510 1488 514 1492
rect 630 1488 634 1492
rect 742 1488 746 1492
rect 846 1488 850 1492
rect 950 1488 954 1492
rect 1222 1488 1226 1492
rect 1398 1488 1402 1492
rect 1582 1488 1586 1492
rect 1710 1488 1714 1492
rect 1974 1488 1978 1492
rect 2326 1488 2330 1492
rect 2358 1488 2362 1492
rect 2382 1488 2386 1492
rect 2478 1488 2482 1492
rect 2694 1488 2698 1492
rect 6 1478 10 1482
rect 134 1478 138 1482
rect 262 1478 266 1482
rect 294 1478 298 1482
rect 438 1478 442 1482
rect 462 1478 466 1482
rect 510 1478 514 1482
rect 574 1478 578 1482
rect 606 1478 610 1482
rect 638 1478 642 1482
rect 958 1478 962 1482
rect 1022 1478 1026 1482
rect 1054 1478 1058 1482
rect 1102 1478 1106 1482
rect 1118 1478 1122 1482
rect 1214 1478 1218 1482
rect 1286 1478 1290 1482
rect 1358 1478 1362 1482
rect 1366 1478 1370 1482
rect 1494 1478 1498 1482
rect 1718 1478 1722 1482
rect 1822 1478 1826 1482
rect 1854 1478 1858 1482
rect 1862 1478 1866 1482
rect 1918 1478 1922 1482
rect 2070 1478 2074 1482
rect 2078 1478 2082 1482
rect 2166 1478 2170 1482
rect 2262 1478 2266 1482
rect 2302 1478 2306 1482
rect 2390 1478 2394 1482
rect 2398 1478 2402 1482
rect 2430 1478 2434 1482
rect 2486 1478 2490 1482
rect 2590 1478 2594 1482
rect 2646 1478 2650 1482
rect 62 1468 66 1472
rect 94 1468 98 1472
rect 198 1468 202 1472
rect 206 1468 210 1472
rect 246 1468 250 1472
rect 278 1468 282 1472
rect 614 1468 618 1472
rect 654 1468 658 1472
rect 822 1468 826 1472
rect 854 1468 858 1472
rect 870 1468 874 1472
rect 958 1468 962 1472
rect 1094 1468 1098 1472
rect 1126 1468 1130 1472
rect 1150 1468 1154 1472
rect 1206 1468 1210 1472
rect 1318 1468 1322 1472
rect 1342 1468 1346 1472
rect 1382 1468 1386 1472
rect 1406 1468 1410 1472
rect 1430 1468 1434 1472
rect 1446 1468 1450 1472
rect 1734 1468 1738 1472
rect 1782 1468 1786 1472
rect 22 1458 26 1462
rect 38 1458 42 1462
rect 54 1458 58 1462
rect 86 1458 90 1462
rect 102 1458 106 1462
rect 118 1458 122 1462
rect 166 1458 170 1462
rect 214 1458 218 1462
rect 230 1458 234 1462
rect 238 1458 242 1462
rect 270 1458 274 1462
rect 326 1459 330 1463
rect 358 1458 362 1462
rect 422 1458 426 1462
rect 438 1458 442 1462
rect 502 1458 506 1462
rect 550 1458 554 1462
rect 678 1458 682 1462
rect 702 1458 706 1462
rect 774 1458 778 1462
rect 798 1458 802 1462
rect 894 1458 898 1462
rect 918 1458 922 1462
rect 998 1458 1002 1462
rect 1038 1458 1042 1462
rect 1078 1458 1082 1462
rect 1118 1458 1122 1462
rect 1182 1458 1186 1462
rect 1278 1458 1282 1462
rect 1422 1458 1426 1462
rect 1438 1458 1442 1462
rect 1518 1458 1522 1462
rect 1534 1458 1538 1462
rect 1598 1458 1602 1462
rect 1654 1458 1658 1462
rect 1670 1458 1674 1462
rect 1806 1466 1810 1470
rect 1814 1468 1818 1472
rect 1854 1468 1858 1472
rect 1886 1468 1890 1472
rect 1934 1468 1938 1472
rect 2030 1468 2034 1472
rect 2118 1468 2122 1472
rect 2134 1468 2138 1472
rect 2182 1468 2186 1472
rect 2230 1468 2234 1472
rect 2254 1468 2258 1472
rect 2286 1468 2290 1472
rect 2334 1468 2338 1472
rect 2518 1468 2522 1472
rect 2526 1468 2530 1472
rect 1774 1458 1778 1462
rect 1790 1458 1794 1462
rect 1878 1458 1882 1462
rect 1894 1458 1898 1462
rect 1910 1458 1914 1462
rect 1934 1458 1938 1462
rect 1942 1458 1946 1462
rect 1966 1458 1970 1462
rect 2038 1459 2042 1463
rect 2094 1458 2098 1462
rect 2142 1458 2146 1462
rect 2222 1458 2226 1462
rect 2230 1458 2234 1462
rect 2278 1458 2282 1462
rect 2286 1458 2290 1462
rect 2310 1458 2314 1462
rect 2374 1458 2378 1462
rect 2414 1458 2418 1462
rect 2430 1458 2434 1462
rect 2446 1458 2450 1462
rect 2470 1458 2474 1462
rect 2510 1458 2514 1462
rect 2542 1458 2546 1462
rect 2574 1466 2578 1470
rect 2582 1468 2586 1472
rect 2638 1468 2642 1472
rect 2702 1478 2706 1482
rect 2662 1468 2666 1472
rect 2686 1468 2690 1472
rect 2590 1458 2594 1462
rect 2614 1458 2618 1462
rect 2622 1458 2626 1462
rect 2630 1458 2634 1462
rect 2646 1458 2650 1462
rect 54 1448 58 1452
rect 86 1448 90 1452
rect 102 1448 106 1452
rect 134 1448 138 1452
rect 182 1448 186 1452
rect 230 1448 234 1452
rect 534 1448 538 1452
rect 982 1448 986 1452
rect 1030 1448 1034 1452
rect 1062 1448 1066 1452
rect 1174 1448 1178 1452
rect 1758 1448 1762 1452
rect 1910 1448 1914 1452
rect 2102 1448 2106 1452
rect 2206 1448 2210 1452
rect 2398 1448 2402 1452
rect 2438 1448 2442 1452
rect 2494 1448 2498 1452
rect 2526 1448 2530 1452
rect 2614 1448 2618 1452
rect 2686 1448 2690 1452
rect 158 1438 162 1442
rect 734 1438 738 1442
rect 838 1438 842 1442
rect 1022 1438 1026 1442
rect 1182 1438 1186 1442
rect 1190 1438 1194 1442
rect 1878 1438 1882 1442
rect 2238 1438 2242 1442
rect 2454 1438 2458 1442
rect 2510 1438 2514 1442
rect 1934 1428 1938 1432
rect 14 1418 18 1422
rect 166 1418 170 1422
rect 262 1418 266 1422
rect 294 1418 298 1422
rect 390 1418 394 1422
rect 950 1418 954 1422
rect 1134 1418 1138 1422
rect 1182 1418 1186 1422
rect 1326 1418 1330 1422
rect 1358 1418 1362 1422
rect 2198 1418 2202 1422
rect 2446 1418 2450 1422
rect 578 1403 582 1407
rect 585 1403 589 1407
rect 1602 1403 1606 1407
rect 1609 1403 1613 1407
rect 22 1388 26 1392
rect 214 1388 218 1392
rect 558 1388 562 1392
rect 622 1388 626 1392
rect 854 1388 858 1392
rect 886 1388 890 1392
rect 926 1388 930 1392
rect 1286 1388 1290 1392
rect 1382 1388 1386 1392
rect 1670 1388 1674 1392
rect 1782 1388 1786 1392
rect 2022 1388 2026 1392
rect 2166 1388 2170 1392
rect 2190 1388 2194 1392
rect 2214 1388 2218 1392
rect 2230 1388 2234 1392
rect 2278 1388 2282 1392
rect 2302 1388 2306 1392
rect 2550 1388 2554 1392
rect 2678 1388 2682 1392
rect 1958 1378 1962 1382
rect 2382 1378 2386 1382
rect 14 1368 18 1372
rect 150 1368 154 1372
rect 222 1368 226 1372
rect 766 1368 770 1372
rect 1518 1368 1522 1372
rect 1774 1368 1778 1372
rect 1982 1368 1986 1372
rect 2006 1368 2010 1372
rect 2342 1368 2346 1372
rect 2590 1368 2594 1372
rect 70 1358 74 1362
rect 166 1358 170 1362
rect 310 1358 314 1362
rect 342 1358 346 1362
rect 22 1348 26 1352
rect 94 1348 98 1352
rect 126 1348 130 1352
rect 214 1348 218 1352
rect 278 1348 282 1352
rect 502 1358 506 1362
rect 998 1358 1002 1362
rect 1022 1358 1026 1362
rect 1758 1358 1762 1362
rect 1966 1358 1970 1362
rect 2014 1358 2018 1362
rect 2062 1358 2066 1362
rect 2078 1358 2082 1362
rect 2174 1358 2178 1362
rect 2198 1358 2202 1362
rect 2222 1358 2226 1362
rect 2270 1358 2274 1362
rect 2286 1358 2290 1362
rect 2310 1358 2314 1362
rect 2318 1358 2322 1362
rect 2334 1358 2338 1362
rect 2358 1358 2362 1362
rect 358 1348 362 1352
rect 422 1347 426 1351
rect 454 1348 458 1352
rect 510 1348 514 1352
rect 558 1348 562 1352
rect 670 1348 674 1352
rect 742 1348 746 1352
rect 790 1348 794 1352
rect 870 1348 874 1352
rect 894 1348 898 1352
rect 1062 1348 1066 1352
rect 1102 1348 1106 1352
rect 1126 1348 1130 1352
rect 1166 1348 1170 1352
rect 1246 1348 1250 1352
rect 1342 1348 1346 1352
rect 1414 1348 1418 1352
rect 1438 1348 1442 1352
rect 1478 1348 1482 1352
rect 1566 1347 1570 1351
rect 1742 1348 1746 1352
rect 1766 1348 1770 1352
rect 1790 1348 1794 1352
rect 1822 1348 1826 1352
rect 1854 1348 1858 1352
rect 1886 1348 1890 1352
rect 1942 1348 1946 1352
rect 1958 1348 1962 1352
rect 1974 1348 1978 1352
rect 2094 1348 2098 1352
rect 2150 1348 2154 1352
rect 2206 1348 2210 1352
rect 2382 1348 2386 1352
rect 2406 1348 2410 1352
rect 2414 1348 2418 1352
rect 2454 1358 2458 1362
rect 2494 1358 2498 1362
rect 2566 1358 2570 1362
rect 2574 1358 2578 1362
rect 2454 1348 2458 1352
rect 2478 1348 2482 1352
rect 2494 1348 2498 1352
rect 2510 1348 2514 1352
rect 2526 1348 2530 1352
rect 2550 1348 2554 1352
rect 2590 1348 2594 1352
rect 2606 1348 2610 1352
rect 2622 1348 2626 1352
rect 2646 1348 2650 1352
rect 2662 1348 2666 1352
rect 54 1338 58 1342
rect 70 1338 74 1342
rect 86 1338 90 1342
rect 126 1338 130 1342
rect 150 1338 154 1342
rect 166 1338 170 1342
rect 182 1338 186 1342
rect 286 1338 290 1342
rect 294 1338 298 1342
rect 318 1338 322 1342
rect 374 1338 378 1342
rect 390 1338 394 1342
rect 406 1338 410 1342
rect 518 1338 522 1342
rect 526 1340 530 1344
rect 582 1338 586 1342
rect 702 1338 706 1342
rect 830 1338 834 1342
rect 982 1338 986 1342
rect 1006 1338 1010 1342
rect 1070 1338 1074 1342
rect 1142 1340 1146 1344
rect 1182 1338 1186 1342
rect 1270 1338 1274 1342
rect 1582 1338 1586 1342
rect 1614 1338 1618 1342
rect 1686 1338 1690 1342
rect 1814 1338 1818 1342
rect 1838 1338 1842 1342
rect 1934 1338 1938 1342
rect 1982 1338 1986 1342
rect 2030 1338 2034 1342
rect 2086 1338 2090 1342
rect 2102 1338 2106 1342
rect 2142 1338 2146 1342
rect 2158 1338 2162 1342
rect 2182 1338 2186 1342
rect 2198 1338 2202 1342
rect 2246 1338 2250 1342
rect 2270 1338 2274 1342
rect 2286 1338 2290 1342
rect 2318 1338 2322 1342
rect 2334 1338 2338 1342
rect 2462 1338 2466 1342
rect 2470 1338 2474 1342
rect 2502 1338 2506 1342
rect 2534 1338 2538 1342
rect 2542 1338 2546 1342
rect 2598 1338 2602 1342
rect 2606 1338 2610 1342
rect 2654 1338 2658 1342
rect 2686 1338 2690 1342
rect 62 1328 66 1332
rect 94 1328 98 1332
rect 110 1328 114 1332
rect 174 1328 178 1332
rect 254 1328 258 1332
rect 606 1328 610 1332
rect 878 1328 882 1332
rect 990 1328 994 1332
rect 1030 1328 1034 1332
rect 1078 1328 1082 1332
rect 1110 1328 1114 1332
rect 1126 1328 1130 1332
rect 1350 1328 1354 1332
rect 1942 1328 1946 1332
rect 2006 1328 2010 1332
rect 2038 1328 2042 1332
rect 2054 1328 2058 1332
rect 2070 1328 2074 1332
rect 2126 1328 2130 1332
rect 2238 1328 2242 1332
rect 2366 1328 2370 1332
rect 2390 1328 2394 1332
rect 2430 1328 2434 1332
rect 2526 1328 2530 1332
rect 2622 1328 2626 1332
rect 86 1318 90 1322
rect 190 1318 194 1322
rect 246 1318 250 1322
rect 262 1318 266 1322
rect 302 1318 306 1322
rect 486 1318 490 1322
rect 622 1318 626 1322
rect 726 1318 730 1322
rect 750 1318 754 1322
rect 1054 1318 1058 1322
rect 1158 1318 1162 1322
rect 1174 1318 1178 1322
rect 1190 1318 1194 1322
rect 1286 1318 1290 1322
rect 1502 1318 1506 1322
rect 1870 1318 1874 1322
rect 1902 1318 1906 1322
rect 2134 1318 2138 1322
rect 2262 1318 2266 1322
rect 2278 1318 2282 1322
rect 2302 1318 2306 1322
rect 2398 1318 2402 1322
rect 30 1308 34 1312
rect 110 1308 114 1312
rect 150 1308 154 1312
rect 1082 1303 1086 1307
rect 1089 1303 1093 1307
rect 2106 1303 2110 1307
rect 2113 1303 2117 1307
rect 94 1298 98 1302
rect 206 1298 210 1302
rect 278 1298 282 1302
rect 894 1298 898 1302
rect 38 1288 42 1292
rect 78 1288 82 1292
rect 230 1288 234 1292
rect 326 1288 330 1292
rect 534 1288 538 1292
rect 574 1288 578 1292
rect 678 1288 682 1292
rect 926 1288 930 1292
rect 1102 1288 1106 1292
rect 1110 1288 1114 1292
rect 1198 1288 1202 1292
rect 1278 1288 1282 1292
rect 1478 1288 1482 1292
rect 1590 1288 1594 1292
rect 1638 1288 1642 1292
rect 1742 1288 1746 1292
rect 1758 1288 1762 1292
rect 1806 1288 1810 1292
rect 1862 1288 1866 1292
rect 1910 1288 1914 1292
rect 2062 1288 2066 1292
rect 2286 1288 2290 1292
rect 2318 1288 2322 1292
rect 2454 1288 2458 1292
rect 2566 1288 2570 1292
rect 2622 1288 2626 1292
rect 54 1268 58 1272
rect 70 1268 74 1272
rect 94 1278 98 1282
rect 126 1278 130 1282
rect 206 1278 210 1282
rect 238 1278 242 1282
rect 246 1278 250 1282
rect 278 1278 282 1282
rect 358 1278 362 1282
rect 382 1278 386 1282
rect 622 1278 626 1282
rect 782 1278 786 1282
rect 918 1278 922 1282
rect 934 1278 938 1282
rect 1062 1278 1066 1282
rect 1206 1278 1210 1282
rect 1230 1278 1234 1282
rect 1470 1278 1474 1282
rect 1502 1278 1506 1282
rect 1542 1278 1546 1282
rect 1598 1278 1602 1282
rect 2054 1278 2058 1282
rect 2110 1278 2114 1282
rect 2150 1278 2154 1282
rect 2174 1278 2178 1282
rect 2206 1278 2210 1282
rect 2230 1278 2234 1282
rect 2350 1278 2354 1282
rect 2358 1278 2362 1282
rect 2382 1278 2386 1282
rect 2430 1278 2434 1282
rect 2478 1278 2482 1282
rect 2502 1278 2506 1282
rect 2534 1278 2538 1282
rect 2550 1278 2554 1282
rect 2558 1278 2562 1282
rect 2590 1278 2594 1282
rect 2598 1278 2602 1282
rect 190 1268 194 1272
rect 214 1268 218 1272
rect 262 1268 266 1272
rect 286 1268 290 1272
rect 326 1268 330 1272
rect 342 1268 346 1272
rect 390 1268 394 1272
rect 422 1268 426 1272
rect 438 1268 442 1272
rect 454 1268 458 1272
rect 542 1268 546 1272
rect 614 1268 618 1272
rect 630 1268 634 1272
rect 654 1268 658 1272
rect 766 1268 770 1272
rect 790 1268 794 1272
rect 838 1268 842 1272
rect 846 1268 850 1272
rect 974 1268 978 1272
rect 62 1258 66 1262
rect 190 1258 194 1262
rect 278 1258 282 1262
rect 302 1258 306 1262
rect 318 1258 322 1262
rect 350 1258 354 1262
rect 470 1259 474 1263
rect 502 1258 506 1262
rect 550 1258 554 1262
rect 582 1258 586 1262
rect 646 1258 650 1262
rect 662 1258 666 1262
rect 750 1259 754 1263
rect 806 1258 810 1262
rect 846 1258 850 1262
rect 982 1266 986 1270
rect 1006 1268 1010 1272
rect 1022 1268 1026 1272
rect 1126 1268 1130 1272
rect 1190 1268 1194 1272
rect 1238 1268 1242 1272
rect 1302 1268 1306 1272
rect 1350 1268 1354 1272
rect 1398 1268 1402 1272
rect 1414 1268 1418 1272
rect 1446 1268 1450 1272
rect 1454 1268 1458 1272
rect 1462 1268 1466 1272
rect 1486 1268 1490 1272
rect 1526 1268 1530 1272
rect 1550 1268 1554 1272
rect 1582 1268 1586 1272
rect 1678 1268 1682 1272
rect 1766 1268 1770 1272
rect 1822 1268 1826 1272
rect 966 1258 970 1262
rect 998 1258 1002 1262
rect 1038 1258 1042 1262
rect 1142 1258 1146 1262
rect 1182 1258 1186 1262
rect 1246 1258 1250 1262
rect 1286 1258 1290 1262
rect 1334 1258 1338 1262
rect 1390 1258 1394 1262
rect 1478 1258 1482 1262
rect 1510 1258 1514 1262
rect 1542 1258 1546 1262
rect 1582 1258 1586 1262
rect 1598 1258 1602 1262
rect 1686 1258 1690 1262
rect 1798 1258 1802 1262
rect 1854 1258 1858 1262
rect 1886 1268 1890 1272
rect 1918 1268 1922 1272
rect 2078 1268 2082 1272
rect 2094 1268 2098 1272
rect 2150 1268 2154 1272
rect 2174 1268 2178 1272
rect 2222 1268 2226 1272
rect 2254 1268 2258 1272
rect 2326 1268 2330 1272
rect 2510 1268 2514 1272
rect 2574 1268 2578 1272
rect 2614 1268 2618 1272
rect 2638 1278 2642 1282
rect 2670 1268 2674 1272
rect 2694 1268 2698 1272
rect 1942 1258 1946 1262
rect 1990 1258 1994 1262
rect 2022 1259 2026 1263
rect 2070 1258 2074 1262
rect 2118 1258 2122 1262
rect 2142 1258 2146 1262
rect 2166 1258 2170 1262
rect 2182 1258 2186 1262
rect 2198 1258 2202 1262
rect 2222 1258 2226 1262
rect 2246 1258 2250 1262
rect 2334 1258 2338 1262
rect 2374 1258 2378 1262
rect 2406 1258 2410 1262
rect 2446 1258 2450 1262
rect 2486 1258 2490 1262
rect 2582 1258 2586 1262
rect 166 1248 170 1252
rect 310 1248 314 1252
rect 398 1248 402 1252
rect 414 1248 418 1252
rect 1022 1248 1026 1252
rect 1054 1248 1058 1252
rect 1110 1248 1114 1252
rect 1134 1248 1138 1252
rect 1262 1248 1266 1252
rect 1422 1248 1426 1252
rect 1526 1248 1530 1252
rect 1574 1248 1578 1252
rect 1750 1248 1754 1252
rect 1806 1248 1810 1252
rect 1862 1248 1866 1252
rect 1950 1248 1954 1252
rect 2086 1248 2090 1252
rect 2270 1248 2274 1252
rect 2430 1248 2434 1252
rect 2438 1248 2442 1252
rect 2670 1248 2674 1252
rect 686 1238 690 1242
rect 702 1238 706 1242
rect 814 1238 818 1242
rect 1150 1238 1154 1242
rect 1166 1238 1170 1242
rect 1382 1238 1386 1242
rect 1902 1238 1906 1242
rect 1934 1238 1938 1242
rect 2382 1238 2386 1242
rect 1142 1228 1146 1232
rect 2406 1228 2410 1232
rect 902 1218 906 1222
rect 1014 1218 1018 1222
rect 1214 1218 1218 1222
rect 1534 1218 1538 1222
rect 1782 1218 1786 1222
rect 1838 1218 1842 1222
rect 1942 1218 1946 1222
rect 1958 1218 1962 1222
rect 2342 1218 2346 1222
rect 578 1203 582 1207
rect 585 1203 589 1207
rect 1602 1203 1606 1207
rect 1609 1203 1613 1207
rect 182 1188 186 1192
rect 270 1188 274 1192
rect 766 1188 770 1192
rect 1254 1188 1258 1192
rect 1566 1188 1570 1192
rect 1694 1188 1698 1192
rect 2134 1188 2138 1192
rect 2166 1188 2170 1192
rect 2238 1188 2242 1192
rect 2646 1188 2650 1192
rect 302 1168 306 1172
rect 462 1168 466 1172
rect 758 1168 762 1172
rect 1294 1168 1298 1172
rect 1318 1168 1322 1172
rect 1678 1168 1682 1172
rect 1982 1168 1986 1172
rect 198 1158 202 1162
rect 222 1158 226 1162
rect 286 1158 290 1162
rect 318 1158 322 1162
rect 1094 1158 1098 1162
rect 1326 1158 1330 1162
rect 1342 1158 1346 1162
rect 1390 1158 1394 1162
rect 1502 1158 1506 1162
rect 1518 1158 1522 1162
rect 110 1148 114 1152
rect 182 1148 186 1152
rect 238 1148 242 1152
rect 270 1148 274 1152
rect 302 1148 306 1152
rect 318 1148 322 1152
rect 342 1148 346 1152
rect 358 1148 362 1152
rect 390 1147 394 1151
rect 422 1148 426 1152
rect 534 1148 538 1152
rect 558 1148 562 1152
rect 606 1148 610 1152
rect 678 1148 682 1152
rect 702 1148 706 1152
rect 750 1148 754 1152
rect 830 1148 834 1152
rect 870 1148 874 1152
rect 918 1147 922 1151
rect 1022 1148 1026 1152
rect 1062 1148 1066 1152
rect 1230 1148 1234 1152
rect 1254 1148 1258 1152
rect 1286 1148 1290 1152
rect 1302 1148 1306 1152
rect 1342 1148 1346 1152
rect 1358 1148 1362 1152
rect 1406 1148 1410 1152
rect 1446 1148 1450 1152
rect 1494 1148 1498 1152
rect 1590 1148 1594 1152
rect 54 1138 58 1142
rect 118 1138 122 1142
rect 174 1138 178 1142
rect 206 1138 210 1142
rect 214 1138 218 1142
rect 222 1138 226 1142
rect 262 1138 266 1142
rect 294 1138 298 1142
rect 334 1138 338 1142
rect 350 1138 354 1142
rect 374 1138 378 1142
rect 462 1138 466 1142
rect 478 1138 482 1142
rect 630 1138 634 1142
rect 854 1138 858 1142
rect 886 1138 890 1142
rect 902 1138 906 1142
rect 1046 1138 1050 1142
rect 1134 1138 1138 1142
rect 1174 1138 1178 1142
rect 1350 1138 1354 1142
rect 1366 1138 1370 1142
rect 1398 1138 1402 1142
rect 1414 1138 1418 1142
rect 1438 1138 1442 1142
rect 1470 1138 1474 1142
rect 1486 1138 1490 1142
rect 1502 1138 1506 1142
rect 1526 1138 1530 1142
rect 1630 1147 1634 1151
rect 1742 1148 1746 1152
rect 1798 1148 1802 1152
rect 1838 1147 1842 1151
rect 1934 1147 1938 1151
rect 2046 1148 2050 1152
rect 2150 1158 2154 1162
rect 2182 1158 2186 1162
rect 2222 1158 2226 1162
rect 2302 1158 2306 1162
rect 2374 1158 2378 1162
rect 2430 1158 2434 1162
rect 2478 1158 2482 1162
rect 2630 1158 2634 1162
rect 2662 1158 2666 1162
rect 2670 1158 2674 1162
rect 2126 1148 2130 1152
rect 2214 1148 2218 1152
rect 2238 1148 2242 1152
rect 2310 1148 2314 1152
rect 2350 1148 2354 1152
rect 2390 1148 2394 1152
rect 2478 1148 2482 1152
rect 2510 1148 2514 1152
rect 2534 1148 2538 1152
rect 2542 1148 2546 1152
rect 2558 1148 2562 1152
rect 2582 1148 2586 1152
rect 2630 1148 2634 1152
rect 1646 1138 1650 1142
rect 1806 1138 1810 1142
rect 1822 1138 1826 1142
rect 1918 1138 1922 1142
rect 1966 1138 1970 1142
rect 2006 1138 2010 1142
rect 2094 1138 2098 1142
rect 2246 1138 2250 1142
rect 2254 1138 2258 1142
rect 2262 1140 2266 1144
rect 2286 1138 2290 1142
rect 2358 1138 2362 1142
rect 2374 1138 2378 1142
rect 2414 1138 2418 1142
rect 2454 1138 2458 1142
rect 2462 1138 2466 1142
rect 2502 1138 2506 1142
rect 2574 1138 2578 1142
rect 2606 1138 2610 1142
rect 2630 1138 2634 1142
rect 2638 1138 2642 1142
rect 2702 1138 2706 1142
rect 6 1128 10 1132
rect 38 1128 42 1132
rect 78 1128 82 1132
rect 110 1128 114 1132
rect 494 1128 498 1132
rect 638 1128 642 1132
rect 886 1128 890 1132
rect 990 1128 994 1132
rect 998 1128 1002 1132
rect 1006 1128 1010 1132
rect 1078 1128 1082 1132
rect 1110 1128 1114 1132
rect 1126 1128 1130 1132
rect 1166 1128 1170 1132
rect 1206 1128 1210 1132
rect 1222 1127 1226 1131
rect 1238 1128 1242 1132
rect 1262 1128 1266 1132
rect 1318 1128 1322 1132
rect 1382 1128 1386 1132
rect 1422 1128 1426 1132
rect 1462 1128 1466 1132
rect 1734 1128 1738 1132
rect 2062 1128 2066 1132
rect 2094 1128 2098 1132
rect 2158 1128 2162 1132
rect 2190 1128 2194 1132
rect 2214 1128 2218 1132
rect 2326 1128 2330 1132
rect 2526 1128 2530 1132
rect 2550 1128 2554 1132
rect 2574 1128 2578 1132
rect 2598 1128 2602 1132
rect 62 1118 66 1122
rect 254 1118 258 1122
rect 590 1118 594 1122
rect 774 1118 778 1122
rect 982 1118 986 1122
rect 1030 1118 1034 1122
rect 1070 1118 1074 1122
rect 1118 1118 1122 1122
rect 1142 1118 1146 1122
rect 1182 1118 1186 1122
rect 1374 1118 1378 1122
rect 1430 1118 1434 1122
rect 1478 1118 1482 1122
rect 1550 1118 1554 1122
rect 1710 1118 1714 1122
rect 1734 1118 1738 1122
rect 1774 1118 1778 1122
rect 1902 1118 1906 1122
rect 1998 1118 2002 1122
rect 2014 1118 2018 1122
rect 2070 1118 2074 1122
rect 2278 1118 2282 1122
rect 2318 1118 2322 1122
rect 2342 1118 2346 1122
rect 2366 1118 2370 1122
rect 2406 1118 2410 1122
rect 2430 1118 2434 1122
rect 2438 1118 2442 1122
rect 2494 1118 2498 1122
rect 2518 1118 2522 1122
rect 2678 1118 2682 1122
rect 38 1108 42 1112
rect 46 1108 50 1112
rect 78 1108 82 1112
rect 126 1108 130 1112
rect 1082 1103 1086 1107
rect 1089 1103 1093 1107
rect 2106 1103 2110 1107
rect 2113 1103 2117 1107
rect 150 1098 154 1102
rect 214 1098 218 1102
rect 30 1088 34 1092
rect 102 1088 106 1092
rect 134 1088 138 1092
rect 414 1088 418 1092
rect 846 1088 850 1092
rect 1238 1088 1242 1092
rect 1334 1088 1338 1092
rect 1494 1088 1498 1092
rect 1598 1088 1602 1092
rect 1654 1088 1658 1092
rect 1798 1088 1802 1092
rect 1918 1088 1922 1092
rect 2046 1088 2050 1092
rect 2078 1088 2082 1092
rect 2230 1088 2234 1092
rect 2286 1088 2290 1092
rect 2430 1088 2434 1092
rect 2646 1088 2650 1092
rect 78 1078 82 1082
rect 110 1078 114 1082
rect 198 1078 202 1082
rect 214 1078 218 1082
rect 302 1078 306 1082
rect 334 1078 338 1082
rect 422 1078 426 1082
rect 446 1078 450 1082
rect 510 1078 514 1082
rect 526 1078 530 1082
rect 582 1078 586 1082
rect 638 1078 642 1082
rect 774 1078 778 1082
rect 838 1078 842 1082
rect 934 1078 938 1082
rect 958 1078 962 1082
rect 990 1078 994 1082
rect 998 1078 1002 1082
rect 1182 1078 1186 1082
rect 1190 1078 1194 1082
rect 1446 1078 1450 1082
rect 1550 1078 1554 1082
rect 1622 1078 1626 1082
rect 1630 1078 1634 1082
rect 1638 1078 1642 1082
rect 1790 1078 1794 1082
rect 1910 1078 1914 1082
rect 2086 1078 2090 1082
rect 2182 1078 2186 1082
rect 2214 1078 2218 1082
rect 2222 1078 2226 1082
rect 2302 1078 2306 1082
rect 2326 1078 2330 1082
rect 2350 1078 2354 1082
rect 2390 1078 2394 1082
rect 6 1068 10 1072
rect 38 1068 42 1072
rect 54 1068 58 1072
rect 94 1068 98 1072
rect 118 1068 122 1072
rect 134 1068 138 1072
rect 198 1068 202 1072
rect 214 1068 218 1072
rect 350 1068 354 1072
rect 454 1068 458 1072
rect 542 1068 546 1072
rect 558 1068 562 1072
rect 598 1068 602 1072
rect 774 1068 778 1072
rect 830 1068 834 1072
rect 894 1068 898 1072
rect 902 1068 906 1072
rect 1006 1068 1010 1072
rect 1030 1068 1034 1072
rect 1062 1068 1066 1072
rect 1110 1068 1114 1072
rect 1158 1068 1162 1072
rect 1230 1068 1234 1072
rect 1270 1068 1274 1072
rect 1294 1068 1298 1072
rect 1502 1068 1506 1072
rect 14 1058 18 1062
rect 86 1058 90 1062
rect 230 1058 234 1062
rect 302 1059 306 1063
rect 366 1058 370 1062
rect 406 1058 410 1062
rect 478 1058 482 1062
rect 486 1058 490 1062
rect 550 1058 554 1062
rect 614 1058 618 1062
rect 662 1058 666 1062
rect 710 1058 714 1062
rect 742 1059 746 1063
rect 1534 1066 1538 1070
rect 1550 1068 1554 1072
rect 1558 1068 1562 1072
rect 1678 1068 1682 1072
rect 1742 1068 1746 1072
rect 1806 1068 1810 1072
rect 1822 1068 1826 1072
rect 1854 1068 1858 1072
rect 1902 1068 1906 1072
rect 1926 1068 1930 1072
rect 1942 1068 1946 1072
rect 1974 1068 1978 1072
rect 2022 1068 2026 1072
rect 2030 1068 2034 1072
rect 2054 1068 2058 1072
rect 2102 1068 2106 1072
rect 2142 1068 2146 1072
rect 2158 1068 2162 1072
rect 2254 1068 2258 1072
rect 2262 1068 2266 1072
rect 2486 1078 2490 1082
rect 2414 1068 2418 1072
rect 2462 1068 2466 1072
rect 2686 1078 2690 1082
rect 2510 1068 2514 1072
rect 2526 1068 2530 1072
rect 2558 1068 2562 1072
rect 2606 1068 2610 1072
rect 2622 1068 2626 1072
rect 2638 1068 2642 1072
rect 798 1058 802 1062
rect 822 1058 826 1062
rect 862 1058 866 1062
rect 894 1058 898 1062
rect 958 1058 962 1062
rect 974 1058 978 1062
rect 1078 1058 1082 1062
rect 1110 1058 1114 1062
rect 1150 1058 1154 1062
rect 1222 1058 1226 1062
rect 1302 1059 1306 1063
rect 1366 1058 1370 1062
rect 1398 1059 1402 1063
rect 1430 1058 1434 1062
rect 1446 1058 1450 1062
rect 1486 1058 1490 1062
rect 1582 1058 1586 1062
rect 1638 1058 1642 1062
rect 1662 1058 1666 1062
rect 1686 1058 1690 1062
rect 1702 1058 1706 1062
rect 1718 1058 1722 1062
rect 1774 1058 1778 1062
rect 1814 1058 1818 1062
rect 1830 1058 1834 1062
rect 1934 1058 1938 1062
rect 1950 1058 1954 1062
rect 2094 1058 2098 1062
rect 2110 1058 2114 1062
rect 2150 1058 2154 1062
rect 2166 1058 2170 1062
rect 2174 1058 2178 1062
rect 2198 1058 2202 1062
rect 2254 1058 2258 1062
rect 2270 1058 2274 1062
rect 2318 1058 2322 1062
rect 2342 1058 2346 1062
rect 2366 1058 2370 1062
rect 2470 1058 2474 1062
rect 2518 1058 2522 1062
rect 2550 1058 2554 1062
rect 2630 1058 2634 1062
rect 2662 1058 2666 1062
rect 30 1048 34 1052
rect 54 1048 58 1052
rect 134 1048 138 1052
rect 158 1048 162 1052
rect 502 1048 506 1052
rect 534 1048 538 1052
rect 870 1048 874 1052
rect 902 1048 906 1052
rect 966 1048 970 1052
rect 1054 1048 1058 1052
rect 1086 1048 1090 1052
rect 1206 1048 1210 1052
rect 1670 1048 1674 1052
rect 1710 1048 1714 1052
rect 1782 1048 1786 1052
rect 1830 1048 1834 1052
rect 1950 1048 1954 1052
rect 2046 1048 2050 1052
rect 2078 1048 2082 1052
rect 2118 1048 2122 1052
rect 2230 1048 2234 1052
rect 2334 1048 2338 1052
rect 2478 1048 2482 1052
rect 2550 1048 2554 1052
rect 2614 1048 2618 1052
rect 2646 1048 2650 1052
rect 238 1038 242 1042
rect 654 1038 658 1042
rect 678 1038 682 1042
rect 806 1038 810 1042
rect 950 1038 954 1042
rect 1070 1038 1074 1042
rect 1118 1038 1122 1042
rect 1654 1038 1658 1042
rect 1726 1038 1730 1042
rect 1750 1038 1754 1042
rect 1766 1038 1770 1042
rect 1886 1038 1890 1042
rect 2006 1038 2010 1042
rect 2494 1038 2498 1042
rect 230 1018 234 1022
rect 470 1018 474 1022
rect 574 1018 578 1022
rect 638 1018 642 1022
rect 662 1018 666 1022
rect 982 1018 986 1022
rect 1038 1018 1042 1022
rect 1662 1018 1666 1022
rect 1718 1018 1722 1022
rect 1774 1018 1778 1022
rect 2358 1018 2362 1022
rect 2406 1018 2410 1022
rect 2574 1018 2578 1022
rect 578 1003 582 1007
rect 585 1003 589 1007
rect 1602 1003 1606 1007
rect 1609 1003 1613 1007
rect 126 988 130 992
rect 238 988 242 992
rect 454 988 458 992
rect 798 988 802 992
rect 846 988 850 992
rect 1246 988 1250 992
rect 1278 988 1282 992
rect 1446 988 1450 992
rect 1630 988 1634 992
rect 1998 988 2002 992
rect 2222 988 2226 992
rect 2254 988 2258 992
rect 2518 988 2522 992
rect 726 978 730 982
rect 406 968 410 972
rect 734 968 738 972
rect 806 968 810 972
rect 838 968 842 972
rect 870 968 874 972
rect 1294 968 1298 972
rect 1614 968 1618 972
rect 1830 968 1834 972
rect 2638 968 2642 972
rect 6 958 10 962
rect 118 958 122 962
rect 254 958 258 962
rect 262 958 266 962
rect 366 958 370 962
rect 526 958 530 962
rect 774 958 778 962
rect 958 958 962 962
rect 1222 958 1226 962
rect 1406 958 1410 962
rect 1462 958 1466 962
rect 1686 958 1690 962
rect 1854 958 1858 962
rect 1870 958 1874 962
rect 2038 958 2042 962
rect 2086 958 2090 962
rect 30 948 34 952
rect 46 948 50 952
rect 94 948 98 952
rect 110 948 114 952
rect 150 948 154 952
rect 238 948 242 952
rect 286 948 290 952
rect 430 948 434 952
rect 494 948 498 952
rect 502 948 506 952
rect 542 948 546 952
rect 614 948 618 952
rect 646 947 650 951
rect 678 948 682 952
rect 726 948 730 952
rect 814 948 818 952
rect 822 948 826 952
rect 846 948 850 952
rect 862 948 866 952
rect 886 948 890 952
rect 918 948 922 952
rect 950 948 954 952
rect 974 948 978 952
rect 1062 947 1066 951
rect 1094 948 1098 952
rect 1174 947 1178 951
rect 1206 948 1210 952
rect 1342 947 1346 951
rect 1374 948 1378 952
rect 1422 948 1426 952
rect 1430 948 1434 952
rect 1574 948 1578 952
rect 1646 948 1650 952
rect 1678 948 1682 952
rect 1710 948 1714 952
rect 1774 948 1778 952
rect 1870 948 1874 952
rect 1950 948 1954 952
rect 1966 948 1970 952
rect 2054 948 2058 952
rect 2094 948 2098 952
rect 2278 958 2282 962
rect 2310 958 2314 962
rect 2398 958 2402 962
rect 2214 948 2218 952
rect 2238 948 2242 952
rect 2326 948 2330 952
rect 2438 948 2442 952
rect 2486 948 2490 952
rect 2494 948 2498 952
rect 2502 948 2506 952
rect 2534 948 2538 952
rect 2558 948 2562 952
rect 2622 948 2626 952
rect 102 938 106 942
rect 134 938 138 942
rect 174 938 178 942
rect 222 938 226 942
rect 230 938 234 942
rect 294 938 298 942
rect 374 938 378 942
rect 422 938 426 942
rect 486 938 490 942
rect 606 938 610 942
rect 790 938 794 942
rect 894 938 898 942
rect 966 938 970 942
rect 982 938 986 942
rect 990 938 994 942
rect 1006 938 1010 942
rect 1014 938 1018 942
rect 1046 938 1050 942
rect 1142 938 1146 942
rect 1358 938 1362 942
rect 1382 938 1386 942
rect 1430 938 1434 942
rect 1438 938 1442 942
rect 1470 938 1474 942
rect 1550 938 1554 942
rect 1702 938 1706 942
rect 1718 938 1722 942
rect 1750 938 1754 942
rect 1838 938 1842 942
rect 1862 938 1866 942
rect 2022 938 2026 942
rect 2062 938 2066 942
rect 2070 938 2074 942
rect 2150 938 2154 942
rect 2158 938 2162 942
rect 2206 938 2210 942
rect 2302 938 2306 942
rect 2326 938 2330 942
rect 2358 938 2362 942
rect 2382 938 2386 942
rect 2414 938 2418 942
rect 2670 938 2674 942
rect 6 928 10 932
rect 62 928 66 932
rect 318 928 322 932
rect 350 928 354 932
rect 358 928 362 932
rect 430 928 434 932
rect 446 928 450 932
rect 462 928 466 932
rect 470 928 474 932
rect 502 928 506 932
rect 558 928 562 932
rect 590 928 594 932
rect 750 928 754 932
rect 934 928 938 932
rect 990 928 994 932
rect 1030 928 1034 932
rect 1262 928 1266 932
rect 1654 928 1658 932
rect 1734 928 1738 932
rect 1902 928 1906 932
rect 2006 928 2010 932
rect 2110 928 2114 932
rect 2126 928 2130 932
rect 2230 928 2234 932
rect 2390 928 2394 932
rect 2422 928 2426 932
rect 2462 928 2466 932
rect 2470 928 2474 932
rect 2542 928 2546 932
rect 2702 928 2706 932
rect 30 918 34 922
rect 46 918 50 922
rect 166 918 170 922
rect 206 918 210 922
rect 270 918 274 922
rect 302 918 306 922
rect 478 918 482 922
rect 574 918 578 922
rect 598 918 602 922
rect 758 918 762 922
rect 1134 918 1138 922
rect 1238 918 1242 922
rect 1270 918 1274 922
rect 1278 918 1282 922
rect 1390 918 1394 922
rect 1526 918 1530 922
rect 1646 918 1650 922
rect 1726 918 1730 922
rect 1854 918 1858 922
rect 2014 918 2018 922
rect 2086 918 2090 922
rect 2174 918 2178 922
rect 2270 918 2274 922
rect 2318 918 2322 922
rect 2366 918 2370 922
rect 2406 918 2410 922
rect 2430 918 2434 922
rect 2454 918 2458 922
rect 2478 918 2482 922
rect 2582 918 2586 922
rect 2686 918 2690 922
rect 286 908 290 912
rect 318 908 322 912
rect 1082 903 1086 907
rect 1089 903 1093 907
rect 2106 903 2110 907
rect 2113 903 2117 907
rect 102 898 106 902
rect 78 888 82 892
rect 142 888 146 892
rect 182 888 186 892
rect 246 888 250 892
rect 294 888 298 892
rect 366 888 370 892
rect 382 888 386 892
rect 486 888 490 892
rect 606 888 610 892
rect 878 888 882 892
rect 886 888 890 892
rect 1054 888 1058 892
rect 1110 888 1114 892
rect 1182 888 1186 892
rect 1206 888 1210 892
rect 1454 888 1458 892
rect 1462 888 1466 892
rect 1574 888 1578 892
rect 1694 888 1698 892
rect 1814 888 1818 892
rect 1822 888 1826 892
rect 1862 888 1866 892
rect 1894 888 1898 892
rect 1982 888 1986 892
rect 2398 888 2402 892
rect 2598 888 2602 892
rect 2654 888 2658 892
rect 102 878 106 882
rect 190 878 194 882
rect 494 878 498 882
rect 558 878 562 882
rect 574 878 578 882
rect 766 878 770 882
rect 1086 878 1090 882
rect 1166 878 1170 882
rect 1302 878 1306 882
rect 1318 878 1322 882
rect 1526 878 1530 882
rect 1630 878 1634 882
rect 1662 878 1666 882
rect 1750 878 1754 882
rect 1830 878 1834 882
rect 1838 878 1842 882
rect 1886 878 1890 882
rect 1934 878 1938 882
rect 62 868 66 872
rect 102 868 106 872
rect 158 868 162 872
rect 214 868 218 872
rect 262 868 266 872
rect 270 868 274 872
rect 374 868 378 872
rect 462 868 466 872
rect 558 868 562 872
rect 582 868 586 872
rect 630 868 634 872
rect 750 868 754 872
rect 766 868 770 872
rect 966 868 970 872
rect 982 868 986 872
rect 1014 868 1018 872
rect 1078 868 1082 872
rect 1118 868 1122 872
rect 1150 868 1154 872
rect 2006 878 2010 882
rect 2070 878 2074 882
rect 2086 878 2090 882
rect 2190 878 2194 882
rect 2246 878 2250 882
rect 2294 878 2298 882
rect 2310 878 2314 882
rect 2374 878 2378 882
rect 2414 878 2418 882
rect 2510 878 2514 882
rect 1302 868 1306 872
rect 1342 868 1346 872
rect 1358 868 1362 872
rect 1558 868 1562 872
rect 1590 868 1594 872
rect 1606 868 1610 872
rect 1646 868 1650 872
rect 1718 868 1722 872
rect 1734 868 1738 872
rect 1878 868 1882 872
rect 1902 868 1906 872
rect 1974 868 1978 872
rect 2014 868 2018 872
rect 2062 868 2066 872
rect 2214 868 2218 872
rect 2222 868 2226 872
rect 2254 868 2258 872
rect 2270 868 2274 872
rect 2318 868 2322 872
rect 2366 868 2370 872
rect 2390 868 2394 872
rect 2406 868 2410 872
rect 2430 868 2434 872
rect 2534 868 2538 872
rect 2550 868 2554 872
rect 2582 868 2586 872
rect 2638 868 2642 872
rect 2686 868 2690 872
rect 30 858 34 862
rect 86 858 90 862
rect 206 858 210 862
rect 326 858 330 862
rect 446 859 450 863
rect 478 858 482 862
rect 518 858 522 862
rect 622 858 626 862
rect 654 858 658 862
rect 734 859 738 863
rect 782 858 786 862
rect 814 859 818 863
rect 846 858 850 862
rect 942 858 946 862
rect 982 858 986 862
rect 1014 858 1018 862
rect 1046 858 1050 862
rect 1126 858 1130 862
rect 1134 858 1138 862
rect 1142 858 1146 862
rect 1246 858 1250 862
rect 1270 859 1274 863
rect 1318 858 1322 862
rect 1358 858 1362 862
rect 1390 859 1394 863
rect 1414 858 1418 862
rect 1526 859 1530 863
rect 1598 858 1602 862
rect 1614 858 1618 862
rect 1654 858 1658 862
rect 1758 858 1762 862
rect 1854 858 1858 862
rect 1918 858 1922 862
rect 1958 858 1962 862
rect 1990 858 1994 862
rect 2006 858 2010 862
rect 2022 858 2026 862
rect 2030 858 2034 862
rect 2070 858 2074 862
rect 2094 858 2098 862
rect 2134 858 2138 862
rect 2174 858 2178 862
rect 2222 858 2226 862
rect 2230 858 2234 862
rect 2262 858 2266 862
rect 2350 858 2354 862
rect 2454 858 2458 862
rect 2526 858 2530 862
rect 2558 858 2562 862
rect 2574 858 2578 862
rect 6 848 10 852
rect 22 848 26 852
rect 166 848 170 852
rect 566 848 570 852
rect 590 848 594 852
rect 510 838 514 842
rect 646 838 650 842
rect 1006 848 1010 852
rect 1582 848 1586 852
rect 1702 848 1706 852
rect 1966 848 1970 852
rect 1998 848 2002 852
rect 2038 848 2042 852
rect 2046 848 2050 852
rect 2150 848 2154 852
rect 2454 848 2458 852
rect 2486 848 2490 852
rect 2542 848 2546 852
rect 2574 848 2578 852
rect 1150 838 1154 842
rect 1950 838 1954 842
rect 2294 838 2298 842
rect 1958 828 1962 832
rect 174 818 178 822
rect 350 818 354 822
rect 518 818 522 822
rect 654 818 658 822
rect 1054 818 1058 822
rect 1814 818 1818 822
rect 2054 818 2058 822
rect 2174 818 2178 822
rect 2422 818 2426 822
rect 578 803 582 807
rect 585 803 589 807
rect 1602 803 1606 807
rect 1609 803 1613 807
rect 582 788 586 792
rect 774 788 778 792
rect 1174 788 1178 792
rect 1398 788 1402 792
rect 1422 788 1426 792
rect 1526 788 1530 792
rect 2198 788 2202 792
rect 2222 788 2226 792
rect 2318 788 2322 792
rect 2518 788 2522 792
rect 2622 788 2626 792
rect 86 778 90 782
rect 102 768 106 772
rect 566 768 570 772
rect 598 768 602 772
rect 1838 768 1842 772
rect 2238 768 2242 772
rect 2686 778 2690 782
rect 2294 768 2298 772
rect 2526 768 2530 772
rect 174 758 178 762
rect 214 758 218 762
rect 238 758 242 762
rect 270 758 274 762
rect 302 758 306 762
rect 310 758 314 762
rect 430 758 434 762
rect 446 758 450 762
rect 542 758 546 762
rect 550 758 554 762
rect 726 758 730 762
rect 758 758 762 762
rect 894 758 898 762
rect 902 758 906 762
rect 950 758 954 762
rect 1438 758 1442 762
rect 1774 758 1778 762
rect 1854 758 1858 762
rect 1886 758 1890 762
rect 1942 758 1946 762
rect 2014 758 2018 762
rect 2030 758 2034 762
rect 2278 758 2282 762
rect 22 748 26 752
rect 38 748 42 752
rect 54 748 58 752
rect 70 748 74 752
rect 86 748 90 752
rect 134 748 138 752
rect 166 748 170 752
rect 190 748 194 752
rect 254 748 258 752
rect 286 748 290 752
rect 350 748 354 752
rect 446 748 450 752
rect 54 738 58 742
rect 62 738 66 742
rect 158 738 162 742
rect 182 738 186 742
rect 222 738 226 742
rect 246 738 250 742
rect 278 738 282 742
rect 294 738 298 742
rect 358 738 362 742
rect 406 738 410 742
rect 414 738 418 742
rect 454 738 458 742
rect 494 748 498 752
rect 510 748 514 752
rect 542 748 546 752
rect 558 748 562 752
rect 470 738 474 742
rect 518 738 522 742
rect 662 747 666 751
rect 718 748 722 752
rect 742 748 746 752
rect 774 748 778 752
rect 854 747 858 751
rect 934 748 938 752
rect 958 748 962 752
rect 1006 748 1010 752
rect 1014 748 1018 752
rect 678 738 682 742
rect 694 738 698 742
rect 750 738 754 742
rect 782 738 786 742
rect 846 738 850 742
rect 1086 747 1090 751
rect 1118 748 1122 752
rect 1158 748 1162 752
rect 1214 747 1218 751
rect 1246 748 1250 752
rect 1350 747 1354 751
rect 1382 748 1386 752
rect 1406 748 1410 752
rect 1614 748 1618 752
rect 1710 748 1714 752
rect 1734 748 1738 752
rect 1822 748 1826 752
rect 1846 748 1850 752
rect 1862 748 1866 752
rect 1958 748 1962 752
rect 2006 748 2010 752
rect 2062 748 2066 752
rect 2078 748 2082 752
rect 2126 747 2130 751
rect 2254 748 2258 752
rect 2270 748 2274 752
rect 2286 748 2290 752
rect 2318 748 2322 752
rect 2342 758 2346 762
rect 2430 758 2434 762
rect 2550 758 2554 762
rect 2574 758 2578 762
rect 2606 758 2610 762
rect 2678 758 2682 762
rect 926 738 930 742
rect 958 738 962 742
rect 974 738 978 742
rect 1022 738 1026 742
rect 1182 738 1186 742
rect 1366 738 1370 742
rect 1446 738 1450 742
rect 1510 738 1514 742
rect 1582 738 1586 742
rect 1606 738 1610 742
rect 1638 738 1642 742
rect 1798 738 1802 742
rect 1814 738 1818 742
rect 1902 738 1906 742
rect 1918 738 1922 742
rect 1934 738 1938 742
rect 1990 738 1994 742
rect 2046 738 2050 742
rect 2070 738 2074 742
rect 2110 738 2114 742
rect 2238 738 2242 742
rect 2398 748 2402 752
rect 2406 748 2410 752
rect 2462 748 2466 752
rect 2534 748 2538 752
rect 2566 748 2570 752
rect 2590 748 2594 752
rect 2654 748 2658 752
rect 2310 738 2314 742
rect 2366 738 2370 742
rect 2390 738 2394 742
rect 2510 738 2514 742
rect 2566 738 2570 742
rect 2598 738 2602 742
rect 2630 738 2634 742
rect 2662 738 2666 742
rect 6 728 10 732
rect 110 728 114 732
rect 118 728 122 732
rect 150 728 154 732
rect 214 728 218 732
rect 334 728 338 732
rect 414 728 418 732
rect 510 728 514 732
rect 694 728 698 732
rect 974 728 978 732
rect 1038 728 1042 732
rect 1670 728 1674 732
rect 1782 728 1786 732
rect 1798 728 1802 732
rect 1846 728 1850 732
rect 1878 728 1882 732
rect 1910 728 1914 732
rect 1998 728 2002 732
rect 2022 728 2026 732
rect 2038 728 2042 732
rect 2054 728 2058 732
rect 2206 728 2210 732
rect 2238 728 2242 732
rect 2374 728 2378 732
rect 2406 728 2410 732
rect 2438 728 2442 732
rect 2638 728 2642 732
rect 2694 728 2698 732
rect 54 718 58 722
rect 86 718 90 722
rect 230 718 234 722
rect 310 718 314 722
rect 374 718 378 722
rect 398 718 402 722
rect 478 718 482 722
rect 790 718 794 722
rect 990 718 994 722
rect 1030 718 1034 722
rect 1150 718 1154 722
rect 1174 718 1178 722
rect 1278 718 1282 722
rect 1286 718 1290 722
rect 1398 718 1402 722
rect 1526 718 1530 722
rect 1630 718 1634 722
rect 1646 718 1650 722
rect 1766 718 1770 722
rect 1806 718 1810 722
rect 1870 718 1874 722
rect 1942 718 1946 722
rect 2190 718 2194 722
rect 2422 718 2426 722
rect 2478 718 2482 722
rect 2678 718 2682 722
rect 118 708 122 712
rect 214 708 218 712
rect 1082 703 1086 707
rect 1089 703 1093 707
rect 2106 703 2110 707
rect 2113 703 2117 707
rect 62 698 66 702
rect 70 698 74 702
rect 22 688 26 692
rect 102 688 106 692
rect 142 688 146 692
rect 174 688 178 692
rect 230 688 234 692
rect 278 688 282 692
rect 310 688 314 692
rect 374 688 378 692
rect 862 688 866 692
rect 958 688 962 692
rect 1198 688 1202 692
rect 1254 688 1258 692
rect 1358 688 1362 692
rect 1438 688 1442 692
rect 1958 688 1962 692
rect 2038 688 2042 692
rect 2198 688 2202 692
rect 2278 688 2282 692
rect 2294 688 2298 692
rect 2342 688 2346 692
rect 2590 688 2594 692
rect 2678 688 2682 692
rect 6 678 10 682
rect 62 678 66 682
rect 22 668 26 672
rect 46 668 50 672
rect 150 678 154 682
rect 182 678 186 682
rect 238 678 242 682
rect 246 678 250 682
rect 270 678 274 682
rect 334 678 338 682
rect 422 678 426 682
rect 470 678 474 682
rect 478 678 482 682
rect 526 678 530 682
rect 614 678 618 682
rect 718 678 722 682
rect 854 678 858 682
rect 1190 678 1194 682
rect 1446 678 1450 682
rect 1510 678 1514 682
rect 1662 678 1666 682
rect 1742 678 1746 682
rect 1750 678 1754 682
rect 1838 678 1842 682
rect 1862 678 1866 682
rect 2006 679 2010 683
rect 2054 678 2058 682
rect 2086 678 2090 682
rect 2142 678 2146 682
rect 2206 678 2210 682
rect 2326 678 2330 682
rect 2430 678 2434 682
rect 2438 678 2442 682
rect 2454 678 2458 682
rect 2478 678 2482 682
rect 2518 678 2522 682
rect 2566 678 2570 682
rect 86 668 90 672
rect 126 668 130 672
rect 166 668 170 672
rect 190 668 194 672
rect 214 668 218 672
rect 222 668 226 672
rect 286 668 290 672
rect 358 668 362 672
rect 366 668 370 672
rect 398 668 402 672
rect 454 668 458 672
rect 606 668 610 672
rect 670 668 674 672
rect 734 668 738 672
rect 846 668 850 672
rect 870 668 874 672
rect 902 668 906 672
rect 982 668 986 672
rect 1206 668 1210 672
rect 1246 668 1250 672
rect 1278 668 1282 672
rect 1342 668 1346 672
rect 1350 668 1354 672
rect 1398 668 1402 672
rect 1414 668 1418 672
rect 1422 668 1426 672
rect 1454 668 1458 672
rect 1510 668 1514 672
rect 1614 668 1618 672
rect 1622 668 1626 672
rect 1750 668 1754 672
rect 1766 668 1770 672
rect 1782 668 1786 672
rect 1854 668 1858 672
rect 1870 668 1874 672
rect 1942 668 1946 672
rect 1990 668 1994 672
rect 2022 668 2026 672
rect 2062 668 2066 672
rect 2182 668 2186 672
rect 2222 668 2226 672
rect 2238 668 2242 672
rect 2270 668 2274 672
rect 2326 668 2330 672
rect 2366 668 2370 672
rect 2374 668 2378 672
rect 2414 668 2418 672
rect 2526 668 2530 672
rect 2542 668 2546 672
rect 2574 668 2578 672
rect 2622 668 2626 672
rect 22 658 26 662
rect 38 658 42 662
rect 78 658 82 662
rect 94 658 98 662
rect 118 658 122 662
rect 126 658 130 662
rect 158 658 162 662
rect 206 658 210 662
rect 246 658 250 662
rect 262 658 266 662
rect 294 658 298 662
rect 342 658 346 662
rect 374 658 378 662
rect 390 658 394 662
rect 422 658 426 662
rect 454 658 458 662
rect 494 658 498 662
rect 534 658 538 662
rect 558 658 562 662
rect 630 658 634 662
rect 646 658 650 662
rect 678 658 682 662
rect 750 659 754 663
rect 782 658 786 662
rect 838 658 842 662
rect 878 658 882 662
rect 894 658 898 662
rect 942 658 946 662
rect 974 658 978 662
rect 1006 658 1010 662
rect 1014 658 1018 662
rect 1046 658 1050 662
rect 1070 658 1074 662
rect 1078 658 1082 662
rect 1118 658 1122 662
rect 1126 658 1130 662
rect 1150 658 1154 662
rect 1166 658 1170 662
rect 1182 658 1186 662
rect 1214 658 1218 662
rect 1238 658 1242 662
rect 1270 658 1274 662
rect 1278 658 1282 662
rect 1318 658 1322 662
rect 1406 658 1410 662
rect 1422 658 1426 662
rect 1462 658 1466 662
rect 1486 658 1490 662
rect 1550 658 1554 662
rect 1558 658 1562 662
rect 1694 658 1698 662
rect 1726 658 1730 662
rect 1782 658 1786 662
rect 1798 658 1802 662
rect 1854 658 1858 662
rect 1894 658 1898 662
rect 1902 658 1906 662
rect 1926 658 1930 662
rect 1934 658 1938 662
rect 2014 658 2018 662
rect 2102 658 2106 662
rect 2126 658 2130 662
rect 2142 658 2146 662
rect 2166 658 2170 662
rect 2214 658 2218 662
rect 2238 658 2242 662
rect 2246 658 2250 662
rect 2310 658 2314 662
rect 2358 658 2362 662
rect 2382 658 2386 662
rect 2478 658 2482 662
rect 2502 658 2506 662
rect 2510 658 2514 662
rect 2518 658 2522 662
rect 2630 658 2634 662
rect 2662 658 2666 662
rect 38 648 42 652
rect 102 648 106 652
rect 190 648 194 652
rect 318 648 322 652
rect 438 648 442 652
rect 638 648 642 652
rect 694 648 698 652
rect 822 648 826 652
rect 838 648 842 652
rect 886 648 890 652
rect 1254 648 1258 652
rect 1390 648 1394 652
rect 1766 648 1770 652
rect 2182 648 2186 652
rect 2198 648 2202 652
rect 2246 648 2250 652
rect 2270 648 2274 652
rect 2286 648 2290 652
rect 2294 648 2298 652
rect 2398 648 2402 652
rect 358 638 362 642
rect 430 638 434 642
rect 590 638 594 642
rect 654 638 658 642
rect 814 638 818 642
rect 902 638 906 642
rect 926 638 930 642
rect 1142 638 1146 642
rect 1174 638 1178 642
rect 1222 638 1226 642
rect 1478 638 1482 642
rect 1518 638 1522 642
rect 2110 638 2114 642
rect 2158 638 2162 642
rect 2486 638 2490 642
rect 710 628 714 632
rect 1054 628 1058 632
rect 2446 628 2450 632
rect 494 618 498 622
rect 662 618 666 622
rect 1238 618 1242 622
rect 1302 618 1306 622
rect 1638 618 1642 622
rect 1678 618 1682 622
rect 1718 618 1722 622
rect 1806 618 1810 622
rect 1910 618 1914 622
rect 2166 618 2170 622
rect 2430 618 2434 622
rect 578 603 582 607
rect 585 603 589 607
rect 1602 603 1606 607
rect 1609 603 1613 607
rect 86 588 90 592
rect 190 588 194 592
rect 262 588 266 592
rect 430 588 434 592
rect 718 588 722 592
rect 1094 588 1098 592
rect 1446 588 1450 592
rect 1486 588 1490 592
rect 1774 588 1778 592
rect 1926 588 1930 592
rect 1934 588 1938 592
rect 2278 588 2282 592
rect 2294 588 2298 592
rect 2334 588 2338 592
rect 2342 588 2346 592
rect 806 568 810 572
rect 846 568 850 572
rect 1230 568 1234 572
rect 1270 568 1274 572
rect 1438 568 1442 572
rect 1454 568 1458 572
rect 2182 568 2186 572
rect 38 558 42 562
rect 118 558 122 562
rect 222 558 226 562
rect 302 558 306 562
rect 526 558 530 562
rect 702 558 706 562
rect 118 548 122 552
rect 126 548 130 552
rect 134 548 138 552
rect 182 548 186 552
rect 310 548 314 552
rect 318 548 322 552
rect 374 548 378 552
rect 406 548 410 552
rect 494 547 498 551
rect 638 547 642 551
rect 670 548 674 552
rect 694 548 698 552
rect 718 548 722 552
rect 1038 558 1042 562
rect 1310 558 1314 562
rect 1470 558 1474 562
rect 1478 558 1482 562
rect 1590 558 1594 562
rect 1726 558 1730 562
rect 1798 558 1802 562
rect 2454 558 2458 562
rect 2614 558 2618 562
rect 2630 558 2634 562
rect 742 548 746 552
rect 750 548 754 552
rect 766 548 770 552
rect 798 548 802 552
rect 814 548 818 552
rect 822 548 826 552
rect 894 547 898 551
rect 950 548 954 552
rect 982 548 986 552
rect 998 548 1002 552
rect 1086 548 1090 552
rect 1158 547 1162 551
rect 1198 548 1202 552
rect 1214 548 1218 552
rect 1222 548 1226 552
rect 1230 548 1234 552
rect 1270 548 1274 552
rect 1318 548 1322 552
rect 6 538 10 542
rect 54 538 58 542
rect 142 538 146 542
rect 166 538 170 542
rect 206 538 210 542
rect 238 538 242 542
rect 246 538 250 542
rect 294 538 298 542
rect 326 538 330 542
rect 366 538 370 542
rect 382 538 386 542
rect 510 538 514 542
rect 542 538 546 542
rect 622 538 626 542
rect 686 538 690 542
rect 726 538 730 542
rect 758 538 762 542
rect 766 538 770 542
rect 910 538 914 542
rect 990 538 994 542
rect 1022 538 1026 542
rect 1102 538 1106 542
rect 1126 538 1130 542
rect 1174 538 1178 542
rect 1206 538 1210 542
rect 1238 538 1242 542
rect 1254 538 1258 542
rect 1374 547 1378 551
rect 1406 548 1410 552
rect 1462 548 1466 552
rect 1486 548 1490 552
rect 1526 548 1530 552
rect 1534 548 1538 552
rect 1574 548 1578 552
rect 1638 547 1642 551
rect 1758 548 1762 552
rect 1830 548 1834 552
rect 1862 547 1866 551
rect 1894 548 1898 552
rect 1982 548 1986 552
rect 2006 548 2010 552
rect 2070 548 2074 552
rect 2118 547 2122 551
rect 2214 547 2218 551
rect 2318 548 2322 552
rect 2406 547 2410 551
rect 2462 548 2466 552
rect 2550 548 2554 552
rect 2598 548 2602 552
rect 2614 548 2618 552
rect 2694 548 2698 552
rect 1286 538 1290 542
rect 1318 538 1322 542
rect 1326 538 1330 542
rect 1342 538 1346 542
rect 1542 538 1546 542
rect 1566 538 1570 542
rect 1582 538 1586 542
rect 1622 538 1626 542
rect 1710 538 1714 542
rect 1726 538 1730 542
rect 1750 538 1754 542
rect 1782 538 1786 542
rect 1798 538 1802 542
rect 1822 538 1826 542
rect 1830 538 1834 542
rect 2046 538 2050 542
rect 2062 538 2066 542
rect 2102 538 2106 542
rect 2222 538 2226 542
rect 2286 538 2290 542
rect 2422 538 2426 542
rect 2454 538 2458 542
rect 2494 538 2498 542
rect 2590 538 2594 542
rect 2606 538 2610 542
rect 2670 538 2674 542
rect 62 528 66 532
rect 94 528 98 532
rect 102 528 106 532
rect 150 528 154 532
rect 166 528 170 532
rect 334 528 338 532
rect 358 528 362 532
rect 422 528 426 532
rect 550 528 554 532
rect 670 528 674 532
rect 790 528 794 532
rect 934 528 938 532
rect 1190 528 1194 532
rect 1270 528 1274 532
rect 1342 528 1346 532
rect 1518 527 1522 531
rect 1558 528 1562 532
rect 1734 528 1738 532
rect 1766 528 1770 532
rect 1806 528 1810 532
rect 2046 528 2050 532
rect 2054 528 2058 532
rect 2302 528 2306 532
rect 2438 528 2442 532
rect 2502 528 2506 532
rect 2566 528 2570 532
rect 2574 528 2578 532
rect 2582 528 2586 532
rect 2638 528 2642 532
rect 2678 528 2682 532
rect 46 518 50 522
rect 238 518 242 522
rect 390 518 394 522
rect 574 518 578 522
rect 782 518 786 522
rect 830 518 834 522
rect 966 518 970 522
rect 1014 518 1018 522
rect 1038 518 1042 522
rect 1054 518 1058 522
rect 1550 518 1554 522
rect 1702 518 1706 522
rect 1742 518 1746 522
rect 1814 518 1818 522
rect 2502 518 2506 522
rect 2558 518 2562 522
rect 78 508 82 512
rect 94 508 98 512
rect 166 508 170 512
rect 422 508 426 512
rect 1082 503 1086 507
rect 1089 503 1093 507
rect 2106 503 2110 507
rect 2113 503 2117 507
rect 14 488 18 492
rect 38 488 42 492
rect 134 488 138 492
rect 142 488 146 492
rect 158 488 162 492
rect 214 488 218 492
rect 222 488 226 492
rect 254 488 258 492
rect 390 488 394 492
rect 398 488 402 492
rect 422 488 426 492
rect 430 488 434 492
rect 662 488 666 492
rect 694 488 698 492
rect 734 488 738 492
rect 766 488 770 492
rect 886 488 890 492
rect 942 488 946 492
rect 1598 488 1602 492
rect 1662 488 1666 492
rect 1766 488 1770 492
rect 1774 488 1778 492
rect 1990 488 1994 492
rect 1998 488 2002 492
rect 2190 488 2194 492
rect 2286 488 2290 492
rect 2294 488 2298 492
rect 2390 488 2394 492
rect 2494 488 2498 492
rect 2510 488 2514 492
rect 2518 488 2522 492
rect 2566 488 2570 492
rect 2590 488 2594 492
rect 2686 488 2690 492
rect 86 478 90 482
rect 150 478 154 482
rect 238 478 242 482
rect 278 478 282 482
rect 310 478 314 482
rect 382 478 386 482
rect 6 468 10 472
rect 54 468 58 472
rect 62 468 66 472
rect 102 468 106 472
rect 174 468 178 472
rect 182 468 186 472
rect 230 468 234 472
rect 270 468 274 472
rect 318 468 322 472
rect 366 468 370 472
rect 390 468 394 472
rect 406 468 410 472
rect 550 478 554 482
rect 574 478 578 482
rect 606 478 610 482
rect 686 478 690 482
rect 718 478 722 482
rect 726 478 730 482
rect 950 478 954 482
rect 982 478 986 482
rect 1078 478 1082 482
rect 510 468 514 472
rect 542 468 546 472
rect 622 468 626 472
rect 662 468 666 472
rect 702 468 706 472
rect 790 468 794 472
rect 902 468 906 472
rect 918 468 922 472
rect 926 468 930 472
rect 966 468 970 472
rect 982 468 986 472
rect 1014 468 1018 472
rect 1174 468 1178 472
rect 1214 468 1218 472
rect 1230 468 1234 472
rect 1278 478 1282 482
rect 1438 478 1442 482
rect 1470 478 1474 482
rect 1654 478 1658 482
rect 1758 478 1762 482
rect 2222 478 2226 482
rect 2574 478 2578 482
rect 2702 478 2706 482
rect 1294 468 1298 472
rect 1310 468 1314 472
rect 62 458 66 462
rect 94 458 98 462
rect 134 458 138 462
rect 270 458 274 462
rect 494 459 498 463
rect 526 458 530 462
rect 558 458 562 462
rect 654 458 658 462
rect 702 458 706 462
rect 742 458 746 462
rect 758 458 762 462
rect 782 458 786 462
rect 822 459 826 463
rect 846 458 850 462
rect 910 458 914 462
rect 926 458 930 462
rect 958 458 962 462
rect 1030 458 1034 462
rect 1054 458 1058 462
rect 1118 458 1122 462
rect 1198 459 1202 463
rect 1830 468 1834 472
rect 1870 468 1874 472
rect 2046 468 2050 472
rect 2094 468 2098 472
rect 2486 468 2490 472
rect 2542 468 2546 472
rect 2558 468 2562 472
rect 1270 458 1274 462
rect 1302 458 1306 462
rect 1318 458 1322 462
rect 1334 458 1338 462
rect 1406 458 1410 462
rect 1438 459 1442 463
rect 1550 458 1554 462
rect 1558 458 1562 462
rect 1694 458 1698 462
rect 1726 459 1730 463
rect 1814 458 1818 462
rect 1878 458 1882 462
rect 1894 458 1898 462
rect 1926 459 1930 463
rect 1958 458 1962 462
rect 2014 458 2018 462
rect 2022 458 2026 462
rect 2038 458 2042 462
rect 2062 458 2066 462
rect 2126 459 2130 463
rect 2158 458 2162 462
rect 2222 459 2226 463
rect 2254 458 2258 462
rect 2326 458 2330 462
rect 2358 459 2362 463
rect 2422 458 2426 462
rect 2454 459 2458 463
rect 2494 458 2498 462
rect 2534 458 2538 462
rect 2550 458 2554 462
rect 2614 458 2618 462
rect 2646 459 2650 463
rect 78 448 82 452
rect 158 448 162 452
rect 894 448 898 452
rect 1094 448 1098 452
rect 766 438 770 442
rect 990 438 994 442
rect 1046 438 1050 442
rect 1110 438 1114 442
rect 1246 448 1250 452
rect 1582 448 1586 452
rect 2510 448 2514 452
rect 2518 448 2522 452
rect 2678 448 2682 452
rect 1350 438 1354 442
rect 334 418 338 422
rect 374 418 378 422
rect 982 418 986 422
rect 1094 418 1098 422
rect 1638 418 1642 422
rect 2294 418 2298 422
rect 2582 418 2586 422
rect 578 403 582 407
rect 585 403 589 407
rect 1602 403 1606 407
rect 1609 403 1613 407
rect 198 388 202 392
rect 318 388 322 392
rect 462 388 466 392
rect 630 388 634 392
rect 694 388 698 392
rect 838 388 842 392
rect 870 388 874 392
rect 1158 388 1162 392
rect 1246 388 1250 392
rect 1742 388 1746 392
rect 2182 388 2186 392
rect 2214 388 2218 392
rect 2310 388 2314 392
rect 2646 388 2650 392
rect 38 368 42 372
rect 502 368 506 372
rect 622 368 626 372
rect 830 368 834 372
rect 862 368 866 372
rect 1238 368 1242 372
rect 1390 368 1394 372
rect 1878 368 1882 372
rect 2038 368 2042 372
rect 150 358 154 362
rect 182 358 186 362
rect 278 358 282 362
rect 334 358 338 362
rect 638 358 642 362
rect 662 358 666 362
rect 710 358 714 362
rect 1014 358 1018 362
rect 1062 358 1066 362
rect 1190 358 1194 362
rect 1238 358 1242 362
rect 1542 358 1546 362
rect 1566 358 1570 362
rect 1942 358 1946 362
rect 2318 358 2322 362
rect 2382 358 2386 362
rect 2558 358 2562 362
rect 2622 358 2626 362
rect 62 348 66 352
rect 118 348 122 352
rect 150 348 154 352
rect 198 348 202 352
rect 230 348 234 352
rect 238 348 242 352
rect 278 348 282 352
rect 302 348 306 352
rect 310 348 314 352
rect 446 348 450 352
rect 494 348 498 352
rect 534 348 538 352
rect 6 338 10 342
rect 54 338 58 342
rect 118 338 122 342
rect 134 338 138 342
rect 150 338 154 342
rect 158 338 162 342
rect 206 338 210 342
rect 254 338 258 342
rect 566 347 570 351
rect 630 348 634 352
rect 694 348 698 352
rect 358 338 362 342
rect 406 338 410 342
rect 454 338 458 342
rect 470 338 474 342
rect 782 347 786 351
rect 814 348 818 352
rect 822 348 826 352
rect 846 348 850 352
rect 854 348 858 352
rect 910 348 914 352
rect 974 348 978 352
rect 998 348 1002 352
rect 1030 348 1034 352
rect 1094 347 1098 351
rect 1126 348 1130 352
rect 1174 348 1178 352
rect 1198 348 1202 352
rect 1214 348 1218 352
rect 1230 348 1234 352
rect 1246 348 1250 352
rect 1294 347 1298 351
rect 1326 348 1330 352
rect 1374 348 1378 352
rect 1398 348 1402 352
rect 1454 347 1458 351
rect 1638 348 1642 352
rect 1670 347 1674 351
rect 1734 348 1738 352
rect 1758 348 1762 352
rect 1814 347 1818 351
rect 1886 348 1890 352
rect 1918 348 1922 352
rect 1974 347 1978 351
rect 2054 348 2058 352
rect 2078 348 2082 352
rect 2118 347 2122 351
rect 2198 348 2202 352
rect 2246 347 2250 351
rect 2334 348 2338 352
rect 2350 348 2354 352
rect 2398 348 2402 352
rect 2430 348 2434 352
rect 2462 348 2466 352
rect 2510 348 2514 352
rect 2542 348 2546 352
rect 2582 348 2586 352
rect 2606 348 2610 352
rect 2614 348 2618 352
rect 966 338 970 342
rect 982 338 986 342
rect 990 338 994 342
rect 1014 338 1018 342
rect 1022 338 1026 342
rect 1166 338 1170 342
rect 1198 338 1202 342
rect 1206 338 1210 342
rect 1222 338 1226 342
rect 1366 338 1370 342
rect 1414 338 1418 342
rect 1526 338 1530 342
rect 1686 338 1690 342
rect 1718 338 1722 342
rect 1774 338 1778 342
rect 1798 338 1802 342
rect 1894 338 1898 342
rect 1910 338 1914 342
rect 1934 338 1938 342
rect 1958 338 1962 342
rect 2046 338 2050 342
rect 2102 338 2106 342
rect 2190 338 2194 342
rect 2254 338 2258 342
rect 2326 338 2330 342
rect 2342 338 2346 342
rect 2358 338 2362 342
rect 2406 338 2410 342
rect 2454 338 2458 342
rect 2470 338 2474 342
rect 2486 338 2490 342
rect 2550 338 2554 342
rect 2590 338 2594 342
rect 2638 338 2642 342
rect 2662 338 2666 342
rect 118 328 122 332
rect 174 328 178 332
rect 214 328 218 332
rect 238 328 242 332
rect 286 328 290 332
rect 414 328 418 332
rect 782 328 786 332
rect 926 328 930 332
rect 950 328 954 332
rect 1422 328 1426 332
rect 1454 328 1458 332
rect 1582 328 1586 332
rect 1702 328 1706 332
rect 1750 328 1754 332
rect 1910 328 1914 332
rect 2006 328 2010 332
rect 2246 328 2250 332
rect 2414 328 2418 332
rect 2422 328 2426 332
rect 2438 328 2442 332
rect 2494 328 2498 332
rect 2638 328 2642 332
rect 2646 328 2650 332
rect 2678 328 2682 332
rect 94 318 98 322
rect 222 318 226 322
rect 230 318 234 322
rect 294 318 298 322
rect 366 318 370 322
rect 438 318 442 322
rect 678 318 682 322
rect 718 318 722 322
rect 918 318 922 322
rect 1062 318 1066 322
rect 1358 318 1362 322
rect 1518 318 1522 322
rect 1558 318 1562 322
rect 1574 318 1578 322
rect 1606 318 1610 322
rect 1902 318 1906 322
rect 2350 318 2354 322
rect 2366 318 2370 322
rect 2446 318 2450 322
rect 2486 318 2490 322
rect 2510 318 2514 322
rect 2566 318 2570 322
rect 118 308 122 312
rect 158 308 162 312
rect 2414 308 2418 312
rect 2494 308 2498 312
rect 1082 303 1086 307
rect 1089 303 1093 307
rect 2106 303 2110 307
rect 2113 303 2117 307
rect 38 298 42 302
rect 326 298 330 302
rect 2238 298 2242 302
rect 46 288 50 292
rect 86 288 90 292
rect 422 288 426 292
rect 822 288 826 292
rect 830 288 834 292
rect 990 288 994 292
rect 1022 288 1026 292
rect 1086 288 1090 292
rect 1214 288 1218 292
rect 1238 288 1242 292
rect 1286 288 1290 292
rect 1326 288 1330 292
rect 1414 288 1418 292
rect 1630 288 1634 292
rect 1678 288 1682 292
rect 1774 288 1778 292
rect 2054 288 2058 292
rect 2158 288 2162 292
rect 2206 288 2210 292
rect 2230 288 2234 292
rect 2326 288 2330 292
rect 2398 288 2402 292
rect 2422 288 2426 292
rect 2582 288 2586 292
rect 2598 288 2602 292
rect 2694 288 2698 292
rect 6 278 10 282
rect 38 278 42 282
rect 118 278 122 282
rect 46 268 50 272
rect 78 268 82 272
rect 118 268 122 272
rect 150 278 154 282
rect 166 278 170 282
rect 206 278 210 282
rect 222 278 226 282
rect 286 278 290 282
rect 326 278 330 282
rect 558 278 562 282
rect 726 278 730 282
rect 926 278 930 282
rect 998 278 1002 282
rect 1118 278 1122 282
rect 1222 278 1226 282
rect 1262 278 1266 282
rect 1278 278 1282 282
rect 1310 278 1314 282
rect 1318 278 1322 282
rect 1406 278 1410 282
rect 1534 278 1538 282
rect 1782 278 1786 282
rect 1814 278 1818 282
rect 2142 278 2146 282
rect 2238 278 2242 282
rect 2286 278 2290 282
rect 2318 278 2322 282
rect 2406 278 2410 282
rect 2550 278 2554 282
rect 2590 278 2594 282
rect 142 268 146 272
rect 182 268 186 272
rect 310 268 314 272
rect 542 268 546 272
rect 678 268 682 272
rect 966 268 970 272
rect 982 268 986 272
rect 1006 268 1010 272
rect 1038 268 1042 272
rect 1046 268 1050 272
rect 1102 268 1106 272
rect 1254 268 1258 272
rect 1310 268 1314 272
rect 1358 268 1362 272
rect 1390 268 1394 272
rect 1454 268 1458 272
rect 1494 268 1498 272
rect 1518 268 1522 272
rect 1534 268 1538 272
rect 1654 268 1658 272
rect 1694 268 1698 272
rect 1822 268 1826 272
rect 1918 268 1922 272
rect 1950 268 1954 272
rect 2006 268 2010 272
rect 2078 268 2082 272
rect 2086 268 2090 272
rect 2102 268 2106 272
rect 2166 268 2170 272
rect 2174 268 2178 272
rect 2190 268 2194 272
rect 2206 268 2210 272
rect 2214 268 2218 272
rect 2262 268 2266 272
rect 2302 268 2306 272
rect 2326 268 2330 272
rect 2342 268 2346 272
rect 2374 268 2378 272
rect 2390 268 2394 272
rect 2430 268 2434 272
rect 2438 268 2442 272
rect 2486 268 2490 272
rect 2502 268 2506 272
rect 2614 268 2618 272
rect 38 258 42 262
rect 102 258 106 262
rect 174 258 178 262
rect 254 258 258 262
rect 270 258 274 262
rect 294 258 298 262
rect 366 258 370 262
rect 390 258 394 262
rect 454 259 458 263
rect 486 258 490 262
rect 526 258 530 262
rect 606 259 610 263
rect 638 258 642 262
rect 686 258 690 262
rect 758 259 762 263
rect 782 258 786 262
rect 862 258 866 262
rect 894 259 898 263
rect 974 258 978 262
rect 1054 258 1058 262
rect 1078 258 1082 262
rect 1150 259 1154 263
rect 1182 258 1186 262
rect 1262 258 1266 262
rect 1278 258 1282 262
rect 1342 258 1346 262
rect 1358 258 1362 262
rect 1470 258 1474 262
rect 1510 258 1514 262
rect 1534 258 1538 262
rect 1566 259 1570 263
rect 1590 258 1594 262
rect 1662 258 1666 262
rect 1718 258 1722 262
rect 1926 258 1930 262
rect 2014 258 2018 262
rect 2038 258 2042 262
rect 2046 258 2050 262
rect 2070 258 2074 262
rect 2094 258 2098 262
rect 2190 258 2194 262
rect 2254 258 2258 262
rect 2270 258 2274 262
rect 2286 258 2290 262
rect 2366 258 2370 262
rect 2382 258 2386 262
rect 2486 258 2490 262
rect 2518 259 2522 263
rect 2638 258 2642 262
rect 62 248 66 252
rect 158 248 162 252
rect 206 248 210 252
rect 238 248 242 252
rect 702 248 706 252
rect 718 248 722 252
rect 934 248 938 252
rect 950 248 954 252
rect 1022 248 1026 252
rect 1070 248 1074 252
rect 1118 248 1122 252
rect 1366 248 1370 252
rect 1382 248 1386 252
rect 1678 248 1682 252
rect 2110 248 2114 252
rect 2126 248 2130 252
rect 2150 248 2154 252
rect 2286 248 2290 252
rect 2326 248 2330 252
rect 2350 248 2354 252
rect 2366 248 2370 252
rect 670 238 674 242
rect 1798 238 1802 242
rect 518 218 522 222
rect 1878 218 1882 222
rect 578 203 582 207
rect 585 203 589 207
rect 1602 203 1606 207
rect 1609 203 1613 207
rect 438 188 442 192
rect 654 188 658 192
rect 782 188 786 192
rect 854 188 858 192
rect 894 188 898 192
rect 918 188 922 192
rect 942 188 946 192
rect 1694 188 1698 192
rect 2150 188 2154 192
rect 2342 188 2346 192
rect 2462 188 2466 192
rect 2558 188 2562 192
rect 2574 188 2578 192
rect 542 168 546 172
rect 1734 168 1738 172
rect 2046 168 2050 172
rect 2182 168 2186 172
rect 2222 168 2226 172
rect 2286 168 2290 172
rect 2510 168 2514 172
rect 630 158 634 162
rect 638 158 642 162
rect 694 158 698 162
rect 710 158 714 162
rect 902 158 906 162
rect 958 158 962 162
rect 1094 158 1098 162
rect 1222 158 1226 162
rect 1366 158 1370 162
rect 1950 158 1954 162
rect 2134 158 2138 162
rect 2246 158 2250 162
rect 2310 158 2314 162
rect 2374 158 2378 162
rect 2430 158 2434 162
rect 2478 158 2482 162
rect 2526 158 2530 162
rect 22 148 26 152
rect 38 148 42 152
rect 102 148 106 152
rect 142 148 146 152
rect 238 148 242 152
rect 278 148 282 152
rect 334 148 338 152
rect 358 148 362 152
rect 398 148 402 152
rect 430 148 434 152
rect 590 148 594 152
rect 614 148 618 152
rect 630 148 634 152
rect 654 148 658 152
rect 670 148 674 152
rect 686 148 690 152
rect 710 148 714 152
rect 750 148 754 152
rect 846 148 850 152
rect 870 148 874 152
rect 918 148 922 152
rect 934 148 938 152
rect 1166 148 1170 152
rect 1182 148 1186 152
rect 126 138 130 142
rect 158 138 162 142
rect 262 138 266 142
rect 310 138 314 142
rect 414 138 418 142
rect 502 138 506 142
rect 558 138 562 142
rect 598 138 602 142
rect 662 138 666 142
rect 726 138 730 142
rect 838 138 842 142
rect 878 138 882 142
rect 950 138 954 142
rect 982 138 986 142
rect 1030 138 1034 142
rect 1054 138 1058 142
rect 1310 147 1314 151
rect 1374 148 1378 152
rect 1470 148 1474 152
rect 1574 148 1578 152
rect 1630 148 1634 152
rect 1726 148 1730 152
rect 1766 148 1770 152
rect 1798 147 1802 151
rect 1846 148 1850 152
rect 1862 148 1866 152
rect 1870 148 1874 152
rect 1934 148 1938 152
rect 1990 148 1994 152
rect 2054 148 2058 152
rect 2086 148 2090 152
rect 2094 148 2098 152
rect 2102 148 2106 152
rect 2150 148 2154 152
rect 2198 148 2202 152
rect 2222 148 2226 152
rect 2246 148 2250 152
rect 2286 148 2290 152
rect 2366 148 2370 152
rect 2390 148 2394 152
rect 2406 148 2410 152
rect 2462 148 2466 152
rect 2518 148 2522 152
rect 2598 148 2602 152
rect 2638 148 2642 152
rect 1118 138 1122 142
rect 1222 138 1226 142
rect 1302 138 1306 142
rect 1382 138 1386 142
rect 1430 138 1434 142
rect 1478 138 1482 142
rect 1550 138 1554 142
rect 1638 138 1642 142
rect 1814 138 1818 142
rect 1886 138 1890 142
rect 1894 138 1898 142
rect 1902 140 1906 144
rect 1982 138 1986 142
rect 2062 138 2066 142
rect 2102 138 2106 142
rect 2158 138 2162 142
rect 2166 138 2170 142
rect 2182 138 2186 142
rect 2190 138 2194 142
rect 2262 138 2266 142
rect 2294 138 2298 142
rect 2342 138 2346 142
rect 2406 138 2410 142
rect 2422 138 2426 142
rect 2454 138 2458 142
rect 2486 138 2490 142
rect 2494 138 2498 142
rect 2502 138 2506 142
rect 2590 138 2594 142
rect 2614 138 2618 142
rect 14 128 18 132
rect 198 128 202 132
rect 286 127 290 131
rect 430 128 434 132
rect 462 128 466 132
rect 470 128 474 132
rect 486 128 490 132
rect 502 128 506 132
rect 574 128 578 132
rect 670 128 674 132
rect 766 128 770 132
rect 862 128 866 132
rect 894 128 898 132
rect 950 128 954 132
rect 998 128 1002 132
rect 1006 128 1010 132
rect 1046 128 1050 132
rect 1126 128 1130 132
rect 1158 128 1162 132
rect 1166 128 1170 132
rect 1190 128 1194 132
rect 1238 128 1242 132
rect 1342 128 1346 132
rect 1438 128 1442 132
rect 1470 128 1474 132
rect 1582 128 1586 132
rect 1630 128 1634 132
rect 1830 128 1834 132
rect 1886 128 1890 132
rect 1966 128 1970 132
rect 2238 128 2242 132
rect 2270 128 2274 132
rect 2550 128 2554 132
rect 2566 128 2570 132
rect 2574 128 2578 132
rect 46 118 50 122
rect 390 118 394 122
rect 742 118 746 122
rect 1214 118 1218 122
rect 1246 118 1250 122
rect 1406 118 1410 122
rect 1534 118 1538 122
rect 1710 118 1714 122
rect 1870 118 1874 122
rect 1950 118 1954 122
rect 2150 118 2154 122
rect 2214 118 2218 122
rect 2414 118 2418 122
rect 2438 118 2442 122
rect 2494 118 2498 122
rect 2510 118 2514 122
rect 2598 118 2602 122
rect 2694 118 2698 122
rect 1886 108 1890 112
rect 2270 108 2274 112
rect 1082 103 1086 107
rect 1089 103 1093 107
rect 2106 103 2110 107
rect 2113 103 2117 107
rect 2406 98 2410 102
rect 2582 98 2586 102
rect 94 88 98 92
rect 342 88 346 92
rect 502 88 506 92
rect 614 88 618 92
rect 678 88 682 92
rect 822 88 826 92
rect 894 88 898 92
rect 926 88 930 92
rect 982 88 986 92
rect 1174 88 1178 92
rect 1230 88 1234 92
rect 1326 88 1330 92
rect 1414 88 1418 92
rect 1430 88 1434 92
rect 1582 88 1586 92
rect 1726 88 1730 92
rect 1846 88 1850 92
rect 2134 88 2138 92
rect 2142 88 2146 92
rect 2166 88 2170 92
rect 2174 88 2178 92
rect 2526 88 2530 92
rect 2550 88 2554 92
rect 2606 88 2610 92
rect 2614 88 2618 92
rect 2646 88 2650 92
rect 2694 88 2698 92
rect 54 78 58 82
rect 158 78 162 82
rect 278 78 282 82
rect 438 78 442 82
rect 606 78 610 82
rect 638 78 642 82
rect 774 78 778 82
rect 782 78 786 82
rect 886 78 890 82
rect 974 78 978 82
rect 1022 78 1026 82
rect 1054 78 1058 82
rect 1102 78 1106 82
rect 1206 78 1210 82
rect 1222 78 1226 82
rect 6 68 10 72
rect 30 68 34 72
rect 246 68 250 72
rect 390 68 394 72
rect 406 68 410 72
rect 534 68 538 72
rect 582 68 586 72
rect 646 68 650 72
rect 22 58 26 62
rect 54 58 58 62
rect 86 58 90 62
rect 150 58 154 62
rect 206 58 210 62
rect 214 58 218 62
rect 278 59 282 63
rect 374 58 378 62
rect 438 59 442 63
rect 702 68 706 72
rect 750 68 754 72
rect 798 68 802 72
rect 830 68 834 72
rect 846 68 850 72
rect 862 68 866 72
rect 910 68 914 72
rect 918 68 922 72
rect 942 68 946 72
rect 990 68 994 72
rect 1006 68 1010 72
rect 1030 68 1034 72
rect 1046 68 1050 72
rect 1110 68 1114 72
rect 1158 68 1162 72
rect 1182 68 1186 72
rect 1246 68 1250 72
rect 1254 68 1258 72
rect 1302 68 1306 72
rect 1318 68 1322 72
rect 1342 78 1346 82
rect 1398 78 1402 82
rect 1694 78 1698 82
rect 1910 78 1914 82
rect 1366 68 1370 72
rect 1382 68 1386 72
rect 1422 68 1426 72
rect 1510 68 1514 72
rect 1526 68 1530 72
rect 2038 78 2042 82
rect 2270 78 2274 82
rect 2334 78 2338 82
rect 2406 78 2410 82
rect 2414 78 2418 82
rect 2494 78 2498 82
rect 2534 78 2538 82
rect 2558 78 2562 82
rect 2574 78 2578 82
rect 2582 78 2586 82
rect 2598 78 2602 82
rect 2654 78 2658 82
rect 2686 78 2690 82
rect 1646 68 1650 72
rect 1702 68 1706 72
rect 1942 68 1946 72
rect 1958 68 1962 72
rect 2022 68 2026 72
rect 2054 68 2058 72
rect 2166 68 2170 72
rect 2222 68 2226 72
rect 2254 68 2258 72
rect 2286 68 2290 72
rect 2294 68 2298 72
rect 2446 68 2450 72
rect 2486 68 2490 72
rect 2518 68 2522 72
rect 2558 68 2562 72
rect 2606 68 2610 72
rect 2638 68 2642 72
rect 598 58 602 62
rect 694 58 698 62
rect 782 58 786 62
rect 806 58 810 62
rect 822 58 826 62
rect 838 58 842 62
rect 870 58 874 62
rect 950 58 954 62
rect 966 58 970 62
rect 998 58 1002 62
rect 1006 58 1010 62
rect 1054 58 1058 62
rect 1222 58 1226 62
rect 1270 58 1274 62
rect 1310 58 1314 62
rect 1358 58 1362 62
rect 1382 58 1386 62
rect 1470 58 1474 62
rect 1638 58 1642 62
rect 1718 58 1722 62
rect 1758 58 1762 62
rect 1782 58 1786 62
rect 1910 59 1914 63
rect 1974 58 1978 62
rect 1982 58 1986 62
rect 2006 58 2010 62
rect 2070 59 2074 63
rect 2166 58 2170 62
rect 2238 59 2242 63
rect 2294 58 2298 62
rect 2318 58 2322 62
rect 2326 58 2330 62
rect 2366 58 2370 62
rect 2390 58 2394 62
rect 2430 58 2434 62
rect 2438 58 2442 62
rect 2454 58 2458 62
rect 2494 58 2498 62
rect 2542 58 2546 62
rect 2606 58 2610 62
rect 2630 58 2634 62
rect 2678 58 2682 62
rect 222 48 226 52
rect 862 48 866 52
rect 894 48 898 52
rect 934 48 938 52
rect 1030 48 1034 52
rect 1126 48 1130 52
rect 1166 48 1170 52
rect 1182 48 1186 52
rect 1230 48 1234 52
rect 1406 48 1410 52
rect 1542 48 1546 52
rect 2398 48 2402 52
rect 2470 48 2474 52
rect 2622 48 2626 52
rect 86 38 90 42
rect 190 18 194 22
rect 366 18 370 22
rect 526 18 530 22
rect 1822 18 1826 22
rect 1998 18 2002 22
rect 2662 18 2666 22
rect 578 3 582 7
rect 585 3 589 7
rect 1602 3 1606 7
rect 1609 3 1613 7
<< metal2 >>
rect 46 1828 50 1832
rect 78 1828 82 1832
rect 102 1828 106 1832
rect 182 1828 186 1832
rect 222 1831 226 1832
rect 214 1828 226 1831
rect 254 1828 258 1832
rect 294 1828 298 1832
rect 366 1828 370 1832
rect 406 1828 410 1832
rect 454 1828 458 1832
rect 502 1831 506 1832
rect 502 1828 513 1831
rect 598 1828 602 1832
rect 638 1828 642 1832
rect 742 1828 746 1832
rect 758 1828 762 1832
rect 774 1831 778 1832
rect 790 1831 794 1832
rect 766 1828 778 1831
rect 782 1828 794 1831
rect 822 1828 826 1832
rect 838 1828 842 1832
rect 862 1828 866 1832
rect 934 1831 938 1832
rect 934 1828 945 1831
rect 102 1762 105 1768
rect 10 1758 14 1761
rect 58 1758 62 1761
rect 90 1758 94 1761
rect 6 1732 9 1738
rect 30 1722 33 1748
rect 6 1662 9 1708
rect 38 1651 41 1738
rect 46 1702 49 1748
rect 86 1742 89 1758
rect 182 1752 185 1828
rect 58 1738 62 1741
rect 34 1648 41 1651
rect 54 1662 57 1728
rect 78 1722 81 1738
rect 102 1722 105 1738
rect 62 1682 65 1698
rect 70 1681 73 1718
rect 70 1678 81 1681
rect 66 1668 70 1671
rect 46 1562 49 1618
rect 26 1548 30 1551
rect 54 1541 57 1658
rect 78 1652 81 1678
rect 86 1662 89 1718
rect 118 1712 121 1728
rect 126 1722 129 1738
rect 158 1732 161 1738
rect 138 1718 142 1721
rect 166 1712 169 1728
rect 182 1711 185 1748
rect 214 1742 217 1828
rect 366 1742 369 1828
rect 406 1742 409 1828
rect 454 1802 457 1828
rect 510 1792 513 1828
rect 576 1803 578 1807
rect 582 1803 585 1807
rect 589 1803 592 1807
rect 742 1802 745 1828
rect 758 1782 761 1828
rect 766 1792 769 1828
rect 782 1782 785 1828
rect 838 1802 841 1828
rect 790 1792 793 1798
rect 742 1772 745 1778
rect 446 1742 449 1748
rect 258 1738 262 1741
rect 306 1738 310 1741
rect 370 1738 374 1741
rect 214 1732 217 1738
rect 250 1728 254 1731
rect 202 1718 206 1721
rect 174 1708 185 1711
rect 110 1662 113 1668
rect 118 1662 121 1668
rect 142 1662 145 1708
rect 158 1682 161 1698
rect 174 1682 177 1708
rect 182 1682 185 1698
rect 238 1682 241 1728
rect 294 1722 297 1738
rect 302 1722 305 1728
rect 174 1662 177 1678
rect 198 1662 201 1668
rect 254 1662 257 1668
rect 194 1658 198 1661
rect 234 1658 238 1661
rect 134 1642 137 1648
rect 98 1638 102 1641
rect 50 1538 57 1541
rect 78 1552 81 1578
rect 6 1512 9 1528
rect 34 1518 38 1521
rect 6 1482 9 1488
rect 38 1472 41 1488
rect 46 1471 49 1538
rect 78 1532 81 1548
rect 54 1492 57 1498
rect 54 1471 57 1478
rect 46 1468 57 1471
rect 62 1472 65 1518
rect 70 1512 73 1528
rect 86 1492 89 1618
rect 134 1562 137 1588
rect 142 1582 145 1658
rect 270 1642 273 1718
rect 278 1652 281 1718
rect 326 1681 329 1718
rect 334 1712 337 1728
rect 326 1678 337 1681
rect 310 1672 313 1678
rect 290 1658 294 1661
rect 166 1592 169 1618
rect 206 1572 209 1618
rect 162 1568 166 1571
rect 142 1562 145 1568
rect 146 1548 150 1551
rect 206 1551 209 1568
rect 246 1552 249 1618
rect 198 1548 209 1551
rect 134 1542 137 1548
rect 94 1472 97 1538
rect 110 1522 113 1538
rect 118 1522 121 1538
rect 190 1532 193 1538
rect 198 1532 201 1548
rect 214 1541 217 1548
rect 210 1538 217 1541
rect 234 1538 238 1541
rect 254 1532 257 1558
rect 262 1532 265 1578
rect 286 1551 289 1618
rect 294 1562 297 1568
rect 318 1561 321 1678
rect 326 1662 329 1668
rect 334 1661 337 1678
rect 342 1672 345 1688
rect 350 1682 353 1718
rect 374 1712 377 1728
rect 382 1682 385 1728
rect 354 1668 358 1671
rect 334 1658 342 1661
rect 350 1582 353 1668
rect 378 1648 382 1651
rect 390 1631 393 1718
rect 398 1672 401 1738
rect 406 1732 409 1738
rect 454 1732 457 1738
rect 418 1668 422 1671
rect 430 1662 433 1678
rect 438 1652 441 1718
rect 454 1681 457 1728
rect 450 1678 457 1681
rect 470 1682 473 1718
rect 486 1712 489 1728
rect 494 1722 497 1748
rect 582 1742 585 1747
rect 494 1672 497 1688
rect 502 1672 505 1738
rect 522 1718 526 1721
rect 514 1678 518 1681
rect 542 1672 545 1688
rect 566 1672 569 1678
rect 522 1668 526 1671
rect 426 1638 430 1641
rect 382 1628 393 1631
rect 358 1572 361 1618
rect 314 1558 321 1561
rect 334 1552 337 1558
rect 350 1552 353 1558
rect 282 1548 289 1551
rect 322 1548 326 1551
rect 362 1548 366 1551
rect 302 1542 305 1548
rect 382 1542 385 1628
rect 390 1562 393 1618
rect 406 1552 409 1618
rect 446 1592 449 1668
rect 550 1662 553 1668
rect 582 1662 585 1668
rect 598 1662 601 1688
rect 622 1682 625 1718
rect 654 1692 657 1748
rect 610 1668 614 1671
rect 506 1658 510 1661
rect 538 1658 542 1661
rect 618 1648 622 1651
rect 550 1642 553 1648
rect 646 1642 649 1668
rect 474 1638 478 1641
rect 576 1603 578 1607
rect 582 1603 585 1607
rect 589 1603 592 1607
rect 506 1578 510 1581
rect 406 1542 409 1548
rect 278 1532 281 1538
rect 382 1532 385 1538
rect 390 1532 393 1538
rect 410 1528 414 1531
rect 422 1522 425 1548
rect 430 1532 433 1538
rect 102 1492 105 1518
rect 54 1462 57 1468
rect 102 1462 105 1468
rect 118 1462 121 1488
rect 130 1478 134 1481
rect 42 1458 46 1461
rect 82 1458 86 1461
rect 14 1382 17 1418
rect 22 1392 25 1458
rect 58 1448 62 1451
rect 90 1448 94 1451
rect 106 1448 110 1451
rect 138 1448 142 1451
rect 14 1292 17 1368
rect 70 1352 73 1358
rect 62 1348 70 1351
rect 22 1332 25 1348
rect 54 1312 57 1338
rect 62 1332 65 1348
rect 70 1332 73 1338
rect 30 1278 33 1308
rect 78 1292 81 1448
rect 158 1442 161 1518
rect 166 1462 169 1488
rect 182 1482 185 1518
rect 198 1472 201 1488
rect 178 1448 182 1451
rect 206 1451 209 1468
rect 214 1462 217 1468
rect 230 1462 233 1468
rect 238 1462 241 1478
rect 246 1472 249 1498
rect 254 1481 257 1518
rect 254 1478 262 1481
rect 270 1462 273 1518
rect 438 1502 441 1558
rect 470 1552 473 1578
rect 494 1562 497 1568
rect 566 1552 569 1558
rect 506 1548 510 1551
rect 470 1532 473 1548
rect 514 1488 518 1491
rect 294 1482 297 1488
rect 438 1482 441 1488
rect 506 1478 510 1481
rect 278 1472 281 1478
rect 438 1462 441 1468
rect 206 1448 217 1451
rect 166 1372 169 1418
rect 214 1392 217 1448
rect 150 1362 153 1368
rect 162 1358 166 1361
rect 98 1348 102 1351
rect 122 1348 126 1351
rect 150 1342 153 1348
rect 166 1342 169 1348
rect 130 1338 134 1341
rect 86 1322 89 1338
rect 174 1332 177 1358
rect 210 1348 214 1351
rect 222 1341 225 1368
rect 214 1338 225 1341
rect 94 1311 97 1328
rect 86 1308 97 1311
rect 42 1288 46 1291
rect 70 1272 73 1288
rect 58 1268 62 1271
rect 54 1252 57 1268
rect 86 1262 89 1308
rect 94 1282 97 1298
rect 66 1258 70 1261
rect 6 1132 9 1168
rect 58 1138 62 1141
rect 38 1112 41 1128
rect 46 1102 49 1108
rect 30 1082 33 1088
rect 54 1082 57 1138
rect 38 1072 41 1078
rect 10 1068 14 1071
rect 50 1068 54 1071
rect 62 1062 65 1118
rect 78 1112 81 1128
rect 102 1092 105 1328
rect 110 1312 113 1328
rect 182 1321 185 1338
rect 182 1318 190 1321
rect 114 1308 118 1311
rect 150 1278 153 1308
rect 126 1272 129 1278
rect 186 1268 190 1271
rect 186 1258 190 1261
rect 166 1252 169 1258
rect 182 1192 185 1228
rect 110 1142 113 1148
rect 118 1132 121 1138
rect 114 1128 118 1131
rect 110 1082 113 1088
rect 126 1081 129 1108
rect 134 1092 137 1118
rect 150 1102 153 1132
rect 126 1078 137 1081
rect 166 1078 169 1168
rect 198 1162 201 1308
rect 206 1282 209 1298
rect 214 1272 217 1338
rect 214 1252 217 1268
rect 222 1162 225 1298
rect 230 1292 233 1448
rect 238 1352 241 1458
rect 262 1392 265 1418
rect 270 1372 273 1458
rect 254 1332 257 1368
rect 274 1348 278 1351
rect 286 1342 289 1378
rect 294 1362 297 1418
rect 310 1362 313 1378
rect 294 1342 297 1348
rect 318 1332 321 1338
rect 246 1302 249 1318
rect 262 1312 265 1318
rect 238 1282 241 1288
rect 278 1282 281 1298
rect 302 1282 305 1318
rect 326 1292 329 1459
rect 358 1442 361 1458
rect 390 1412 393 1418
rect 342 1362 345 1388
rect 246 1272 249 1278
rect 262 1272 265 1278
rect 286 1272 289 1278
rect 326 1272 329 1278
rect 302 1262 305 1268
rect 174 1132 177 1138
rect 182 1092 185 1148
rect 206 1142 209 1148
rect 222 1142 225 1158
rect 238 1152 241 1238
rect 270 1192 273 1248
rect 270 1142 273 1148
rect 214 1132 217 1138
rect 262 1132 265 1138
rect 278 1122 281 1258
rect 310 1252 313 1268
rect 302 1172 305 1178
rect 290 1158 294 1161
rect 310 1161 313 1248
rect 318 1232 321 1258
rect 334 1162 337 1358
rect 342 1282 345 1358
rect 362 1348 366 1351
rect 406 1342 409 1438
rect 422 1371 425 1458
rect 462 1442 465 1478
rect 506 1458 510 1461
rect 534 1452 537 1498
rect 606 1482 609 1518
rect 574 1472 577 1478
rect 614 1472 617 1638
rect 646 1551 649 1558
rect 630 1492 633 1548
rect 662 1542 665 1738
rect 678 1692 681 1748
rect 710 1718 718 1721
rect 710 1682 713 1718
rect 674 1678 678 1681
rect 722 1678 726 1681
rect 634 1478 638 1481
rect 654 1472 657 1538
rect 670 1482 673 1678
rect 686 1642 689 1668
rect 722 1658 726 1661
rect 710 1592 713 1618
rect 726 1592 729 1648
rect 734 1642 737 1668
rect 750 1622 753 1748
rect 766 1592 769 1778
rect 894 1762 897 1768
rect 934 1752 937 1758
rect 834 1748 838 1751
rect 922 1748 926 1751
rect 774 1672 777 1748
rect 910 1742 913 1748
rect 822 1672 825 1728
rect 810 1658 814 1661
rect 822 1592 825 1658
rect 846 1562 849 1638
rect 886 1622 889 1678
rect 894 1662 897 1668
rect 918 1662 921 1738
rect 886 1592 889 1618
rect 910 1592 913 1648
rect 742 1542 745 1548
rect 750 1532 753 1548
rect 774 1532 777 1538
rect 742 1528 750 1531
rect 706 1518 710 1521
rect 726 1492 729 1518
rect 742 1492 745 1528
rect 538 1448 542 1451
rect 550 1442 553 1458
rect 558 1392 561 1458
rect 576 1403 578 1407
rect 582 1403 585 1407
rect 589 1403 592 1407
rect 622 1392 625 1438
rect 422 1368 433 1371
rect 422 1351 425 1358
rect 342 1262 345 1268
rect 350 1262 353 1278
rect 358 1272 361 1278
rect 374 1272 377 1338
rect 390 1332 393 1338
rect 382 1282 385 1288
rect 390 1272 393 1308
rect 422 1272 425 1288
rect 394 1248 398 1251
rect 414 1242 417 1248
rect 350 1172 353 1228
rect 430 1222 433 1368
rect 502 1362 505 1368
rect 558 1352 561 1358
rect 438 1272 441 1278
rect 454 1272 457 1348
rect 510 1332 513 1348
rect 518 1342 521 1348
rect 526 1332 529 1340
rect 486 1322 489 1328
rect 470 1252 473 1259
rect 462 1172 465 1218
rect 310 1158 318 1161
rect 306 1148 310 1151
rect 290 1138 294 1141
rect 214 1082 217 1098
rect 18 1058 25 1061
rect 42 1058 49 1061
rect 10 958 14 961
rect 6 932 9 938
rect 6 872 9 928
rect 22 852 25 1058
rect 34 1048 38 1051
rect 46 952 49 1058
rect 58 1048 62 1051
rect 78 1042 81 1078
rect 134 1072 137 1078
rect 198 1072 201 1078
rect 114 1068 118 1071
rect 86 1062 89 1068
rect 94 1062 97 1068
rect 158 1052 161 1058
rect 198 1052 201 1068
rect 214 1062 217 1068
rect 226 1058 230 1061
rect 134 1042 137 1048
rect 126 992 129 1038
rect 110 952 113 958
rect 118 952 121 958
rect 146 948 150 951
rect 30 922 33 948
rect 94 942 97 948
rect 222 942 225 1048
rect 242 1038 246 1041
rect 230 962 233 1018
rect 238 992 241 1028
rect 254 962 257 1118
rect 302 1082 305 1088
rect 302 1063 305 1068
rect 318 1032 321 1148
rect 334 1142 337 1158
rect 342 1142 345 1148
rect 350 1142 353 1168
rect 390 1151 393 1158
rect 422 1152 425 1168
rect 358 1142 361 1148
rect 462 1142 465 1168
rect 474 1138 478 1141
rect 334 1042 337 1078
rect 350 1062 353 1068
rect 366 1062 369 1108
rect 374 1082 377 1138
rect 418 1088 422 1091
rect 486 1082 489 1238
rect 494 1132 497 1288
rect 526 1282 529 1328
rect 574 1292 577 1348
rect 582 1322 585 1338
rect 534 1282 537 1288
rect 542 1262 545 1268
rect 554 1258 558 1261
rect 578 1258 582 1261
rect 502 1172 505 1258
rect 606 1222 609 1328
rect 614 1318 622 1321
rect 614 1272 617 1318
rect 622 1282 625 1288
rect 630 1282 633 1468
rect 678 1462 681 1488
rect 698 1458 702 1461
rect 726 1452 729 1488
rect 774 1462 777 1468
rect 738 1438 742 1441
rect 742 1398 750 1401
rect 742 1352 745 1398
rect 666 1348 670 1351
rect 678 1292 681 1348
rect 630 1272 633 1278
rect 646 1262 649 1268
rect 654 1232 657 1268
rect 662 1262 665 1268
rect 702 1242 705 1338
rect 726 1292 729 1318
rect 690 1238 694 1241
rect 576 1203 578 1207
rect 582 1203 585 1207
rect 589 1203 592 1207
rect 702 1172 705 1238
rect 742 1192 745 1348
rect 750 1282 753 1318
rect 766 1272 769 1368
rect 782 1282 785 1538
rect 798 1462 801 1518
rect 822 1472 825 1478
rect 838 1462 841 1548
rect 846 1492 849 1558
rect 866 1548 870 1551
rect 866 1538 870 1541
rect 894 1532 897 1548
rect 910 1542 913 1548
rect 854 1472 857 1488
rect 870 1472 873 1478
rect 854 1452 857 1468
rect 890 1458 894 1461
rect 838 1442 841 1448
rect 838 1382 841 1438
rect 870 1422 873 1458
rect 902 1442 905 1538
rect 918 1462 921 1658
rect 926 1552 929 1558
rect 942 1552 945 1828
rect 950 1828 954 1832
rect 966 1831 970 1832
rect 966 1828 977 1831
rect 950 1792 953 1828
rect 974 1792 977 1828
rect 1102 1828 1106 1832
rect 1126 1831 1130 1832
rect 1126 1828 1137 1831
rect 1102 1792 1105 1828
rect 1134 1792 1137 1828
rect 1222 1828 1226 1832
rect 1246 1831 1250 1832
rect 1238 1828 1250 1831
rect 1278 1828 1282 1832
rect 1310 1831 1314 1832
rect 1310 1828 1321 1831
rect 1350 1828 1354 1832
rect 1430 1831 1434 1832
rect 1454 1831 1458 1832
rect 1478 1831 1482 1832
rect 1502 1831 1506 1832
rect 1526 1831 1530 1832
rect 1430 1828 1441 1831
rect 1454 1828 1465 1831
rect 1478 1828 1489 1831
rect 1502 1828 1513 1831
rect 1142 1752 1145 1768
rect 1074 1748 1078 1751
rect 958 1682 961 1748
rect 1014 1742 1017 1748
rect 990 1732 993 1738
rect 1038 1672 1041 1738
rect 1062 1692 1065 1748
rect 1118 1722 1121 1748
rect 1206 1742 1209 1747
rect 1074 1718 1078 1721
rect 1118 1712 1121 1718
rect 1080 1703 1082 1707
rect 1086 1703 1089 1707
rect 1093 1703 1096 1707
rect 1154 1688 1158 1691
rect 1062 1682 1065 1688
rect 1166 1682 1169 1708
rect 1198 1692 1201 1738
rect 1206 1722 1209 1728
rect 1214 1692 1217 1698
rect 1222 1681 1225 1828
rect 1238 1792 1241 1828
rect 1318 1792 1321 1828
rect 1438 1792 1441 1828
rect 1462 1792 1465 1828
rect 1486 1792 1489 1828
rect 1510 1792 1513 1828
rect 1518 1828 1530 1831
rect 1558 1828 1562 1832
rect 1678 1831 1682 1832
rect 1702 1831 1706 1832
rect 1678 1828 1689 1831
rect 1518 1792 1521 1828
rect 1542 1752 1545 1768
rect 1254 1692 1257 1748
rect 1214 1678 1225 1681
rect 1078 1672 1081 1678
rect 974 1662 977 1668
rect 986 1658 990 1661
rect 990 1632 993 1658
rect 998 1652 1001 1658
rect 998 1562 1001 1568
rect 934 1492 937 1538
rect 950 1532 953 1558
rect 998 1532 1001 1538
rect 1006 1532 1009 1668
rect 1014 1662 1017 1668
rect 1022 1642 1025 1668
rect 1098 1659 1102 1662
rect 1190 1642 1193 1668
rect 1206 1622 1209 1678
rect 1214 1592 1217 1678
rect 1262 1632 1265 1748
rect 1274 1738 1278 1741
rect 1294 1732 1297 1748
rect 1334 1722 1337 1738
rect 1294 1672 1297 1718
rect 1358 1692 1361 1748
rect 1410 1718 1414 1721
rect 1310 1682 1313 1688
rect 1398 1682 1401 1718
rect 1346 1678 1350 1681
rect 1278 1663 1281 1668
rect 1014 1562 1017 1568
rect 1034 1558 1038 1561
rect 1046 1532 1049 1558
rect 1078 1552 1081 1558
rect 1174 1552 1177 1558
rect 1294 1552 1297 1668
rect 1326 1662 1329 1668
rect 1326 1592 1329 1618
rect 1334 1552 1337 1678
rect 1342 1632 1345 1658
rect 1366 1642 1369 1668
rect 1414 1662 1417 1668
rect 1358 1562 1361 1568
rect 1070 1542 1073 1548
rect 1078 1532 1081 1548
rect 1094 1542 1097 1548
rect 946 1488 950 1491
rect 950 1472 953 1488
rect 958 1482 961 1528
rect 982 1522 985 1528
rect 958 1462 961 1468
rect 858 1388 862 1391
rect 870 1352 873 1418
rect 886 1392 889 1438
rect 918 1421 921 1458
rect 918 1418 929 1421
rect 926 1392 929 1418
rect 790 1342 793 1348
rect 750 1263 753 1268
rect 766 1192 769 1258
rect 754 1168 758 1171
rect 558 1152 561 1168
rect 702 1152 705 1168
rect 538 1148 542 1151
rect 602 1148 606 1151
rect 630 1122 633 1138
rect 594 1118 598 1121
rect 638 1112 641 1128
rect 526 1082 529 1088
rect 450 1078 454 1081
rect 514 1078 518 1081
rect 422 1072 425 1078
rect 410 1058 414 1061
rect 242 948 246 951
rect 262 942 265 958
rect 286 952 289 958
rect 358 942 361 1038
rect 454 992 457 1068
rect 486 1062 489 1078
rect 558 1072 561 1088
rect 582 1072 585 1078
rect 598 1072 601 1088
rect 638 1082 641 1098
rect 546 1068 550 1071
rect 366 962 369 968
rect 406 952 409 968
rect 470 962 473 1018
rect 430 952 433 958
rect 370 938 374 941
rect 62 922 65 928
rect 30 862 33 868
rect 10 848 14 851
rect 30 822 33 858
rect 46 852 49 918
rect 78 892 81 928
rect 62 822 65 868
rect 86 862 89 918
rect 102 902 105 938
rect 134 932 137 938
rect 102 882 105 898
rect 138 888 142 891
rect 102 872 105 878
rect 90 858 97 861
rect 82 778 86 781
rect 6 732 9 758
rect 54 752 57 768
rect 94 762 97 858
rect 158 852 161 868
rect 166 852 169 918
rect 174 861 177 938
rect 222 921 225 938
rect 230 932 233 938
rect 214 918 225 921
rect 182 862 185 888
rect 190 882 193 888
rect 206 862 209 918
rect 214 882 217 918
rect 246 892 249 938
rect 270 892 273 918
rect 214 872 217 878
rect 286 875 289 908
rect 294 892 297 938
rect 358 932 361 938
rect 302 902 305 918
rect 318 912 321 928
rect 350 922 353 928
rect 422 922 425 938
rect 470 932 473 938
rect 478 932 481 1058
rect 506 1048 510 1051
rect 506 948 510 951
rect 486 942 489 948
rect 434 928 438 931
rect 494 931 497 948
rect 526 942 529 958
rect 534 942 537 1048
rect 550 1042 553 1058
rect 614 1042 617 1058
rect 654 1042 657 1088
rect 662 1062 665 1098
rect 678 1082 681 1148
rect 682 1038 686 1041
rect 578 1018 582 1021
rect 576 1003 578 1007
rect 582 1003 585 1007
rect 589 1003 592 1007
rect 638 992 641 1018
rect 662 982 665 1018
rect 614 952 617 958
rect 486 928 497 931
rect 502 932 505 938
rect 446 922 449 928
rect 462 922 465 928
rect 382 892 385 918
rect 478 892 481 918
rect 486 892 489 928
rect 542 922 545 948
rect 650 947 654 950
rect 554 928 558 931
rect 594 928 598 931
rect 370 888 377 891
rect 374 872 377 888
rect 494 872 497 878
rect 262 862 265 868
rect 174 858 182 861
rect 270 852 273 868
rect 326 862 329 868
rect 446 863 449 868
rect 102 772 105 778
rect 110 752 113 818
rect 174 782 177 818
rect 174 762 177 768
rect 270 762 273 768
rect 302 762 305 768
rect 310 762 313 768
rect 210 758 214 761
rect 234 758 238 761
rect 134 752 137 758
rect 166 752 169 758
rect 254 752 257 758
rect 350 752 353 818
rect 42 748 46 751
rect 186 748 190 751
rect 282 748 286 751
rect 22 742 25 748
rect 62 742 65 748
rect 54 722 57 738
rect 70 702 73 748
rect 86 722 89 748
rect 6 672 9 678
rect 22 672 25 688
rect 62 682 65 698
rect 102 692 105 748
rect 110 732 113 748
rect 158 742 161 748
rect 358 742 361 848
rect 462 792 465 868
rect 518 862 521 878
rect 478 832 481 858
rect 506 838 510 841
rect 446 762 449 768
rect 178 738 182 741
rect 262 738 270 741
rect 274 738 278 741
rect 418 738 422 741
rect 222 732 225 738
rect 246 732 249 738
rect 146 728 150 731
rect 118 712 121 728
rect 142 692 145 718
rect 214 712 217 728
rect 226 718 230 721
rect 174 692 177 708
rect 230 692 233 708
rect 182 682 185 688
rect 238 682 241 718
rect 246 682 249 688
rect 150 672 153 678
rect 90 668 94 671
rect 186 668 190 671
rect 46 662 49 668
rect 22 652 25 658
rect 38 652 41 658
rect 38 562 41 568
rect 6 532 9 538
rect 54 521 57 538
rect 50 518 57 521
rect 62 511 65 528
rect 54 508 65 511
rect 6 488 14 491
rect 34 488 38 491
rect 6 472 9 488
rect 54 472 57 508
rect 70 472 73 668
rect 126 662 129 668
rect 90 658 94 661
rect 78 652 81 658
rect 98 648 102 651
rect 118 642 121 658
rect 86 592 89 628
rect 114 558 118 561
rect 126 552 129 658
rect 158 652 161 658
rect 166 641 169 668
rect 202 658 206 661
rect 194 648 198 651
rect 158 638 169 641
rect 134 552 137 558
rect 114 548 118 551
rect 94 512 97 528
rect 66 468 70 471
rect 34 368 38 371
rect 54 351 57 468
rect 66 458 70 461
rect 78 452 81 508
rect 86 482 89 488
rect 102 472 105 528
rect 142 492 145 538
rect 150 522 153 528
rect 158 492 161 638
rect 190 592 193 638
rect 178 548 182 551
rect 166 542 169 548
rect 166 512 169 528
rect 102 462 105 468
rect 134 462 137 488
rect 146 478 150 481
rect 182 472 185 528
rect 206 522 209 538
rect 214 492 217 668
rect 222 662 225 668
rect 262 662 265 738
rect 278 692 281 728
rect 294 692 297 738
rect 334 722 337 728
rect 314 718 318 721
rect 378 718 382 721
rect 406 721 409 738
rect 402 718 409 721
rect 310 692 313 698
rect 374 692 377 708
rect 270 682 273 688
rect 414 682 417 728
rect 430 712 433 758
rect 450 748 454 751
rect 470 742 473 748
rect 450 738 454 741
rect 286 672 289 678
rect 250 658 254 661
rect 290 658 294 661
rect 262 592 265 648
rect 222 552 225 558
rect 294 542 297 578
rect 302 562 305 568
rect 310 552 313 668
rect 318 642 321 648
rect 334 592 337 678
rect 366 672 369 678
rect 342 662 345 668
rect 358 662 361 668
rect 390 662 393 678
rect 422 672 425 678
rect 378 658 382 661
rect 358 642 361 648
rect 398 642 401 668
rect 422 652 425 658
rect 430 642 433 688
rect 454 672 457 678
rect 454 652 457 658
rect 442 648 446 651
rect 438 642 441 648
rect 434 588 438 591
rect 378 548 382 551
rect 238 522 241 538
rect 246 502 249 538
rect 226 488 233 491
rect 230 472 233 488
rect 174 462 177 468
rect 94 452 97 458
rect 154 448 158 451
rect 182 451 185 468
rect 238 462 241 478
rect 246 462 249 498
rect 254 492 257 518
rect 294 482 297 538
rect 318 522 321 548
rect 326 542 329 548
rect 370 538 374 541
rect 354 528 358 531
rect 282 478 289 481
rect 306 478 310 481
rect 334 478 337 528
rect 366 482 369 538
rect 382 532 385 538
rect 390 522 393 528
rect 398 492 401 548
rect 406 502 409 548
rect 422 512 425 528
rect 422 492 425 498
rect 434 488 438 491
rect 378 478 382 481
rect 274 468 278 471
rect 286 462 289 478
rect 366 472 369 478
rect 390 472 393 488
rect 318 462 321 468
rect 174 448 185 451
rect 54 348 62 351
rect 122 348 126 351
rect 6 342 9 348
rect 62 342 65 348
rect 134 342 137 358
rect 150 352 153 358
rect 146 338 150 341
rect 162 338 166 341
rect 6 282 9 338
rect 38 282 41 298
rect 54 291 57 338
rect 118 332 121 338
rect 50 288 57 291
rect 86 292 89 298
rect 46 272 49 288
rect 94 272 97 318
rect 118 312 121 328
rect 134 312 137 338
rect 174 332 177 448
rect 198 392 201 458
rect 270 362 273 458
rect 278 362 281 368
rect 182 352 185 358
rect 198 352 201 358
rect 274 348 278 351
rect 202 338 206 341
rect 118 282 121 308
rect 142 272 145 318
rect 174 312 177 328
rect 150 282 153 288
rect 74 268 78 271
rect 38 262 41 268
rect 118 262 121 268
rect 106 258 110 261
rect 62 252 65 258
rect 158 252 161 308
rect 182 282 185 328
rect 214 322 217 328
rect 230 322 233 348
rect 238 342 241 348
rect 250 338 254 341
rect 286 332 289 458
rect 318 392 321 438
rect 334 362 337 418
rect 374 362 377 418
rect 302 352 305 358
rect 310 342 313 348
rect 406 342 409 468
rect 462 392 465 728
rect 470 682 473 738
rect 478 732 481 828
rect 510 752 513 758
rect 494 742 497 748
rect 518 742 521 818
rect 478 692 481 718
rect 470 492 473 678
rect 478 672 481 678
rect 494 662 497 718
rect 510 662 513 728
rect 518 722 521 738
rect 526 682 529 788
rect 534 761 537 888
rect 542 852 545 918
rect 574 902 577 918
rect 574 882 577 888
rect 562 878 569 881
rect 558 772 561 868
rect 566 852 569 878
rect 578 868 582 871
rect 598 862 601 918
rect 606 892 609 938
rect 678 882 681 948
rect 710 882 713 1058
rect 726 962 729 978
rect 734 972 737 1168
rect 754 1148 758 1151
rect 774 1102 777 1118
rect 782 1082 785 1278
rect 790 1272 793 1278
rect 802 1258 806 1261
rect 814 1242 817 1248
rect 814 1122 817 1238
rect 778 1078 782 1081
rect 774 1062 777 1068
rect 822 1062 825 1218
rect 830 1162 833 1338
rect 846 1272 849 1338
rect 878 1332 881 1378
rect 894 1302 897 1348
rect 926 1292 929 1348
rect 950 1332 953 1418
rect 838 1262 841 1268
rect 830 1112 833 1148
rect 838 1101 841 1258
rect 846 1222 849 1258
rect 918 1222 921 1278
rect 934 1272 937 1278
rect 966 1271 969 1518
rect 998 1492 1001 1528
rect 1022 1482 1025 1528
rect 998 1462 1001 1468
rect 978 1448 982 1451
rect 1022 1442 1025 1478
rect 1030 1452 1033 1528
rect 1082 1518 1086 1521
rect 1050 1478 1054 1481
rect 1042 1458 1046 1461
rect 1062 1452 1065 1518
rect 1080 1503 1082 1507
rect 1086 1503 1089 1507
rect 1093 1503 1096 1507
rect 1098 1478 1102 1481
rect 1098 1468 1102 1471
rect 1074 1458 1078 1461
rect 1034 1448 1038 1451
rect 1002 1358 1006 1361
rect 1026 1358 1030 1361
rect 986 1338 990 1341
rect 986 1328 990 1331
rect 1006 1322 1009 1338
rect 1034 1328 1038 1331
rect 966 1268 974 1271
rect 966 1232 969 1258
rect 974 1252 977 1268
rect 986 1266 990 1269
rect 998 1262 1001 1278
rect 1006 1272 1009 1318
rect 1022 1252 1025 1268
rect 1038 1262 1041 1318
rect 1054 1312 1057 1318
rect 1062 1292 1065 1348
rect 1070 1332 1073 1338
rect 1078 1332 1081 1378
rect 1110 1372 1113 1538
rect 1198 1532 1201 1538
rect 1118 1522 1121 1528
rect 1118 1502 1121 1518
rect 1118 1482 1121 1488
rect 1122 1478 1126 1481
rect 1150 1472 1153 1498
rect 1222 1482 1225 1488
rect 1210 1478 1214 1481
rect 1202 1468 1206 1471
rect 1118 1352 1121 1458
rect 1126 1452 1129 1468
rect 1150 1462 1153 1468
rect 1174 1452 1177 1458
rect 1182 1442 1185 1458
rect 1190 1442 1193 1468
rect 1126 1352 1129 1358
rect 1080 1303 1082 1307
rect 1086 1303 1089 1307
rect 1093 1303 1096 1307
rect 1102 1292 1105 1348
rect 1118 1341 1121 1348
rect 1118 1338 1129 1341
rect 1126 1332 1129 1338
rect 1114 1328 1118 1331
rect 1134 1292 1137 1418
rect 1166 1352 1169 1438
rect 1182 1432 1185 1438
rect 1182 1382 1185 1418
rect 1230 1392 1233 1548
rect 1270 1512 1273 1548
rect 1294 1532 1297 1548
rect 1334 1532 1337 1548
rect 1346 1538 1350 1541
rect 1286 1528 1294 1531
rect 1286 1482 1289 1528
rect 1330 1518 1334 1521
rect 1358 1482 1361 1548
rect 1366 1532 1369 1548
rect 1374 1542 1377 1548
rect 1382 1542 1385 1638
rect 1398 1632 1401 1658
rect 1422 1622 1425 1748
rect 1446 1672 1449 1748
rect 1470 1722 1473 1748
rect 1482 1658 1486 1661
rect 1366 1482 1369 1518
rect 1382 1472 1385 1538
rect 1406 1532 1409 1558
rect 1470 1552 1473 1658
rect 1442 1547 1446 1550
rect 1398 1492 1401 1508
rect 1346 1468 1350 1471
rect 1278 1452 1281 1458
rect 1286 1392 1289 1428
rect 1318 1392 1321 1468
rect 1406 1462 1409 1468
rect 1422 1462 1425 1538
rect 1470 1532 1473 1548
rect 1494 1482 1497 1748
rect 1534 1692 1537 1748
rect 1558 1711 1561 1828
rect 1600 1803 1602 1807
rect 1606 1803 1609 1807
rect 1613 1803 1616 1807
rect 1686 1792 1689 1828
rect 1694 1828 1706 1831
rect 1726 1828 1730 1832
rect 1750 1828 1754 1832
rect 1766 1828 1770 1832
rect 1782 1828 1786 1832
rect 1830 1828 1834 1832
rect 1886 1831 1890 1832
rect 1886 1828 1897 1831
rect 1942 1828 1946 1832
rect 1958 1828 1962 1832
rect 1982 1828 1986 1832
rect 2086 1828 2090 1832
rect 2382 1828 2386 1832
rect 2582 1828 2586 1832
rect 2686 1831 2690 1832
rect 2686 1828 2697 1831
rect 1694 1792 1697 1828
rect 1782 1802 1785 1828
rect 1734 1792 1737 1798
rect 1894 1792 1897 1828
rect 2694 1792 2697 1828
rect 2154 1778 2158 1781
rect 1834 1768 1838 1771
rect 1870 1752 1873 1768
rect 2022 1762 2025 1778
rect 2054 1762 2057 1768
rect 2222 1762 2225 1768
rect 2382 1762 2385 1768
rect 1666 1748 1670 1751
rect 1830 1748 1838 1751
rect 2086 1751 2089 1758
rect 2230 1752 2233 1758
rect 1606 1742 1609 1747
rect 1646 1732 1649 1738
rect 1654 1732 1657 1748
rect 1558 1708 1569 1711
rect 1546 1688 1550 1691
rect 1534 1682 1537 1688
rect 1534 1662 1537 1668
rect 1518 1592 1521 1658
rect 1502 1562 1505 1568
rect 1510 1552 1513 1568
rect 1542 1552 1545 1618
rect 1566 1592 1569 1708
rect 1582 1662 1585 1668
rect 1602 1658 1606 1661
rect 1550 1552 1553 1558
rect 1582 1542 1585 1648
rect 1600 1603 1602 1607
rect 1606 1603 1609 1607
rect 1613 1603 1616 1607
rect 1594 1568 1598 1571
rect 1646 1542 1649 1728
rect 1662 1682 1665 1718
rect 1670 1692 1673 1738
rect 1710 1731 1713 1748
rect 1718 1742 1721 1748
rect 1750 1732 1753 1738
rect 1774 1732 1777 1748
rect 1710 1728 1721 1731
rect 1718 1692 1721 1728
rect 1810 1688 1814 1691
rect 1718 1682 1721 1688
rect 1734 1672 1737 1678
rect 1702 1662 1705 1668
rect 1750 1663 1753 1668
rect 1678 1652 1681 1658
rect 1822 1652 1825 1658
rect 1718 1562 1721 1568
rect 1722 1558 1726 1561
rect 1818 1558 1822 1561
rect 1654 1551 1657 1558
rect 1686 1542 1689 1548
rect 1522 1538 1526 1541
rect 1706 1538 1710 1541
rect 1442 1468 1446 1471
rect 1430 1462 1433 1468
rect 1518 1462 1521 1528
rect 1534 1472 1537 1538
rect 1582 1492 1585 1538
rect 1670 1462 1673 1538
rect 1690 1528 1694 1531
rect 1734 1522 1737 1548
rect 1750 1542 1753 1548
rect 1798 1542 1801 1558
rect 1770 1538 1774 1541
rect 1786 1538 1790 1541
rect 1750 1512 1753 1538
rect 1766 1522 1769 1528
rect 1798 1522 1801 1538
rect 1710 1482 1713 1488
rect 1722 1478 1726 1481
rect 1734 1462 1737 1468
rect 1442 1458 1446 1461
rect 1530 1458 1534 1461
rect 1658 1458 1662 1461
rect 1142 1322 1145 1340
rect 1182 1332 1185 1338
rect 1186 1318 1190 1321
rect 1114 1288 1118 1291
rect 1158 1282 1161 1318
rect 1058 1278 1062 1281
rect 1018 1248 1022 1251
rect 902 1162 905 1218
rect 1014 1182 1017 1218
rect 1054 1212 1057 1248
rect 1062 1172 1065 1278
rect 1130 1268 1134 1271
rect 1142 1262 1145 1278
rect 1110 1252 1113 1258
rect 1174 1252 1177 1318
rect 1198 1292 1201 1328
rect 1206 1282 1209 1368
rect 1230 1282 1233 1388
rect 1242 1348 1246 1351
rect 1238 1272 1241 1278
rect 1194 1268 1198 1271
rect 1246 1262 1249 1288
rect 1270 1272 1273 1338
rect 1278 1292 1281 1318
rect 1286 1292 1289 1318
rect 1302 1272 1305 1278
rect 1186 1258 1190 1261
rect 1138 1248 1142 1251
rect 1154 1238 1158 1241
rect 1166 1232 1169 1238
rect 1138 1228 1142 1231
rect 1214 1202 1217 1218
rect 1254 1192 1257 1258
rect 1262 1242 1265 1248
rect 1090 1158 1094 1161
rect 854 1142 857 1158
rect 870 1132 873 1148
rect 886 1142 889 1148
rect 902 1142 905 1158
rect 1062 1152 1065 1158
rect 922 1147 926 1150
rect 882 1128 886 1131
rect 902 1112 905 1118
rect 830 1098 841 1101
rect 830 1072 833 1098
rect 846 1092 849 1108
rect 870 1092 873 1098
rect 742 1052 745 1059
rect 798 992 801 1058
rect 822 1052 825 1058
rect 806 1042 809 1048
rect 838 1012 841 1078
rect 862 1042 865 1058
rect 870 1052 873 1088
rect 902 1072 905 1108
rect 934 1082 937 1138
rect 998 1132 1001 1148
rect 1022 1142 1025 1148
rect 1050 1138 1054 1141
rect 1078 1132 1081 1138
rect 1126 1132 1129 1148
rect 1174 1142 1177 1148
rect 1134 1132 1137 1138
rect 1166 1132 1169 1138
rect 986 1128 990 1131
rect 1106 1128 1110 1131
rect 1230 1131 1233 1148
rect 998 1122 1001 1128
rect 986 1118 990 1121
rect 1006 1112 1009 1128
rect 1002 1078 1006 1081
rect 890 1068 894 1071
rect 894 1052 897 1058
rect 906 1048 910 1051
rect 846 992 849 1038
rect 738 968 742 971
rect 586 848 590 851
rect 566 832 569 848
rect 622 822 625 858
rect 630 852 633 868
rect 654 842 657 858
rect 726 842 729 948
rect 750 932 753 988
rect 774 962 777 978
rect 810 968 814 971
rect 842 968 846 971
rect 870 962 873 968
rect 790 921 793 938
rect 814 932 817 948
rect 790 918 801 921
rect 758 892 761 918
rect 766 882 769 898
rect 750 872 753 878
rect 734 863 737 868
rect 766 862 769 868
rect 774 858 782 861
rect 576 803 578 807
rect 582 803 585 807
rect 589 803 592 807
rect 578 788 582 791
rect 602 768 606 771
rect 534 758 542 761
rect 542 742 545 748
rect 550 682 553 758
rect 558 752 561 768
rect 534 662 537 668
rect 558 662 561 708
rect 566 702 569 768
rect 646 741 649 838
rect 654 762 657 818
rect 726 762 729 768
rect 718 752 721 758
rect 726 752 729 758
rect 742 752 745 818
rect 658 747 662 750
rect 694 742 697 748
rect 646 738 657 741
rect 614 672 617 678
rect 602 668 606 671
rect 594 638 598 641
rect 490 618 494 621
rect 576 603 578 607
rect 582 603 585 607
rect 589 603 592 607
rect 526 562 529 568
rect 494 551 497 558
rect 510 542 513 548
rect 542 542 545 588
rect 510 472 513 538
rect 494 463 497 468
rect 526 462 529 468
rect 494 352 497 358
rect 502 352 505 368
rect 534 352 537 538
rect 542 472 545 488
rect 550 482 553 528
rect 574 512 577 518
rect 574 482 577 488
rect 606 482 609 658
rect 614 522 617 668
rect 622 542 625 708
rect 630 612 633 658
rect 646 652 649 658
rect 638 642 641 648
rect 654 642 657 738
rect 678 712 681 738
rect 694 672 697 728
rect 666 668 670 671
rect 682 658 686 661
rect 702 651 705 718
rect 698 648 705 651
rect 654 592 657 638
rect 662 572 665 618
rect 694 552 697 568
rect 702 562 705 648
rect 718 702 721 738
rect 742 732 745 748
rect 750 742 753 848
rect 774 792 777 858
rect 798 772 801 918
rect 822 892 825 948
rect 846 932 849 948
rect 862 902 865 948
rect 886 942 889 948
rect 894 942 897 1048
rect 950 1042 953 1078
rect 958 1072 961 1078
rect 990 1072 993 1078
rect 1014 1071 1017 1098
rect 1030 1082 1033 1118
rect 1070 1102 1073 1118
rect 1080 1103 1082 1107
rect 1086 1103 1089 1107
rect 1093 1103 1096 1107
rect 1010 1068 1017 1071
rect 1034 1068 1038 1071
rect 974 1062 977 1068
rect 958 1052 961 1058
rect 1054 1052 1057 1078
rect 1110 1072 1113 1088
rect 1066 1068 1070 1071
rect 1078 1062 1081 1068
rect 1118 1061 1121 1118
rect 1114 1058 1121 1061
rect 1134 1062 1137 1128
rect 1146 1118 1150 1121
rect 1158 1062 1161 1068
rect 970 1048 974 1051
rect 1074 1038 1078 1041
rect 1086 1022 1089 1048
rect 1118 1042 1121 1048
rect 1150 1032 1153 1058
rect 1166 1042 1169 1128
rect 1182 1082 1185 1118
rect 1206 1092 1209 1128
rect 1226 1128 1233 1131
rect 1242 1128 1246 1131
rect 1238 1092 1241 1128
rect 1254 1092 1257 1148
rect 1262 1132 1265 1138
rect 1182 1072 1185 1078
rect 1190 1072 1193 1078
rect 1270 1072 1273 1268
rect 1286 1252 1289 1258
rect 1286 1172 1289 1228
rect 1326 1202 1329 1418
rect 1358 1402 1361 1418
rect 1378 1388 1382 1391
rect 1438 1352 1441 1398
rect 1518 1372 1521 1458
rect 1598 1452 1601 1458
rect 1598 1422 1601 1448
rect 1600 1403 1602 1407
rect 1606 1403 1609 1407
rect 1613 1403 1616 1407
rect 1418 1348 1422 1351
rect 1342 1322 1345 1348
rect 1350 1332 1353 1348
rect 1350 1272 1353 1328
rect 1478 1292 1481 1348
rect 1566 1322 1569 1347
rect 1582 1342 1585 1348
rect 1502 1282 1505 1318
rect 1590 1292 1593 1318
rect 1614 1292 1617 1338
rect 1638 1292 1641 1418
rect 1670 1392 1673 1458
rect 1758 1422 1761 1448
rect 1758 1392 1761 1418
rect 1766 1402 1769 1518
rect 1782 1472 1785 1508
rect 1806 1492 1809 1518
rect 1814 1502 1817 1558
rect 1822 1522 1825 1528
rect 1806 1470 1809 1478
rect 1814 1472 1817 1498
rect 1822 1482 1825 1488
rect 1774 1442 1777 1458
rect 1782 1392 1785 1468
rect 1790 1462 1793 1468
rect 1830 1462 1833 1748
rect 1838 1732 1841 1738
rect 1854 1682 1857 1738
rect 1870 1732 1873 1748
rect 1910 1722 1913 1738
rect 1910 1672 1913 1718
rect 1934 1702 1937 1748
rect 2006 1742 2009 1748
rect 2194 1748 2198 1751
rect 2250 1748 2254 1751
rect 2174 1742 2177 1748
rect 1994 1738 1998 1741
rect 2194 1738 2198 1741
rect 2038 1722 2041 1738
rect 1838 1662 1841 1668
rect 1914 1658 1918 1661
rect 1982 1652 1985 1659
rect 1990 1652 1993 1718
rect 1846 1592 1849 1648
rect 2030 1642 2033 1708
rect 2054 1682 2057 1728
rect 2070 1712 2073 1738
rect 2062 1692 2065 1698
rect 2070 1682 2073 1708
rect 2104 1703 2106 1707
rect 2110 1703 2113 1707
rect 2117 1703 2120 1707
rect 2086 1682 2089 1688
rect 2094 1678 2102 1681
rect 2042 1638 2046 1641
rect 1878 1562 1881 1638
rect 1914 1568 1918 1571
rect 1838 1552 1841 1558
rect 1934 1552 1937 1608
rect 1958 1562 1961 1578
rect 1998 1562 2001 1568
rect 1922 1548 1926 1551
rect 1994 1548 1998 1551
rect 1838 1492 1841 1528
rect 1778 1368 1782 1371
rect 1762 1358 1766 1361
rect 1682 1338 1686 1341
rect 1474 1278 1478 1281
rect 1538 1278 1542 1281
rect 1594 1278 1598 1281
rect 1526 1272 1529 1278
rect 1410 1268 1414 1271
rect 1466 1268 1470 1271
rect 1334 1262 1337 1268
rect 1386 1258 1390 1261
rect 1382 1242 1385 1258
rect 1298 1168 1302 1171
rect 1314 1168 1318 1171
rect 1286 1152 1289 1168
rect 1342 1162 1345 1168
rect 1390 1162 1393 1248
rect 1398 1232 1401 1268
rect 1422 1242 1425 1248
rect 1446 1232 1449 1268
rect 1454 1262 1457 1268
rect 1474 1258 1478 1261
rect 1486 1232 1489 1268
rect 1542 1262 1545 1278
rect 1582 1272 1585 1278
rect 1510 1252 1513 1258
rect 1526 1252 1529 1258
rect 1302 1142 1305 1148
rect 1318 1132 1321 1138
rect 1326 1132 1329 1158
rect 1358 1152 1361 1158
rect 1346 1148 1350 1151
rect 1342 1142 1345 1148
rect 1406 1142 1409 1148
rect 1414 1142 1417 1198
rect 1446 1152 1449 1198
rect 1486 1142 1489 1228
rect 1518 1162 1521 1168
rect 1494 1152 1497 1158
rect 1502 1152 1505 1158
rect 1526 1142 1529 1178
rect 1534 1162 1537 1218
rect 1550 1182 1553 1268
rect 1590 1258 1598 1261
rect 1582 1252 1585 1258
rect 1566 1248 1574 1251
rect 1566 1242 1569 1248
rect 1566 1192 1569 1238
rect 1590 1192 1593 1258
rect 1600 1203 1602 1207
rect 1606 1203 1609 1207
rect 1613 1203 1616 1207
rect 1590 1152 1593 1188
rect 1354 1138 1358 1141
rect 1442 1138 1446 1141
rect 1366 1132 1369 1138
rect 1398 1132 1401 1138
rect 1470 1132 1473 1138
rect 1418 1128 1422 1131
rect 1338 1088 1342 1091
rect 1374 1082 1377 1118
rect 1234 1068 1238 1071
rect 1202 1048 1206 1051
rect 918 912 921 948
rect 934 932 937 938
rect 878 892 881 898
rect 886 892 889 898
rect 934 892 937 928
rect 814 863 817 888
rect 846 862 849 878
rect 942 862 945 1018
rect 982 1002 985 1018
rect 950 952 953 958
rect 958 941 961 958
rect 974 952 977 958
rect 982 942 985 978
rect 1006 942 1009 978
rect 1014 942 1017 948
rect 950 938 961 941
rect 994 938 998 941
rect 758 762 761 768
rect 718 682 721 698
rect 718 642 721 678
rect 734 672 737 708
rect 750 692 753 738
rect 758 722 761 758
rect 770 748 774 751
rect 782 742 785 748
rect 846 742 849 858
rect 950 772 953 938
rect 966 932 969 938
rect 986 928 990 931
rect 966 872 969 878
rect 986 868 990 871
rect 950 762 953 768
rect 894 752 897 758
rect 790 712 793 718
rect 838 712 841 728
rect 854 711 857 747
rect 902 742 905 758
rect 954 748 958 751
rect 922 738 926 741
rect 854 708 865 711
rect 750 632 753 659
rect 714 628 718 631
rect 718 592 721 608
rect 706 558 713 561
rect 634 547 638 550
rect 674 548 678 551
rect 686 542 689 548
rect 670 532 673 538
rect 662 492 665 498
rect 694 492 697 518
rect 554 478 558 481
rect 690 478 694 481
rect 702 472 705 478
rect 626 468 630 471
rect 658 468 662 471
rect 650 458 654 461
rect 698 458 702 461
rect 558 422 561 458
rect 558 362 561 418
rect 576 403 578 407
rect 582 403 585 407
rect 589 403 592 407
rect 630 392 633 458
rect 450 348 454 351
rect 566 351 569 388
rect 622 362 625 368
rect 638 362 641 428
rect 470 342 473 348
rect 450 338 454 341
rect 238 322 241 328
rect 358 321 361 338
rect 358 318 366 321
rect 222 292 225 318
rect 206 282 209 288
rect 286 282 289 308
rect 218 278 222 281
rect 166 272 169 278
rect 182 272 185 278
rect 294 272 297 318
rect 406 312 409 338
rect 414 332 417 338
rect 326 282 329 298
rect 414 291 417 328
rect 414 288 422 291
rect 438 272 441 318
rect 254 262 257 268
rect 310 262 313 268
rect 366 262 369 268
rect 274 258 278 261
rect 470 262 473 338
rect 174 252 177 258
rect 294 252 297 258
rect 202 248 206 251
rect 242 248 246 251
rect 390 232 393 258
rect 358 152 361 228
rect 438 192 441 258
rect 454 252 457 259
rect 398 152 401 158
rect 26 148 30 151
rect 98 148 102 151
rect 234 148 238 151
rect 338 148 342 151
rect 434 148 438 151
rect 14 122 17 128
rect 6 72 9 78
rect 22 62 25 118
rect 30 52 33 68
rect 38 62 41 148
rect 46 122 49 128
rect 126 92 129 138
rect 90 88 94 91
rect 54 82 57 88
rect 54 62 57 78
rect 142 62 145 148
rect 158 142 161 148
rect 262 142 265 148
rect 158 82 161 88
rect 90 58 94 61
rect 198 61 201 128
rect 262 92 265 138
rect 278 131 281 148
rect 310 142 313 148
rect 278 128 286 131
rect 414 122 417 138
rect 430 132 433 148
rect 462 132 465 218
rect 470 152 473 258
rect 486 232 489 258
rect 502 142 505 348
rect 634 348 638 351
rect 662 282 665 358
rect 670 281 673 428
rect 694 392 697 448
rect 710 362 713 558
rect 738 548 742 551
rect 718 512 721 548
rect 730 538 737 541
rect 718 482 721 508
rect 734 492 737 538
rect 726 462 729 478
rect 750 472 753 548
rect 758 542 761 688
rect 782 632 785 658
rect 798 571 801 668
rect 838 662 841 708
rect 862 692 865 708
rect 846 672 849 688
rect 854 672 857 678
rect 822 652 825 658
rect 870 651 873 668
rect 894 662 897 698
rect 934 682 937 748
rect 974 742 977 748
rect 902 662 905 668
rect 942 662 945 718
rect 882 658 886 661
rect 894 652 897 658
rect 842 648 873 651
rect 886 642 889 648
rect 926 642 929 648
rect 818 638 822 641
rect 906 638 910 641
rect 790 568 801 571
rect 806 572 809 588
rect 846 572 849 628
rect 902 592 905 638
rect 950 612 953 738
rect 958 732 961 738
rect 970 728 974 731
rect 982 712 985 858
rect 1006 852 1009 898
rect 1022 872 1025 1008
rect 1038 982 1041 1018
rect 1062 942 1065 947
rect 1094 942 1097 948
rect 1030 902 1033 928
rect 1046 882 1049 938
rect 1054 892 1057 908
rect 1080 903 1082 907
rect 1086 903 1089 907
rect 1093 903 1096 907
rect 1110 892 1113 948
rect 1174 942 1177 947
rect 1138 938 1142 941
rect 1078 872 1081 888
rect 1086 872 1089 878
rect 1018 868 1022 871
rect 1118 862 1121 868
rect 1126 862 1129 868
rect 1134 862 1137 918
rect 1182 892 1185 1018
rect 1222 962 1225 1058
rect 1246 1032 1249 1068
rect 1294 1062 1297 1068
rect 1302 1063 1305 1078
rect 1366 1062 1369 1068
rect 1246 992 1249 1028
rect 1278 992 1281 1038
rect 1294 972 1297 1058
rect 1382 1051 1385 1128
rect 1430 1102 1433 1118
rect 1446 1082 1449 1118
rect 1394 1059 1398 1062
rect 1430 1062 1433 1078
rect 1442 1058 1446 1061
rect 1382 1048 1393 1051
rect 1206 942 1209 948
rect 1206 892 1209 898
rect 1142 862 1145 888
rect 1150 862 1153 868
rect 1018 858 1022 861
rect 1014 752 1017 798
rect 1006 742 1009 748
rect 962 688 966 691
rect 982 672 985 708
rect 990 702 993 718
rect 1014 681 1017 748
rect 1022 732 1025 738
rect 1038 732 1041 738
rect 1014 678 1025 681
rect 1014 662 1017 668
rect 978 658 982 661
rect 1002 658 1006 661
rect 770 548 774 551
rect 790 542 793 568
rect 798 552 801 558
rect 766 492 769 538
rect 790 532 793 538
rect 814 532 817 548
rect 782 481 785 518
rect 774 478 785 481
rect 746 458 750 461
rect 758 452 761 458
rect 698 348 702 351
rect 678 292 681 318
rect 670 278 681 281
rect 542 262 545 268
rect 522 258 526 261
rect 558 242 561 278
rect 678 272 681 278
rect 606 263 609 268
rect 514 218 518 221
rect 538 168 542 171
rect 558 142 561 238
rect 638 232 641 258
rect 576 203 578 207
rect 582 203 585 207
rect 589 203 592 207
rect 654 192 657 268
rect 666 238 670 241
rect 678 182 681 268
rect 686 262 689 278
rect 710 262 713 358
rect 766 352 769 438
rect 774 392 777 478
rect 790 472 793 498
rect 822 492 825 548
rect 830 482 833 518
rect 782 462 785 468
rect 822 452 825 459
rect 830 432 833 478
rect 846 462 849 568
rect 950 552 953 608
rect 982 602 985 658
rect 982 552 985 598
rect 990 562 993 618
rect 894 512 897 547
rect 910 542 913 548
rect 990 542 993 558
rect 1022 552 1025 678
rect 1030 572 1033 718
rect 1046 662 1049 858
rect 1166 852 1169 878
rect 1238 852 1241 918
rect 1246 862 1249 948
rect 1262 902 1265 928
rect 1282 918 1286 921
rect 1270 882 1273 918
rect 1302 882 1305 888
rect 1318 882 1321 918
rect 1342 872 1345 947
rect 1358 872 1361 938
rect 1270 863 1273 868
rect 1302 862 1305 868
rect 1150 832 1153 838
rect 1054 662 1057 818
rect 1174 792 1177 828
rect 1086 751 1089 758
rect 1246 752 1249 858
rect 1318 822 1321 858
rect 1358 822 1361 858
rect 1374 832 1377 948
rect 1390 941 1393 1048
rect 1446 992 1449 1048
rect 1462 972 1465 1128
rect 1470 1092 1473 1128
rect 1478 1082 1481 1118
rect 1402 958 1406 961
rect 1422 952 1425 968
rect 1390 938 1398 941
rect 1382 932 1385 938
rect 1390 863 1393 918
rect 1398 792 1401 938
rect 1406 752 1409 948
rect 1430 942 1433 948
rect 1438 932 1441 938
rect 1414 842 1417 858
rect 1422 792 1425 928
rect 1454 892 1457 968
rect 1462 892 1465 958
rect 1470 942 1473 1068
rect 1486 1062 1489 1108
rect 1494 1092 1497 1138
rect 1502 1132 1505 1138
rect 1550 1122 1553 1128
rect 1534 1070 1537 1098
rect 1550 1072 1553 1078
rect 1558 1072 1561 1098
rect 1502 1062 1505 1068
rect 1550 1052 1553 1068
rect 1582 1062 1585 1078
rect 1590 962 1593 1148
rect 1598 1092 1601 1188
rect 1630 1142 1633 1147
rect 1630 1082 1633 1088
rect 1638 1082 1641 1128
rect 1622 1062 1625 1078
rect 1600 1003 1602 1007
rect 1606 1003 1609 1007
rect 1613 1003 1616 1007
rect 1614 972 1617 978
rect 1578 948 1582 951
rect 1454 882 1457 888
rect 1114 748 1118 751
rect 1158 722 1161 748
rect 1182 742 1185 748
rect 1070 662 1073 718
rect 1080 703 1082 707
rect 1086 703 1089 707
rect 1093 703 1096 707
rect 1078 662 1081 688
rect 1118 662 1121 668
rect 1150 662 1153 718
rect 1174 702 1177 718
rect 1198 692 1201 748
rect 1214 742 1217 747
rect 1246 742 1249 748
rect 1290 718 1294 721
rect 1190 672 1193 678
rect 1206 672 1209 708
rect 1046 652 1049 658
rect 1078 652 1081 658
rect 1054 632 1057 638
rect 1098 588 1102 591
rect 1126 582 1129 658
rect 1142 642 1145 648
rect 1166 622 1169 658
rect 1182 652 1185 658
rect 1174 632 1177 638
rect 1034 558 1038 561
rect 1002 548 1006 551
rect 1022 542 1025 548
rect 934 522 937 528
rect 882 488 886 491
rect 782 351 785 368
rect 822 352 825 398
rect 838 392 841 458
rect 894 452 897 478
rect 902 472 905 478
rect 918 472 921 488
rect 926 472 929 478
rect 910 462 913 468
rect 934 462 937 518
rect 942 492 945 508
rect 966 492 969 518
rect 1014 501 1017 518
rect 1014 498 1025 501
rect 954 478 958 481
rect 986 478 990 481
rect 1014 472 1017 488
rect 970 468 982 471
rect 922 458 926 461
rect 958 452 961 458
rect 870 392 873 448
rect 830 372 833 378
rect 862 372 865 378
rect 982 372 985 418
rect 854 352 857 358
rect 990 352 993 438
rect 1022 361 1025 498
rect 1030 462 1033 468
rect 1018 358 1025 361
rect 1038 351 1041 518
rect 1054 472 1057 518
rect 1054 452 1057 458
rect 1046 392 1049 438
rect 1034 348 1041 351
rect 722 318 726 321
rect 726 282 729 288
rect 702 252 705 258
rect 758 252 761 259
rect 718 242 721 248
rect 630 162 633 168
rect 590 152 593 158
rect 638 152 641 158
rect 654 152 657 158
rect 686 152 689 218
rect 694 162 697 168
rect 714 158 718 161
rect 674 148 678 151
rect 706 148 710 151
rect 490 128 494 131
rect 470 122 473 128
rect 502 122 505 128
rect 394 118 398 121
rect 470 102 473 118
rect 278 82 281 88
rect 342 82 345 88
rect 438 82 441 88
rect 502 82 505 88
rect 246 72 249 78
rect 406 72 409 78
rect 526 72 529 118
rect 558 92 561 138
rect 570 128 574 131
rect 582 72 585 98
rect 530 68 534 71
rect 198 58 206 61
rect 218 58 222 61
rect 390 62 393 68
rect 150 52 153 58
rect 278 52 281 59
rect 378 58 382 61
rect 598 62 601 138
rect 606 82 609 138
rect 614 92 617 148
rect 630 142 633 148
rect 686 142 689 148
rect 658 138 662 141
rect 722 138 726 141
rect 674 128 678 131
rect 750 122 753 148
rect 766 132 769 318
rect 782 262 785 328
rect 814 291 817 348
rect 846 292 849 348
rect 910 312 913 348
rect 950 332 953 348
rect 930 328 934 331
rect 950 322 953 328
rect 814 288 822 291
rect 834 288 838 291
rect 918 291 921 318
rect 918 288 929 291
rect 926 282 929 288
rect 966 272 969 338
rect 974 332 977 348
rect 974 282 977 328
rect 982 312 985 338
rect 990 332 993 338
rect 990 292 993 318
rect 998 282 1001 348
rect 1014 342 1017 348
rect 1022 322 1025 338
rect 1038 332 1041 348
rect 1018 288 1022 291
rect 998 272 1001 278
rect 1038 272 1041 318
rect 1054 312 1057 428
rect 1062 362 1065 568
rect 1086 552 1089 578
rect 1154 547 1158 550
rect 1080 503 1082 507
rect 1086 503 1089 507
rect 1093 503 1096 507
rect 1082 478 1086 481
rect 1090 448 1094 451
rect 1094 351 1097 418
rect 1102 322 1105 538
rect 1114 458 1118 461
rect 1110 442 1113 448
rect 1126 352 1129 538
rect 1174 472 1177 538
rect 1190 532 1193 668
rect 1210 658 1214 661
rect 1222 592 1225 638
rect 1230 582 1233 698
rect 1254 692 1257 708
rect 1278 682 1281 718
rect 1242 668 1246 671
rect 1238 642 1241 658
rect 1254 652 1257 678
rect 1274 668 1278 671
rect 1270 642 1273 658
rect 1230 572 1233 578
rect 1238 572 1241 618
rect 1278 612 1281 658
rect 1274 568 1278 571
rect 1198 542 1201 548
rect 1206 542 1209 568
rect 1230 552 1233 558
rect 1286 552 1289 718
rect 1350 712 1353 747
rect 1366 742 1369 748
rect 1382 692 1385 748
rect 1354 688 1358 691
rect 1338 668 1342 671
rect 1214 542 1217 548
rect 1190 482 1193 528
rect 1222 492 1225 548
rect 1238 542 1241 548
rect 1254 542 1257 548
rect 1270 542 1273 548
rect 1282 538 1286 541
rect 1274 528 1278 531
rect 1274 478 1278 481
rect 1198 463 1201 468
rect 1214 442 1217 468
rect 1230 432 1233 468
rect 1238 392 1241 478
rect 1266 458 1270 461
rect 1278 452 1281 468
rect 1286 462 1289 538
rect 1294 532 1297 638
rect 1302 562 1305 618
rect 1318 602 1321 658
rect 1350 622 1353 668
rect 1390 652 1393 718
rect 1398 692 1401 718
rect 1406 702 1409 748
rect 1438 732 1441 758
rect 1446 742 1449 748
rect 1470 742 1473 938
rect 1526 922 1529 938
rect 1550 932 1553 938
rect 1622 932 1625 1058
rect 1630 992 1633 1068
rect 1638 1052 1641 1058
rect 1646 972 1649 1138
rect 1654 1092 1657 1118
rect 1662 1072 1665 1328
rect 1678 1172 1681 1268
rect 1686 1192 1689 1258
rect 1694 1192 1697 1358
rect 1790 1352 1793 1448
rect 1746 1348 1750 1351
rect 1758 1292 1761 1338
rect 1766 1332 1769 1348
rect 1806 1292 1809 1438
rect 1814 1342 1817 1458
rect 1826 1348 1830 1351
rect 1834 1338 1838 1341
rect 1742 1262 1745 1288
rect 1770 1268 1774 1271
rect 1678 1162 1681 1168
rect 1694 1152 1697 1188
rect 1734 1132 1737 1178
rect 1742 1122 1745 1148
rect 1710 1102 1713 1118
rect 1734 1112 1737 1118
rect 1674 1068 1678 1071
rect 1662 1062 1665 1068
rect 1702 1062 1705 1068
rect 1690 1058 1694 1061
rect 1654 1042 1657 1058
rect 1710 1052 1713 1078
rect 1718 1062 1721 1068
rect 1674 1048 1678 1051
rect 1642 948 1646 951
rect 1662 942 1665 1018
rect 1690 958 1694 961
rect 1710 952 1713 1048
rect 1726 1042 1729 1088
rect 1742 1072 1745 1078
rect 1750 1052 1753 1248
rect 1766 1102 1769 1268
rect 1794 1258 1798 1261
rect 1806 1252 1809 1278
rect 1782 1222 1785 1228
rect 1782 1132 1785 1218
rect 1814 1172 1817 1338
rect 1826 1268 1830 1271
rect 1838 1182 1841 1218
rect 1794 1148 1798 1151
rect 1806 1142 1809 1148
rect 1822 1142 1825 1158
rect 1838 1142 1841 1147
rect 1774 1092 1777 1118
rect 1774 1062 1777 1068
rect 1782 1062 1785 1098
rect 1798 1092 1801 1138
rect 1790 1082 1793 1088
rect 1826 1068 1830 1071
rect 1782 1052 1785 1058
rect 1750 1042 1753 1048
rect 1762 1038 1766 1041
rect 1806 1041 1809 1068
rect 1826 1058 1830 1061
rect 1814 1052 1817 1058
rect 1826 1048 1830 1051
rect 1806 1038 1817 1041
rect 1718 952 1721 1018
rect 1774 982 1777 1018
rect 1682 948 1686 951
rect 1650 928 1654 931
rect 1526 882 1529 918
rect 1574 892 1577 928
rect 1558 872 1561 878
rect 1590 872 1593 878
rect 1526 863 1529 868
rect 1526 792 1529 838
rect 1558 752 1561 868
rect 1598 862 1601 888
rect 1646 882 1649 918
rect 1626 878 1630 881
rect 1610 868 1614 871
rect 1610 858 1614 861
rect 1586 848 1590 851
rect 1600 803 1602 807
rect 1606 803 1609 807
rect 1613 803 1616 807
rect 1614 752 1617 758
rect 1606 742 1609 748
rect 1502 738 1510 741
rect 1578 738 1582 741
rect 1438 692 1441 708
rect 1446 682 1449 688
rect 1398 678 1425 681
rect 1398 672 1401 678
rect 1422 672 1425 678
rect 1410 668 1414 671
rect 1450 668 1454 671
rect 1402 658 1406 661
rect 1458 658 1462 661
rect 1422 592 1425 658
rect 1478 642 1481 648
rect 1486 592 1489 658
rect 1442 588 1446 591
rect 1454 572 1457 578
rect 1442 568 1446 571
rect 1478 562 1481 568
rect 1294 472 1297 528
rect 1310 472 1313 558
rect 1462 552 1465 558
rect 1322 548 1326 551
rect 1342 542 1345 548
rect 1378 547 1382 550
rect 1406 542 1409 548
rect 1330 538 1334 541
rect 1318 532 1321 538
rect 1338 528 1342 531
rect 1438 482 1441 548
rect 1470 482 1473 558
rect 1486 552 1489 558
rect 1502 472 1505 738
rect 1510 682 1513 688
rect 1526 672 1529 718
rect 1510 662 1513 668
rect 1550 662 1553 668
rect 1558 652 1561 658
rect 1514 638 1518 641
rect 1526 531 1529 548
rect 1522 528 1529 531
rect 1306 468 1310 471
rect 1406 462 1409 468
rect 1314 458 1318 461
rect 1302 452 1305 458
rect 1334 452 1337 458
rect 1438 452 1441 459
rect 1250 448 1254 451
rect 1246 392 1249 428
rect 1154 388 1158 391
rect 1190 362 1193 378
rect 1238 372 1241 388
rect 1242 358 1246 361
rect 1194 348 1198 351
rect 1166 332 1169 338
rect 1046 272 1049 278
rect 1054 272 1057 308
rect 782 252 785 258
rect 862 252 865 258
rect 894 252 897 259
rect 950 252 953 258
rect 782 232 785 248
rect 934 242 937 248
rect 782 192 785 228
rect 854 192 857 218
rect 894 192 897 208
rect 918 192 921 228
rect 942 192 945 248
rect 974 222 977 258
rect 982 232 985 268
rect 1006 222 1009 268
rect 1018 248 1022 251
rect 638 82 641 88
rect 638 62 641 78
rect 646 72 649 98
rect 742 92 745 118
rect 674 88 678 91
rect 750 72 753 78
rect 694 62 697 68
rect 702 62 705 68
rect 766 62 769 128
rect 782 82 785 138
rect 774 72 777 78
rect 798 72 801 78
rect 782 62 785 68
rect 806 62 809 128
rect 822 92 825 158
rect 838 142 841 168
rect 906 158 910 161
rect 870 152 873 158
rect 922 148 926 151
rect 938 148 942 151
rect 846 142 849 148
rect 822 62 825 68
rect 438 52 441 59
rect 818 58 822 61
rect 830 52 833 68
rect 838 62 841 78
rect 846 72 849 128
rect 862 102 865 128
rect 870 112 873 148
rect 950 142 953 148
rect 882 138 886 141
rect 898 128 902 131
rect 946 128 950 131
rect 886 82 889 118
rect 894 92 897 98
rect 926 92 929 128
rect 910 72 913 88
rect 918 72 921 78
rect 942 72 945 88
rect 858 68 862 71
rect 862 52 865 58
rect 870 52 873 58
rect 894 52 897 58
rect 934 52 937 68
rect 946 58 950 61
rect 958 52 961 158
rect 1026 138 1030 141
rect 982 132 985 138
rect 998 132 1001 138
rect 1010 128 1014 131
rect 982 92 985 108
rect 1038 82 1041 268
rect 1054 262 1057 268
rect 1062 252 1065 318
rect 1080 303 1082 307
rect 1086 303 1089 307
rect 1093 303 1096 307
rect 1174 292 1177 348
rect 1206 342 1209 358
rect 1218 348 1222 351
rect 1234 348 1241 351
rect 1194 338 1198 341
rect 1218 338 1222 341
rect 1222 332 1225 338
rect 1238 292 1241 348
rect 1246 342 1249 348
rect 1218 288 1222 291
rect 1086 282 1089 288
rect 1114 278 1118 281
rect 1226 278 1230 281
rect 1078 262 1081 278
rect 1106 268 1110 271
rect 1070 252 1073 258
rect 1150 252 1153 259
rect 1182 252 1185 258
rect 1118 242 1121 248
rect 1098 158 1102 161
rect 1182 152 1185 158
rect 1162 148 1166 151
rect 1118 142 1121 148
rect 1054 132 1057 138
rect 1046 112 1049 128
rect 1110 122 1113 138
rect 1158 132 1161 138
rect 1190 132 1193 218
rect 1222 152 1225 158
rect 1226 138 1230 141
rect 1246 132 1249 338
rect 1254 272 1257 308
rect 1262 282 1265 288
rect 1278 282 1281 448
rect 1350 442 1353 448
rect 1534 442 1537 548
rect 1542 542 1545 558
rect 1566 542 1569 698
rect 1622 672 1625 748
rect 1638 742 1641 748
rect 1646 742 1649 868
rect 1654 862 1657 888
rect 1666 878 1670 881
rect 1670 762 1673 878
rect 1686 752 1689 948
rect 1698 938 1702 941
rect 1694 892 1697 918
rect 1710 871 1713 948
rect 1718 942 1721 948
rect 1750 942 1753 968
rect 1774 942 1777 948
rect 1730 928 1734 931
rect 1726 902 1729 918
rect 1750 882 1753 938
rect 1814 932 1817 1038
rect 1830 952 1833 968
rect 1838 942 1841 1098
rect 1846 1092 1849 1528
rect 1854 1482 1857 1488
rect 1862 1482 1865 1488
rect 1858 1468 1862 1471
rect 1854 1262 1857 1348
rect 1862 1292 1865 1418
rect 1870 1402 1873 1538
rect 1894 1522 1897 1548
rect 1878 1462 1881 1498
rect 1886 1462 1889 1468
rect 1894 1452 1897 1458
rect 1878 1442 1881 1448
rect 1902 1352 1905 1538
rect 1926 1532 1929 1548
rect 1934 1542 1937 1548
rect 2030 1542 2033 1638
rect 2046 1542 2049 1547
rect 1978 1538 1982 1541
rect 1994 1538 1998 1541
rect 1986 1528 1990 1531
rect 1918 1482 1921 1518
rect 1910 1462 1913 1468
rect 1918 1462 1921 1478
rect 1934 1472 1937 1508
rect 1978 1488 1982 1491
rect 1934 1462 1937 1468
rect 1962 1458 1966 1461
rect 1910 1442 1913 1448
rect 1882 1348 1886 1351
rect 1858 1248 1862 1251
rect 1854 1072 1857 1118
rect 1870 1112 1873 1318
rect 1890 1268 1894 1271
rect 1902 1251 1905 1318
rect 1918 1312 1921 1458
rect 1942 1452 1945 1458
rect 1930 1428 1934 1431
rect 2014 1412 2017 1538
rect 2030 1472 2033 1538
rect 2054 1532 2057 1678
rect 2094 1671 2097 1678
rect 2142 1672 2145 1698
rect 2174 1672 2177 1738
rect 2190 1722 2193 1728
rect 2206 1722 2209 1748
rect 2222 1742 2225 1748
rect 2278 1742 2281 1748
rect 2314 1747 2318 1750
rect 2382 1742 2385 1758
rect 2398 1752 2401 1758
rect 2430 1742 2433 1748
rect 2470 1742 2473 1748
rect 2502 1744 2505 1778
rect 2666 1758 2670 1761
rect 2234 1738 2238 1741
rect 2258 1738 2262 1741
rect 2386 1738 2390 1741
rect 2490 1738 2494 1741
rect 2246 1722 2249 1738
rect 2274 1728 2278 1731
rect 2182 1682 2185 1688
rect 2090 1668 2097 1671
rect 2170 1668 2174 1671
rect 2102 1662 2105 1668
rect 2182 1662 2185 1678
rect 2082 1658 2086 1661
rect 2146 1658 2150 1661
rect 2102 1612 2105 1658
rect 2154 1648 2158 1651
rect 2190 1622 2193 1718
rect 2206 1692 2209 1698
rect 2222 1672 2225 1718
rect 2230 1672 2233 1688
rect 2270 1682 2273 1688
rect 2294 1682 2297 1738
rect 2406 1732 2409 1738
rect 2422 1732 2425 1738
rect 2458 1728 2462 1731
rect 2430 1722 2433 1728
rect 2394 1718 2398 1721
rect 2458 1718 2462 1721
rect 2470 1692 2473 1738
rect 2502 1732 2505 1740
rect 2490 1728 2494 1731
rect 2478 1692 2481 1718
rect 2354 1688 2358 1691
rect 2402 1688 2406 1691
rect 2390 1672 2393 1688
rect 2454 1672 2457 1688
rect 2290 1668 2294 1671
rect 2322 1668 2326 1671
rect 2450 1668 2454 1671
rect 2466 1668 2473 1671
rect 2198 1632 2201 1658
rect 2114 1578 2118 1581
rect 2178 1568 2182 1571
rect 2198 1562 2201 1618
rect 2222 1592 2225 1668
rect 2230 1652 2233 1668
rect 2270 1662 2273 1668
rect 2358 1662 2361 1668
rect 2366 1662 2369 1668
rect 2278 1652 2281 1658
rect 2246 1622 2249 1648
rect 2294 1622 2297 1658
rect 2302 1652 2305 1658
rect 2310 1652 2313 1658
rect 2146 1548 2150 1551
rect 2070 1482 2073 1528
rect 2134 1522 2137 1528
rect 2104 1503 2106 1507
rect 2110 1503 2113 1507
rect 2117 1503 2120 1507
rect 2142 1492 2145 1548
rect 2158 1542 2161 1558
rect 2198 1552 2201 1558
rect 2214 1552 2217 1558
rect 2222 1552 2225 1568
rect 2182 1542 2185 1548
rect 2190 1542 2193 1548
rect 2210 1538 2214 1541
rect 2230 1541 2233 1598
rect 2278 1552 2281 1558
rect 2294 1552 2297 1608
rect 2310 1592 2313 1618
rect 2334 1592 2337 1658
rect 2346 1648 2350 1651
rect 2358 1642 2361 1658
rect 2398 1652 2401 1658
rect 2370 1648 2374 1651
rect 2382 1642 2385 1648
rect 2226 1538 2233 1541
rect 2162 1528 2166 1531
rect 2254 1528 2262 1531
rect 2246 1502 2249 1518
rect 2082 1478 2086 1481
rect 2038 1463 2041 1478
rect 2118 1472 2121 1478
rect 2130 1468 2134 1471
rect 2142 1462 2145 1468
rect 2090 1458 2094 1461
rect 2166 1452 2169 1478
rect 2182 1472 2185 1498
rect 2230 1472 2233 1488
rect 2254 1472 2257 1528
rect 2270 1522 2273 1548
rect 2290 1528 2294 1531
rect 2262 1482 2265 1488
rect 2234 1458 2238 1461
rect 2206 1452 2209 1458
rect 2102 1432 2105 1448
rect 2022 1392 2025 1398
rect 1954 1378 1958 1381
rect 1986 1368 1990 1371
rect 2002 1368 2006 1371
rect 1942 1352 1945 1368
rect 2014 1362 2017 1378
rect 2062 1362 2065 1368
rect 2078 1362 2081 1388
rect 1962 1358 1966 1361
rect 1962 1348 1966 1351
rect 1942 1342 1945 1348
rect 1974 1342 1977 1348
rect 1982 1342 1985 1348
rect 2030 1342 2033 1348
rect 1930 1338 1934 1341
rect 1910 1292 1913 1308
rect 1934 1292 1937 1338
rect 1942 1312 1945 1328
rect 1918 1272 1921 1278
rect 1938 1258 1942 1261
rect 1950 1252 1953 1278
rect 1974 1262 1977 1338
rect 2038 1332 2041 1358
rect 2010 1328 2014 1331
rect 1902 1248 1913 1251
rect 1898 1238 1902 1241
rect 1910 1172 1913 1248
rect 1930 1238 1934 1241
rect 1990 1221 1993 1258
rect 2022 1252 2025 1259
rect 1982 1218 1993 1221
rect 1942 1162 1945 1218
rect 1918 1142 1921 1158
rect 1934 1132 1937 1147
rect 1898 1118 1902 1121
rect 1918 1092 1921 1128
rect 1910 1082 1913 1088
rect 1926 1072 1929 1078
rect 1942 1072 1945 1158
rect 1958 1152 1961 1218
rect 1982 1172 1985 1218
rect 2006 1142 2009 1148
rect 1906 1068 1910 1071
rect 1838 912 1841 938
rect 1718 872 1721 878
rect 1710 868 1718 871
rect 1702 852 1705 858
rect 1734 752 1737 868
rect 1758 862 1761 898
rect 1798 852 1801 908
rect 1814 882 1817 888
rect 1822 882 1825 888
rect 1830 882 1833 888
rect 1846 881 1849 1058
rect 1934 1052 1937 1058
rect 1882 1038 1886 1041
rect 1854 962 1857 968
rect 1862 942 1865 978
rect 1870 962 1873 968
rect 1854 912 1857 918
rect 1862 892 1865 928
rect 1870 902 1873 948
rect 1842 878 1849 881
rect 1814 862 1817 878
rect 1878 872 1881 888
rect 1886 882 1889 908
rect 1894 892 1897 938
rect 1902 932 1905 948
rect 1902 872 1905 888
rect 1918 872 1921 978
rect 1934 882 1937 898
rect 1942 872 1945 1068
rect 1954 1058 1958 1061
rect 1954 1048 1958 1051
rect 1966 952 1969 1138
rect 2038 1132 2041 1328
rect 2054 1282 2057 1328
rect 2062 1292 2065 1348
rect 2086 1332 2089 1338
rect 2074 1328 2078 1331
rect 2094 1291 2097 1348
rect 2102 1342 2105 1368
rect 2142 1342 2145 1418
rect 2166 1392 2169 1438
rect 2190 1382 2193 1388
rect 2198 1372 2201 1418
rect 2214 1392 2217 1458
rect 2222 1451 2225 1458
rect 2222 1448 2233 1451
rect 2230 1392 2233 1448
rect 2238 1442 2241 1448
rect 2270 1442 2273 1518
rect 2286 1492 2289 1528
rect 2326 1492 2329 1528
rect 2302 1482 2305 1488
rect 2290 1468 2294 1471
rect 2302 1461 2305 1478
rect 2334 1462 2337 1468
rect 2294 1458 2305 1461
rect 2314 1458 2318 1461
rect 2278 1452 2281 1458
rect 2286 1452 2289 1458
rect 2278 1392 2281 1438
rect 2286 1362 2289 1368
rect 2274 1358 2281 1361
rect 2174 1352 2177 1358
rect 2198 1352 2201 1358
rect 2150 1332 2153 1348
rect 2198 1342 2201 1348
rect 2122 1328 2126 1331
rect 2134 1322 2137 1328
rect 2104 1303 2106 1307
rect 2110 1303 2113 1307
rect 2117 1303 2120 1307
rect 2094 1288 2105 1291
rect 2078 1272 2081 1278
rect 2090 1268 2094 1271
rect 2070 1242 2073 1258
rect 2086 1252 2089 1258
rect 2102 1212 2105 1288
rect 2146 1278 2150 1281
rect 2110 1272 2113 1278
rect 2158 1271 2161 1338
rect 2182 1312 2185 1338
rect 2170 1278 2174 1281
rect 2154 1268 2161 1271
rect 2182 1271 2185 1308
rect 2178 1268 2185 1271
rect 2122 1258 2126 1261
rect 2162 1258 2166 1261
rect 2190 1261 2193 1328
rect 2206 1282 2209 1348
rect 2222 1332 2225 1358
rect 2246 1342 2249 1348
rect 2266 1338 2270 1341
rect 2222 1272 2225 1328
rect 2238 1282 2241 1328
rect 2258 1318 2262 1321
rect 2230 1262 2233 1278
rect 2270 1272 2273 1338
rect 2278 1331 2281 1358
rect 2286 1342 2289 1358
rect 2278 1328 2286 1331
rect 2254 1262 2257 1268
rect 2278 1262 2281 1318
rect 2286 1292 2289 1328
rect 2186 1258 2193 1261
rect 2142 1252 2145 1258
rect 2198 1242 2201 1258
rect 2222 1242 2225 1258
rect 2246 1252 2249 1258
rect 2266 1248 2270 1251
rect 2134 1192 2137 1218
rect 2166 1192 2169 1238
rect 2238 1192 2241 1208
rect 2222 1162 2225 1168
rect 2142 1158 2150 1161
rect 2046 1152 2049 1158
rect 2122 1148 2126 1151
rect 1998 1112 2001 1118
rect 1974 1072 1977 1108
rect 2014 1092 2017 1118
rect 2046 1092 2049 1118
rect 2022 1072 2025 1078
rect 2030 1072 2033 1078
rect 2006 1042 2009 1048
rect 2038 992 2041 1078
rect 2054 1072 2057 1078
rect 2046 1052 2049 1068
rect 2062 1062 2065 1128
rect 2070 1102 2073 1118
rect 2078 1092 2081 1148
rect 2098 1138 2105 1141
rect 2094 1122 2097 1128
rect 2102 1122 2105 1138
rect 2104 1103 2106 1107
rect 2110 1103 2113 1107
rect 2117 1103 2120 1107
rect 2086 1082 2089 1088
rect 2002 988 2006 991
rect 2038 962 2041 988
rect 2046 962 2049 1048
rect 2062 972 2065 1058
rect 2070 1042 2073 1068
rect 2086 1051 2089 1078
rect 2142 1072 2145 1158
rect 2182 1152 2185 1158
rect 2214 1142 2217 1148
rect 2158 1132 2161 1138
rect 2186 1128 2190 1131
rect 2210 1128 2214 1131
rect 2214 1082 2217 1088
rect 2222 1082 2225 1108
rect 2230 1092 2233 1138
rect 2238 1092 2241 1148
rect 2246 1142 2249 1148
rect 2254 1142 2257 1148
rect 2286 1142 2289 1268
rect 2294 1182 2297 1458
rect 2342 1452 2345 1548
rect 2350 1542 2353 1578
rect 2406 1561 2409 1668
rect 2470 1662 2473 1668
rect 2518 1671 2521 1718
rect 2526 1712 2529 1748
rect 2542 1732 2545 1758
rect 2550 1742 2553 1748
rect 2590 1742 2593 1747
rect 2554 1728 2558 1731
rect 2558 1692 2561 1718
rect 2518 1668 2526 1671
rect 2494 1662 2497 1668
rect 2534 1662 2537 1688
rect 2574 1682 2577 1738
rect 2670 1732 2673 1748
rect 2654 1722 2657 1728
rect 2450 1658 2454 1661
rect 2482 1658 2486 1661
rect 2414 1652 2417 1658
rect 2414 1592 2417 1638
rect 2462 1622 2465 1658
rect 2478 1648 2486 1651
rect 2438 1592 2441 1618
rect 2478 1592 2481 1648
rect 2518 1612 2521 1658
rect 2398 1558 2409 1561
rect 2366 1552 2369 1558
rect 2398 1542 2401 1558
rect 2382 1508 2390 1511
rect 2358 1492 2361 1498
rect 2382 1492 2385 1508
rect 2390 1482 2393 1498
rect 2398 1472 2401 1478
rect 2406 1462 2409 1548
rect 2430 1532 2433 1548
rect 2462 1542 2465 1548
rect 2478 1532 2481 1578
rect 2494 1562 2497 1568
rect 2542 1562 2545 1658
rect 2550 1642 2553 1648
rect 2558 1631 2561 1678
rect 2574 1662 2577 1668
rect 2590 1642 2593 1678
rect 2606 1672 2609 1718
rect 2638 1692 2641 1698
rect 2670 1672 2673 1688
rect 2550 1628 2561 1631
rect 2550 1592 2553 1628
rect 2558 1602 2561 1618
rect 2562 1558 2566 1561
rect 2534 1552 2537 1558
rect 2574 1552 2577 1558
rect 2546 1548 2550 1551
rect 2422 1502 2425 1528
rect 2446 1502 2449 1528
rect 2478 1492 2481 1528
rect 2486 1492 2489 1528
rect 2502 1522 2505 1548
rect 2526 1532 2529 1538
rect 2510 1522 2513 1528
rect 2518 1512 2521 1518
rect 2494 1481 2497 1498
rect 2490 1478 2497 1481
rect 2430 1472 2433 1478
rect 2446 1462 2449 1468
rect 2426 1458 2430 1461
rect 2302 1392 2305 1448
rect 2374 1442 2377 1458
rect 2378 1378 2382 1381
rect 2346 1368 2350 1371
rect 2334 1362 2337 1368
rect 2322 1358 2326 1361
rect 2310 1332 2313 1358
rect 2334 1342 2337 1358
rect 2358 1352 2361 1358
rect 2390 1351 2393 1458
rect 2402 1448 2406 1451
rect 2414 1392 2417 1458
rect 2434 1448 2438 1451
rect 2458 1438 2462 1441
rect 2446 1422 2449 1428
rect 2422 1392 2425 1408
rect 2386 1348 2393 1351
rect 2406 1352 2409 1358
rect 2414 1352 2417 1368
rect 2322 1338 2326 1341
rect 2370 1328 2374 1331
rect 2302 1272 2305 1318
rect 2310 1162 2313 1328
rect 2382 1322 2385 1348
rect 2318 1292 2321 1298
rect 2326 1272 2329 1288
rect 2350 1282 2353 1288
rect 2334 1262 2337 1268
rect 2342 1212 2345 1218
rect 2350 1172 2353 1278
rect 2358 1242 2361 1278
rect 2382 1272 2385 1278
rect 2370 1258 2374 1261
rect 2382 1242 2385 1248
rect 2390 1232 2393 1328
rect 2398 1312 2401 1318
rect 2402 1258 2406 1261
rect 2406 1232 2409 1238
rect 2298 1158 2302 1161
rect 2370 1158 2374 1161
rect 2302 1152 2305 1158
rect 2310 1142 2313 1148
rect 2350 1142 2353 1148
rect 2358 1142 2361 1148
rect 2374 1142 2377 1158
rect 2262 1132 2265 1140
rect 2158 1072 2161 1078
rect 2098 1068 2102 1071
rect 2166 1062 2169 1078
rect 2182 1072 2185 1078
rect 2250 1068 2254 1071
rect 2082 1048 2089 1051
rect 2114 1058 2118 1061
rect 2154 1058 2158 1061
rect 2202 1058 2206 1061
rect 2262 1061 2265 1068
rect 2258 1058 2265 1061
rect 2270 1062 2273 1068
rect 2094 1051 2097 1058
rect 2174 1052 2177 1058
rect 2094 1048 2118 1051
rect 2222 992 2225 1058
rect 2230 1042 2233 1048
rect 2254 992 2257 1058
rect 2054 952 2057 968
rect 2090 958 2094 961
rect 1950 922 1953 948
rect 1966 912 1969 948
rect 2006 932 2009 938
rect 2022 932 2025 938
rect 2014 922 2017 928
rect 1982 882 1985 888
rect 2006 882 2009 898
rect 1974 872 1977 878
rect 1846 852 1849 868
rect 1854 862 1857 868
rect 1918 862 1921 868
rect 1990 862 1993 878
rect 2006 862 2009 878
rect 2018 868 2022 871
rect 1954 858 1958 861
rect 1962 848 1966 851
rect 1798 802 1801 848
rect 1710 732 1713 748
rect 1666 728 1670 731
rect 1614 621 1617 668
rect 1614 618 1625 621
rect 1590 592 1593 618
rect 1600 603 1602 607
rect 1606 603 1609 607
rect 1613 603 1616 607
rect 1590 562 1593 588
rect 1622 552 1625 618
rect 1630 602 1633 718
rect 1638 551 1641 618
rect 1562 528 1566 531
rect 1550 462 1553 518
rect 1574 502 1577 548
rect 1622 542 1625 548
rect 1582 532 1585 538
rect 1598 492 1601 498
rect 1390 362 1393 368
rect 1398 352 1401 358
rect 1378 348 1382 351
rect 1454 351 1457 368
rect 1294 342 1297 347
rect 1290 288 1294 291
rect 1258 258 1262 261
rect 1282 258 1286 261
rect 1302 252 1305 298
rect 1310 282 1313 288
rect 1318 282 1321 308
rect 1326 302 1329 348
rect 1542 342 1545 358
rect 1558 352 1561 458
rect 1570 358 1574 361
rect 1410 338 1414 341
rect 1330 288 1334 291
rect 1314 268 1318 271
rect 1342 262 1345 338
rect 1366 332 1369 338
rect 1418 328 1422 331
rect 1358 312 1361 318
rect 1390 282 1393 328
rect 1454 302 1457 328
rect 1518 322 1521 338
rect 1526 312 1529 338
rect 1582 332 1585 448
rect 1634 418 1638 421
rect 1600 403 1602 407
rect 1606 403 1609 407
rect 1613 403 1616 407
rect 1646 372 1649 718
rect 1658 678 1662 681
rect 1654 482 1657 588
rect 1662 542 1665 678
rect 1670 552 1673 728
rect 1694 662 1697 708
rect 1734 682 1737 738
rect 1774 722 1777 758
rect 1798 742 1801 798
rect 1814 772 1817 818
rect 1834 768 1838 771
rect 1846 752 1849 848
rect 1990 842 1993 858
rect 1998 842 2001 848
rect 1946 838 1950 841
rect 1950 822 1953 838
rect 1958 832 1961 838
rect 1854 762 1857 768
rect 1886 762 1889 808
rect 1814 742 1817 748
rect 1782 732 1785 738
rect 1794 728 1798 731
rect 1762 718 1766 721
rect 1750 682 1753 718
rect 1738 678 1742 681
rect 1766 672 1769 678
rect 1754 668 1758 671
rect 1678 592 1681 618
rect 1706 538 1710 541
rect 1662 492 1665 538
rect 1702 512 1705 518
rect 1718 482 1721 618
rect 1726 562 1729 658
rect 1774 651 1777 718
rect 1786 668 1790 671
rect 1806 671 1809 718
rect 1822 712 1825 748
rect 1862 742 1865 748
rect 1898 738 1902 741
rect 1846 732 1849 738
rect 1862 682 1865 738
rect 1910 732 1913 768
rect 1942 762 1945 768
rect 1918 742 1921 748
rect 1934 742 1937 748
rect 1958 742 1961 748
rect 1990 742 1993 808
rect 2014 781 2017 868
rect 2006 778 2017 781
rect 2006 752 2009 778
rect 2014 762 2017 768
rect 1870 722 1873 728
rect 1838 672 1841 678
rect 1806 668 1817 671
rect 1858 668 1862 671
rect 1878 671 1881 728
rect 1910 702 1913 728
rect 1918 672 1921 738
rect 1998 732 2001 748
rect 2022 742 2025 858
rect 2030 762 2033 858
rect 2054 852 2057 948
rect 2070 942 2073 948
rect 2094 942 2097 948
rect 2062 882 2065 938
rect 2070 882 2073 938
rect 2110 932 2113 968
rect 2158 942 2161 948
rect 2206 942 2209 988
rect 2238 952 2241 978
rect 2254 962 2257 988
rect 2278 962 2281 1118
rect 2318 1112 2321 1118
rect 2290 1088 2294 1091
rect 2302 1082 2305 1088
rect 2326 1082 2329 1128
rect 2342 1102 2345 1118
rect 2322 1078 2326 1081
rect 2346 1078 2350 1081
rect 2366 1062 2369 1118
rect 2382 1101 2385 1228
rect 2390 1132 2393 1148
rect 2414 1142 2417 1148
rect 2422 1131 2425 1388
rect 2470 1372 2473 1458
rect 2502 1451 2505 1508
rect 2534 1492 2537 1548
rect 2590 1542 2593 1588
rect 2614 1582 2617 1658
rect 2542 1502 2545 1538
rect 2590 1532 2593 1538
rect 2610 1528 2614 1531
rect 2622 1522 2625 1668
rect 2678 1612 2681 1658
rect 2694 1562 2697 1618
rect 2642 1558 2646 1561
rect 2638 1502 2641 1558
rect 2650 1538 2654 1541
rect 2682 1538 2686 1541
rect 2678 1528 2686 1531
rect 2510 1462 2513 1488
rect 2586 1478 2590 1481
rect 2530 1468 2534 1471
rect 2574 1470 2577 1478
rect 2518 1452 2521 1468
rect 2542 1462 2545 1468
rect 2582 1462 2585 1468
rect 2590 1462 2593 1468
rect 2614 1462 2617 1498
rect 2638 1472 2641 1488
rect 2662 1481 2665 1518
rect 2662 1478 2673 1481
rect 2646 1472 2649 1478
rect 2630 1462 2633 1468
rect 2650 1458 2654 1461
rect 2526 1452 2529 1458
rect 2498 1448 2505 1451
rect 2510 1442 2513 1448
rect 2550 1392 2553 1448
rect 2458 1358 2462 1361
rect 2478 1352 2481 1368
rect 2494 1362 2497 1368
rect 2510 1352 2513 1358
rect 2550 1352 2553 1378
rect 2566 1362 2569 1398
rect 2582 1362 2585 1458
rect 2614 1422 2617 1448
rect 2622 1402 2625 1458
rect 2662 1392 2665 1468
rect 2590 1372 2593 1378
rect 2458 1348 2462 1351
rect 2498 1348 2502 1351
rect 2522 1348 2526 1351
rect 2462 1332 2465 1338
rect 2430 1292 2433 1328
rect 2454 1292 2457 1318
rect 2470 1282 2473 1338
rect 2478 1282 2481 1338
rect 2430 1252 2433 1278
rect 2450 1258 2454 1261
rect 2430 1242 2433 1248
rect 2438 1242 2441 1248
rect 2478 1201 2481 1278
rect 2486 1262 2489 1348
rect 2534 1342 2537 1348
rect 2502 1322 2505 1338
rect 2542 1332 2545 1338
rect 2526 1322 2529 1328
rect 2534 1282 2537 1288
rect 2550 1282 2553 1308
rect 2566 1292 2569 1338
rect 2574 1312 2577 1358
rect 2606 1352 2609 1358
rect 2662 1352 2665 1358
rect 2590 1332 2593 1348
rect 2598 1342 2601 1348
rect 2622 1342 2625 1348
rect 2606 1332 2609 1338
rect 2646 1332 2649 1348
rect 2658 1338 2662 1341
rect 2626 1328 2630 1331
rect 2558 1282 2561 1288
rect 2494 1278 2502 1281
rect 2494 1272 2497 1278
rect 2574 1272 2577 1298
rect 2622 1292 2625 1298
rect 2598 1282 2601 1288
rect 2634 1278 2638 1281
rect 2490 1258 2494 1261
rect 2510 1232 2513 1268
rect 2582 1252 2585 1258
rect 2590 1212 2593 1278
rect 2618 1268 2622 1271
rect 2478 1198 2486 1201
rect 2430 1162 2433 1198
rect 2646 1192 2649 1268
rect 2662 1262 2665 1338
rect 2670 1272 2673 1478
rect 2678 1392 2681 1528
rect 2690 1488 2694 1491
rect 2702 1482 2705 1488
rect 2686 1472 2689 1478
rect 2686 1452 2689 1458
rect 2682 1338 2686 1341
rect 2698 1268 2702 1271
rect 2662 1251 2665 1258
rect 2662 1248 2670 1251
rect 2474 1158 2478 1161
rect 2482 1148 2486 1151
rect 2462 1142 2465 1148
rect 2478 1142 2481 1148
rect 2510 1142 2513 1148
rect 2414 1128 2425 1131
rect 2454 1132 2457 1138
rect 2502 1132 2505 1138
rect 2526 1132 2529 1178
rect 2534 1152 2537 1158
rect 2542 1152 2545 1158
rect 2550 1132 2553 1188
rect 2558 1152 2561 1168
rect 2670 1162 2673 1248
rect 2582 1152 2585 1158
rect 2630 1152 2633 1158
rect 2662 1142 2665 1158
rect 2702 1142 2705 1148
rect 2578 1138 2582 1141
rect 2602 1138 2606 1141
rect 2626 1138 2630 1141
rect 2642 1138 2649 1141
rect 2570 1128 2574 1131
rect 2382 1098 2393 1101
rect 2390 1082 2393 1098
rect 2314 1058 2318 1061
rect 2322 1058 2329 1061
rect 2218 948 2222 951
rect 2130 928 2134 931
rect 2150 922 2153 938
rect 2086 882 2089 918
rect 2104 903 2106 907
rect 2110 903 2113 907
rect 2117 903 2120 907
rect 2066 868 2070 871
rect 2074 858 2078 861
rect 2130 858 2134 861
rect 2038 832 2041 848
rect 2046 842 2049 848
rect 2046 742 2049 798
rect 2054 772 2057 818
rect 2086 812 2089 848
rect 2078 752 2081 758
rect 2058 748 2062 751
rect 2074 738 2078 741
rect 2022 732 2025 738
rect 2034 728 2038 731
rect 2050 728 2054 731
rect 1942 692 1945 718
rect 1958 692 1961 708
rect 1998 701 2001 728
rect 1990 698 2001 701
rect 2022 702 2025 718
rect 1990 672 1993 698
rect 1874 668 1881 671
rect 1938 668 1942 671
rect 1770 648 1777 651
rect 1802 658 1806 661
rect 1782 641 1785 658
rect 1774 638 1785 641
rect 1774 592 1777 638
rect 1806 572 1809 618
rect 1758 552 1761 568
rect 1794 558 1798 561
rect 1814 552 1817 668
rect 1902 662 1905 668
rect 1858 658 1862 661
rect 1890 658 1894 661
rect 1922 658 1926 661
rect 1910 572 1913 618
rect 1926 592 1929 598
rect 1934 592 1937 658
rect 1942 592 1945 668
rect 1990 662 1993 668
rect 2006 661 2009 679
rect 2022 672 2025 698
rect 2038 692 2041 708
rect 2062 702 2065 738
rect 2054 682 2057 688
rect 2062 672 2065 698
rect 2086 692 2089 808
rect 2094 762 2097 858
rect 2150 852 2153 898
rect 2130 747 2134 750
rect 2110 732 2113 738
rect 2158 732 2161 938
rect 2178 918 2182 921
rect 2194 878 2198 881
rect 2214 872 2217 948
rect 2302 942 2305 998
rect 2310 962 2313 968
rect 2326 952 2329 1058
rect 2346 1058 2350 1061
rect 2334 1052 2337 1058
rect 2398 1031 2401 1038
rect 2406 1031 2409 1118
rect 2398 1028 2409 1031
rect 2414 1072 2417 1128
rect 2426 1118 2430 1121
rect 2438 1112 2441 1118
rect 2430 1092 2433 1108
rect 2462 1072 2465 1108
rect 2358 962 2361 1018
rect 2398 962 2401 1028
rect 2406 962 2409 1018
rect 2414 952 2417 1068
rect 2470 1062 2473 1118
rect 2486 1082 2489 1088
rect 2478 1052 2481 1058
rect 2494 1051 2497 1118
rect 2486 1048 2497 1051
rect 2438 952 2441 1008
rect 2330 938 2334 941
rect 2354 938 2358 941
rect 2378 938 2382 941
rect 2382 932 2385 938
rect 2390 932 2393 938
rect 2234 928 2241 931
rect 2222 862 2225 868
rect 2230 862 2233 868
rect 2178 858 2182 861
rect 2174 742 2177 818
rect 2086 682 2089 688
rect 2006 658 2014 661
rect 2094 661 2097 718
rect 2104 703 2106 707
rect 2110 703 2113 707
rect 2117 703 2120 707
rect 2142 672 2145 678
rect 2182 672 2185 818
rect 2198 792 2201 828
rect 2222 792 2225 858
rect 2238 772 2241 928
rect 2366 922 2369 928
rect 2246 872 2249 878
rect 2254 872 2257 878
rect 2262 862 2265 888
rect 2270 882 2273 918
rect 2294 882 2297 898
rect 2310 882 2313 918
rect 2318 912 2321 918
rect 2374 882 2377 908
rect 2398 892 2401 948
rect 2414 932 2417 938
rect 2462 932 2465 968
rect 2470 932 2473 998
rect 2486 952 2489 1048
rect 2494 1032 2497 1038
rect 2494 952 2497 958
rect 2502 952 2505 968
rect 2486 942 2489 948
rect 2418 928 2422 931
rect 2406 881 2409 918
rect 2430 902 2433 918
rect 2454 892 2457 918
rect 2406 878 2414 881
rect 2318 872 2321 878
rect 2366 872 2369 878
rect 2430 872 2433 888
rect 2274 868 2278 871
rect 2390 862 2393 868
rect 2346 858 2350 861
rect 2294 772 2297 838
rect 2318 792 2321 848
rect 2206 722 2209 728
rect 2194 718 2198 721
rect 2198 692 2201 698
rect 2202 678 2206 681
rect 2222 672 2225 768
rect 2258 748 2262 751
rect 2270 742 2273 748
rect 2234 738 2238 741
rect 2238 712 2241 728
rect 2278 692 2281 758
rect 2294 752 2297 768
rect 2342 762 2345 838
rect 2406 762 2409 868
rect 2450 858 2454 861
rect 2422 792 2425 818
rect 2446 782 2449 858
rect 2454 842 2457 848
rect 2434 758 2438 761
rect 2342 752 2345 758
rect 2322 748 2326 751
rect 2286 712 2289 748
rect 2366 742 2369 748
rect 2306 738 2310 741
rect 2382 741 2385 758
rect 2462 752 2465 878
rect 2478 772 2481 918
rect 2510 912 2513 1068
rect 2518 1062 2521 1118
rect 2526 1092 2529 1128
rect 2598 1112 2601 1128
rect 2558 1072 2561 1098
rect 2646 1092 2649 1138
rect 2678 1081 2681 1118
rect 2702 1082 2705 1138
rect 2678 1078 2686 1081
rect 2606 1072 2609 1078
rect 2638 1072 2641 1078
rect 2618 1068 2622 1071
rect 2526 1051 2529 1068
rect 2662 1062 2665 1068
rect 2554 1058 2558 1061
rect 2518 1048 2529 1051
rect 2610 1048 2614 1051
rect 2518 992 2521 1048
rect 2550 1042 2553 1048
rect 2630 1042 2633 1058
rect 2646 1052 2649 1058
rect 2578 1018 2582 1021
rect 2558 962 2561 988
rect 2642 968 2646 971
rect 2558 952 2561 958
rect 2510 882 2513 888
rect 2534 872 2537 948
rect 2622 942 2625 948
rect 2670 942 2673 1038
rect 2546 928 2550 931
rect 2586 918 2590 921
rect 2654 892 2657 908
rect 2602 888 2606 891
rect 2638 872 2641 888
rect 2670 878 2673 938
rect 2686 902 2689 918
rect 2554 868 2558 871
rect 2582 862 2585 868
rect 2530 858 2534 861
rect 2570 858 2574 861
rect 2486 802 2489 848
rect 2518 792 2521 848
rect 2542 832 2545 848
rect 2526 772 2529 788
rect 2394 748 2398 751
rect 2538 748 2545 751
rect 2406 742 2409 748
rect 2382 738 2390 741
rect 2514 738 2518 741
rect 2374 732 2377 738
rect 2294 692 2297 718
rect 2342 692 2345 708
rect 2234 668 2238 671
rect 2094 658 2102 661
rect 2122 658 2126 661
rect 2138 658 2142 661
rect 2162 658 2166 661
rect 1830 552 1833 568
rect 1862 551 1865 558
rect 2006 552 2009 658
rect 2182 652 2185 668
rect 2246 662 2249 688
rect 2270 672 2273 688
rect 2326 682 2329 688
rect 2374 672 2377 698
rect 2330 668 2334 671
rect 2362 668 2366 671
rect 2198 652 2201 658
rect 2114 638 2118 641
rect 2154 638 2158 641
rect 1730 538 1734 541
rect 1746 538 1750 541
rect 1762 528 1766 531
rect 1734 522 1737 528
rect 1722 459 1726 462
rect 1742 462 1745 518
rect 1766 492 1769 518
rect 1774 492 1777 548
rect 1782 542 1785 548
rect 1802 538 1806 541
rect 1818 538 1822 541
rect 1806 522 1809 528
rect 1758 482 1761 488
rect 1814 462 1817 518
rect 1830 472 1833 538
rect 1894 512 1897 548
rect 1982 512 1985 548
rect 2062 542 2065 548
rect 2050 538 2054 541
rect 1870 472 1873 478
rect 1878 462 1881 508
rect 1694 421 1697 458
rect 1894 452 1897 458
rect 1926 452 1929 459
rect 1686 418 1697 421
rect 1562 318 1566 321
rect 1390 272 1393 278
rect 1406 272 1409 278
rect 1354 268 1358 271
rect 1414 271 1417 288
rect 1410 268 1417 271
rect 1454 272 1457 298
rect 1534 282 1537 288
rect 1574 282 1577 318
rect 1494 272 1497 278
rect 1510 262 1513 278
rect 1530 268 1534 271
rect 1518 262 1521 268
rect 1362 258 1366 261
rect 1590 262 1593 348
rect 1638 342 1641 348
rect 1670 342 1673 347
rect 1686 342 1689 418
rect 1742 392 1745 438
rect 1734 352 1737 358
rect 1758 352 1761 418
rect 1878 362 1881 368
rect 1942 362 1945 478
rect 1958 462 1961 508
rect 1998 492 2001 508
rect 1990 472 1993 488
rect 2046 472 2049 528
rect 2054 522 2057 528
rect 2070 512 2073 548
rect 2102 542 2105 548
rect 2118 532 2121 547
rect 2166 542 2169 618
rect 2182 552 2185 568
rect 2214 551 2217 658
rect 2238 651 2241 658
rect 2270 652 2273 668
rect 2286 652 2289 658
rect 2294 652 2297 658
rect 2238 648 2246 651
rect 2270 591 2273 648
rect 2310 622 2313 658
rect 2294 592 2297 618
rect 2334 592 2337 668
rect 2358 642 2361 658
rect 2366 652 2369 668
rect 2378 658 2382 661
rect 2358 622 2361 638
rect 2270 588 2278 591
rect 2346 588 2350 591
rect 2314 548 2318 551
rect 2286 542 2289 548
rect 2104 503 2106 507
rect 2110 503 2113 507
rect 2117 503 2120 507
rect 2190 492 2193 518
rect 2222 482 2225 538
rect 2390 532 2393 718
rect 2398 652 2401 738
rect 2434 728 2438 731
rect 2406 722 2409 728
rect 2426 718 2430 721
rect 2482 718 2486 721
rect 2438 682 2441 698
rect 2426 678 2430 681
rect 2454 672 2457 678
rect 2478 672 2481 678
rect 2414 662 2417 668
rect 2482 658 2486 661
rect 2398 592 2401 648
rect 2486 632 2489 638
rect 2446 622 2449 628
rect 2430 572 2433 618
rect 2406 551 2409 568
rect 2454 551 2457 558
rect 2454 548 2462 551
rect 2494 542 2497 678
rect 2510 662 2513 668
rect 2518 662 2521 678
rect 2542 672 2545 748
rect 2550 682 2553 758
rect 2558 732 2561 858
rect 2570 848 2574 851
rect 2686 841 2689 868
rect 2678 838 2689 841
rect 2566 752 2569 798
rect 2622 792 2625 828
rect 2574 762 2577 778
rect 2590 752 2593 758
rect 2598 742 2601 778
rect 2606 762 2609 768
rect 2678 762 2681 838
rect 2686 782 2689 788
rect 2674 758 2678 761
rect 2654 752 2657 758
rect 2638 742 2641 748
rect 2566 692 2569 738
rect 2630 732 2633 738
rect 2638 732 2641 738
rect 2590 692 2593 728
rect 2654 712 2657 748
rect 2662 742 2665 748
rect 2686 728 2694 731
rect 2674 718 2678 721
rect 2566 682 2569 688
rect 2574 672 2577 678
rect 2502 652 2505 658
rect 2518 642 2521 658
rect 2526 652 2529 668
rect 2622 592 2625 668
rect 2630 662 2633 668
rect 2614 562 2617 568
rect 2622 561 2625 588
rect 2622 558 2630 561
rect 2634 558 2641 561
rect 2598 552 2601 558
rect 2618 548 2622 551
rect 2450 538 2454 541
rect 2302 522 2305 528
rect 2294 492 2297 508
rect 2390 492 2393 528
rect 2282 488 2286 491
rect 2014 462 2017 468
rect 2062 462 2065 478
rect 2094 462 2097 468
rect 2126 463 2129 468
rect 2034 458 2038 461
rect 2154 458 2158 461
rect 1738 348 1742 351
rect 1814 351 1817 358
rect 1718 342 1721 348
rect 1774 342 1777 348
rect 1798 342 1801 348
rect 1886 342 1889 348
rect 1894 342 1897 358
rect 1918 352 1921 358
rect 1914 338 1918 341
rect 1934 332 1937 338
rect 1914 328 1918 331
rect 1702 322 1705 328
rect 1610 318 1614 321
rect 1470 252 1473 258
rect 1534 252 1537 258
rect 1566 252 1569 259
rect 1362 248 1366 251
rect 1302 142 1305 248
rect 1382 242 1385 248
rect 1370 158 1374 161
rect 1310 151 1313 158
rect 1374 142 1377 148
rect 1382 142 1385 148
rect 1430 142 1433 218
rect 1574 152 1577 158
rect 1474 148 1478 151
rect 1470 142 1473 148
rect 1550 142 1553 148
rect 1482 138 1486 141
rect 1550 132 1553 138
rect 1130 128 1134 131
rect 1242 128 1246 131
rect 1080 103 1082 107
rect 1086 103 1089 107
rect 1093 103 1096 107
rect 1166 102 1169 128
rect 1210 118 1214 121
rect 1054 82 1057 88
rect 1102 82 1105 98
rect 978 78 982 81
rect 1026 78 1030 81
rect 1006 72 1009 78
rect 986 68 990 71
rect 1026 68 1030 71
rect 1038 71 1041 78
rect 1110 72 1113 88
rect 1126 75 1129 98
rect 1174 92 1177 118
rect 1230 92 1233 128
rect 1250 118 1257 121
rect 1158 72 1161 88
rect 1218 78 1222 81
rect 1038 68 1046 71
rect 966 62 969 68
rect 998 62 1001 68
rect 1054 62 1057 68
rect 1010 58 1014 61
rect 1030 52 1033 58
rect 1166 52 1169 78
rect 1182 62 1185 68
rect 1206 62 1209 78
rect 1130 48 1134 51
rect 1174 51 1177 58
rect 1222 52 1225 58
rect 1230 52 1233 78
rect 1246 72 1249 98
rect 1254 92 1257 118
rect 1326 92 1329 118
rect 1342 92 1345 128
rect 1254 72 1257 78
rect 1302 72 1305 88
rect 1366 82 1369 128
rect 1398 82 1401 88
rect 1346 78 1350 81
rect 1318 72 1321 78
rect 1366 72 1369 78
rect 1378 68 1382 71
rect 1310 62 1313 68
rect 1270 52 1273 58
rect 1358 52 1361 58
rect 1382 52 1385 58
rect 1406 52 1409 118
rect 1414 92 1417 118
rect 1438 112 1441 128
rect 1438 91 1441 108
rect 1434 88 1441 91
rect 1422 52 1425 68
rect 1470 62 1473 128
rect 1534 102 1537 118
rect 1510 72 1513 98
rect 1582 92 1585 128
rect 1590 102 1593 258
rect 1614 222 1617 318
rect 1750 302 1753 328
rect 1630 292 1633 298
rect 1654 272 1657 278
rect 1662 262 1665 298
rect 1774 292 1777 328
rect 1678 282 1681 288
rect 1782 282 1785 298
rect 1818 278 1822 281
rect 1600 203 1602 207
rect 1606 203 1609 207
rect 1613 203 1616 207
rect 1622 148 1630 151
rect 1622 132 1625 148
rect 1638 142 1641 258
rect 1674 248 1678 251
rect 1694 192 1697 268
rect 1718 262 1721 268
rect 1814 252 1817 278
rect 1822 262 1825 268
rect 1794 238 1798 241
rect 1694 162 1697 188
rect 1734 152 1737 168
rect 1766 152 1769 158
rect 1862 152 1865 308
rect 1902 272 1905 318
rect 1942 282 1945 358
rect 1958 342 1961 458
rect 2022 392 2025 458
rect 1974 351 1977 368
rect 2038 352 2041 368
rect 2062 362 2065 458
rect 2222 421 2225 459
rect 2214 418 2225 421
rect 2214 392 2217 418
rect 2178 388 2182 391
rect 2046 342 2049 358
rect 2058 348 2062 351
rect 2082 348 2086 351
rect 2118 351 2121 358
rect 1958 321 1961 338
rect 2006 332 2009 338
rect 2102 332 2105 338
rect 2190 332 2193 338
rect 1950 318 1961 321
rect 1950 272 1953 318
rect 2054 292 2057 318
rect 2198 312 2201 348
rect 2246 342 2249 347
rect 2254 342 2257 458
rect 2326 452 2329 458
rect 2294 362 2297 418
rect 2314 388 2318 391
rect 2334 372 2337 488
rect 2422 462 2425 538
rect 2506 528 2510 531
rect 2438 522 2441 528
rect 2550 522 2553 548
rect 2606 542 2609 548
rect 2594 538 2598 541
rect 2574 532 2577 538
rect 2582 532 2585 538
rect 2606 532 2609 538
rect 2638 532 2641 558
rect 2358 452 2361 459
rect 2422 452 2425 458
rect 2318 351 2321 358
rect 2310 348 2321 351
rect 2334 352 2337 368
rect 2310 332 2313 348
rect 2342 342 2345 348
rect 2322 338 2326 341
rect 2104 303 2106 307
rect 2110 303 2113 307
rect 2117 303 2120 307
rect 2158 292 2161 308
rect 2230 292 2233 328
rect 2010 268 2014 271
rect 1878 162 1881 218
rect 1730 148 1734 151
rect 1798 142 1801 147
rect 1634 138 1638 141
rect 1526 72 1529 78
rect 1542 75 1545 88
rect 1630 81 1633 128
rect 1630 78 1641 81
rect 1638 62 1641 78
rect 1646 72 1649 98
rect 1694 82 1697 128
rect 1702 72 1705 88
rect 1702 62 1705 68
rect 1174 48 1182 51
rect 86 42 89 48
rect 222 42 225 48
rect 1542 42 1545 48
rect 46 -22 50 -18
rect 190 -19 193 18
rect 198 -19 202 -18
rect 190 -22 202 -19
rect 358 -19 362 -18
rect 366 -19 369 18
rect 526 12 529 18
rect 550 -18 553 8
rect 576 3 578 7
rect 582 3 585 7
rect 589 3 592 7
rect 838 -18 841 8
rect 1600 3 1602 7
rect 1606 3 1609 7
rect 1613 3 1616 7
rect 358 -22 369 -19
rect 534 -22 538 -18
rect 550 -22 554 -18
rect 598 -22 602 -18
rect 614 -22 618 -18
rect 734 -22 738 -18
rect 758 -22 762 -18
rect 838 -22 842 -18
rect 1238 -22 1242 -18
rect 1486 -22 1490 -18
rect 1566 -22 1570 -18
rect 1710 -19 1713 118
rect 1814 102 1817 138
rect 1830 132 1833 148
rect 1846 142 1849 148
rect 1722 88 1726 91
rect 1758 62 1761 98
rect 1846 82 1849 88
rect 1778 58 1782 61
rect 1718 52 1721 58
rect 1862 52 1865 148
rect 1870 122 1873 148
rect 1886 142 1889 148
rect 1894 131 1897 138
rect 1890 128 1897 131
rect 1882 108 1886 111
rect 1894 92 1897 128
rect 1902 112 1905 140
rect 1918 101 1921 268
rect 1926 262 1929 268
rect 2046 262 2049 288
rect 2078 272 2081 278
rect 2102 272 2105 278
rect 2010 258 2014 261
rect 1930 148 1934 151
rect 1950 142 1953 158
rect 1982 142 1985 158
rect 1994 148 1998 151
rect 1966 132 1969 138
rect 1950 122 1953 128
rect 1914 98 1921 101
rect 1910 82 1913 98
rect 1982 82 1985 138
rect 1942 72 1945 78
rect 1910 63 1913 68
rect 1958 62 1961 68
rect 1982 62 1985 68
rect 2006 62 2009 158
rect 2038 142 2041 258
rect 2070 242 2073 258
rect 2070 192 2073 238
rect 2050 168 2054 171
rect 2086 152 2089 268
rect 2094 252 2097 258
rect 2122 248 2126 251
rect 2110 232 2113 248
rect 2142 242 2145 278
rect 2174 272 2177 278
rect 2206 272 2209 288
rect 2238 282 2241 298
rect 2194 268 2198 271
rect 2150 192 2153 248
rect 2166 242 2169 268
rect 2214 262 2217 268
rect 2094 152 2097 168
rect 2082 148 2086 151
rect 2106 148 2110 151
rect 2054 142 2057 148
rect 2062 142 2065 148
rect 2102 132 2105 138
rect 2134 122 2137 158
rect 2150 152 2153 178
rect 2182 172 2185 178
rect 2104 103 2106 107
rect 2110 103 2113 107
rect 2117 103 2120 107
rect 2038 72 2041 78
rect 2054 72 2057 98
rect 2142 92 2145 138
rect 2150 122 2153 148
rect 2182 142 2185 148
rect 2190 142 2193 258
rect 2246 251 2249 328
rect 2350 322 2353 348
rect 2358 332 2361 338
rect 2254 262 2257 318
rect 2366 312 2369 318
rect 2382 302 2385 358
rect 2390 341 2393 448
rect 2398 352 2401 368
rect 2430 352 2433 468
rect 2454 463 2457 478
rect 2486 462 2489 468
rect 2494 462 2497 488
rect 2502 482 2505 518
rect 2518 492 2521 518
rect 2558 492 2561 518
rect 2566 492 2569 528
rect 2510 482 2513 488
rect 2538 468 2542 471
rect 2510 452 2513 458
rect 2534 452 2537 458
rect 2522 448 2526 451
rect 2502 432 2505 448
rect 2462 352 2465 358
rect 2390 338 2401 341
rect 2398 292 2401 338
rect 2406 302 2409 338
rect 2422 332 2425 338
rect 2414 312 2417 328
rect 2430 321 2433 348
rect 2470 342 2473 348
rect 2458 338 2462 341
rect 2442 328 2446 331
rect 2486 322 2489 338
rect 2426 318 2433 321
rect 2422 292 2425 318
rect 2330 288 2334 291
rect 2290 278 2294 281
rect 2314 278 2318 281
rect 2326 272 2329 278
rect 2374 272 2377 278
rect 2390 272 2393 288
rect 2298 268 2302 271
rect 2262 262 2265 268
rect 2270 262 2273 268
rect 2282 258 2286 261
rect 2246 248 2257 251
rect 2226 168 2230 171
rect 2246 162 2249 188
rect 2226 148 2230 151
rect 2242 148 2246 151
rect 2198 142 2201 148
rect 2158 112 2161 138
rect 2166 132 2169 138
rect 2242 128 2246 131
rect 2214 102 2217 118
rect 2178 88 2182 91
rect 2134 72 2137 88
rect 2166 72 2169 88
rect 2222 72 2225 78
rect 2022 62 2025 68
rect 2238 63 2241 78
rect 2254 72 2257 248
rect 2342 251 2345 268
rect 2370 258 2374 261
rect 2382 252 2385 258
rect 2342 248 2350 251
rect 2370 248 2374 251
rect 2286 241 2289 248
rect 2286 238 2297 241
rect 2282 168 2286 171
rect 2286 142 2289 148
rect 2294 142 2297 238
rect 2310 162 2313 168
rect 2266 138 2270 141
rect 2294 132 2297 138
rect 2270 112 2273 128
rect 2326 101 2329 248
rect 2342 192 2345 228
rect 2350 172 2353 248
rect 2406 172 2409 278
rect 2430 272 2433 298
rect 2446 292 2449 318
rect 2494 312 2497 328
rect 2486 272 2489 278
rect 2502 272 2505 428
rect 2542 382 2545 468
rect 2550 462 2553 488
rect 2570 478 2574 481
rect 2550 361 2553 458
rect 2558 452 2561 468
rect 2590 462 2593 488
rect 2558 402 2561 448
rect 2586 418 2590 421
rect 2550 358 2558 361
rect 2582 352 2585 358
rect 2510 322 2513 348
rect 2542 292 2545 348
rect 2590 342 2593 378
rect 2554 338 2558 341
rect 2566 312 2569 318
rect 2578 288 2582 291
rect 2542 282 2545 288
rect 2590 282 2593 298
rect 2598 292 2601 508
rect 2654 502 2657 708
rect 2678 692 2681 708
rect 2662 662 2665 668
rect 2666 538 2670 541
rect 2674 528 2678 531
rect 2614 432 2617 458
rect 2614 362 2617 398
rect 2646 392 2649 459
rect 2678 452 2681 498
rect 2686 492 2689 728
rect 2694 552 2697 558
rect 2702 482 2705 928
rect 2614 352 2617 358
rect 2622 352 2625 358
rect 2606 342 2609 348
rect 2622 301 2625 348
rect 2634 338 2638 341
rect 2638 322 2641 328
rect 2622 298 2633 301
rect 2550 272 2553 278
rect 2422 268 2430 271
rect 2362 148 2366 151
rect 2342 112 2345 138
rect 2374 132 2377 158
rect 2406 152 2409 168
rect 2394 148 2398 151
rect 2326 98 2334 101
rect 2270 82 2273 88
rect 2334 82 2337 98
rect 2294 72 2297 78
rect 2282 68 2286 71
rect 1974 52 1977 58
rect 2006 52 2009 58
rect 2070 52 2073 59
rect 2162 58 2166 61
rect 2318 62 2321 68
rect 2390 62 2393 148
rect 2422 142 2425 268
rect 2438 262 2441 268
rect 2430 162 2433 238
rect 2410 138 2414 141
rect 2422 132 2425 138
rect 2414 102 2417 118
rect 2406 82 2409 98
rect 2414 82 2417 88
rect 2438 62 2441 118
rect 2446 72 2449 238
rect 2462 192 2465 258
rect 2486 252 2489 258
rect 2518 252 2521 259
rect 2558 192 2561 218
rect 2574 192 2577 278
rect 2614 262 2617 268
rect 2478 162 2481 188
rect 2466 148 2470 151
rect 2486 142 2489 148
rect 2502 142 2505 188
rect 2510 172 2513 178
rect 2518 152 2521 158
rect 2526 152 2529 158
rect 2590 142 2593 148
rect 2458 138 2462 141
rect 2486 72 2489 128
rect 2494 122 2497 138
rect 2454 62 2457 68
rect 2494 62 2497 78
rect 2502 72 2505 138
rect 2566 132 2569 138
rect 2510 82 2513 118
rect 2526 92 2529 128
rect 2550 122 2553 128
rect 2534 82 2537 98
rect 2550 92 2553 108
rect 2574 102 2577 128
rect 2598 122 2601 148
rect 2614 142 2617 258
rect 2574 82 2577 88
rect 2582 82 2585 98
rect 2618 88 2622 91
rect 2530 78 2534 81
rect 2562 78 2566 81
rect 2594 78 2598 81
rect 2606 72 2609 88
rect 2518 62 2521 68
rect 2558 62 2561 68
rect 2630 62 2633 298
rect 2638 262 2641 268
rect 2638 152 2641 158
rect 2646 92 2649 328
rect 2654 82 2657 318
rect 2662 282 2665 338
rect 2678 332 2681 358
rect 2694 292 2697 478
rect 2702 472 2705 478
rect 2690 118 2694 121
rect 2638 72 2641 78
rect 2290 58 2294 61
rect 2330 58 2334 61
rect 2362 58 2366 61
rect 2426 58 2430 61
rect 2546 58 2550 61
rect 2398 52 2401 58
rect 2606 52 2609 58
rect 2654 52 2657 78
rect 2678 62 2681 118
rect 2694 92 2697 108
rect 2686 82 2689 88
rect 2466 48 2470 51
rect 2618 48 2622 51
rect 1822 -18 1825 18
rect 1718 -19 1722 -18
rect 1710 -22 1722 -19
rect 1822 -22 1826 -18
rect 1838 -22 1842 -18
rect 1934 -22 1938 -18
rect 1990 -19 1994 -18
rect 1998 -19 2001 18
rect 1990 -22 2001 -19
rect 2054 -22 2058 -18
rect 2182 -22 2186 -18
rect 2334 -22 2338 -18
rect 2406 -22 2410 -18
rect 2518 -22 2522 -18
rect 2662 -19 2665 18
rect 2670 -19 2674 -18
rect 2662 -22 2674 -19
<< m3contact >>
rect 14 1758 18 1762
rect 54 1758 58 1762
rect 94 1758 98 1762
rect 102 1758 106 1762
rect 6 1738 10 1742
rect 62 1738 66 1742
rect 86 1738 90 1742
rect 158 1738 162 1742
rect 54 1728 58 1732
rect 62 1668 66 1672
rect 54 1658 58 1662
rect 46 1558 50 1562
rect 30 1548 34 1552
rect 134 1718 138 1722
rect 118 1708 122 1712
rect 142 1708 146 1712
rect 454 1798 458 1802
rect 578 1803 582 1807
rect 585 1803 589 1807
rect 742 1798 746 1802
rect 790 1798 794 1802
rect 838 1798 842 1802
rect 758 1778 762 1782
rect 766 1778 770 1782
rect 782 1778 786 1782
rect 742 1768 746 1772
rect 262 1738 266 1742
rect 302 1738 306 1742
rect 374 1738 378 1742
rect 398 1738 402 1742
rect 446 1738 450 1742
rect 214 1728 218 1732
rect 238 1728 242 1732
rect 246 1728 250 1732
rect 206 1718 210 1722
rect 110 1668 114 1672
rect 382 1728 386 1732
rect 270 1718 274 1722
rect 302 1718 306 1722
rect 198 1668 202 1672
rect 118 1658 122 1662
rect 174 1658 178 1662
rect 190 1658 194 1662
rect 238 1658 242 1662
rect 254 1658 258 1662
rect 134 1648 138 1652
rect 102 1638 106 1642
rect 78 1578 82 1582
rect 78 1548 82 1552
rect 30 1518 34 1522
rect 6 1488 10 1492
rect 38 1468 42 1472
rect 54 1498 58 1502
rect 54 1478 58 1482
rect 134 1588 138 1592
rect 318 1678 322 1682
rect 310 1668 314 1672
rect 294 1658 298 1662
rect 166 1588 170 1592
rect 142 1578 146 1582
rect 142 1568 146 1572
rect 166 1568 170 1572
rect 206 1568 210 1572
rect 134 1548 138 1552
rect 142 1548 146 1552
rect 262 1578 266 1582
rect 214 1548 218 1552
rect 246 1548 250 1552
rect 190 1538 194 1542
rect 86 1488 90 1492
rect 238 1538 242 1542
rect 294 1558 298 1562
rect 326 1658 330 1662
rect 350 1678 354 1682
rect 358 1668 362 1672
rect 382 1648 386 1652
rect 406 1728 410 1732
rect 454 1728 458 1732
rect 430 1678 434 1682
rect 422 1668 426 1672
rect 654 1748 658 1752
rect 502 1738 506 1742
rect 582 1738 586 1742
rect 494 1718 498 1722
rect 470 1678 474 1682
rect 526 1718 530 1722
rect 622 1718 626 1722
rect 510 1678 514 1682
rect 446 1668 450 1672
rect 526 1668 530 1672
rect 550 1668 554 1672
rect 566 1668 570 1672
rect 430 1638 434 1642
rect 350 1578 354 1582
rect 358 1568 362 1572
rect 334 1558 338 1562
rect 350 1558 354 1562
rect 326 1548 330 1552
rect 366 1548 370 1552
rect 390 1558 394 1562
rect 614 1668 618 1672
rect 502 1658 506 1662
rect 534 1658 538 1662
rect 582 1658 586 1662
rect 550 1648 554 1652
rect 622 1648 626 1652
rect 478 1638 482 1642
rect 614 1638 618 1642
rect 646 1638 650 1642
rect 578 1603 582 1607
rect 585 1603 589 1607
rect 470 1578 474 1582
rect 502 1578 506 1582
rect 406 1548 410 1552
rect 278 1538 282 1542
rect 302 1538 306 1542
rect 382 1538 386 1542
rect 254 1528 258 1532
rect 390 1528 394 1532
rect 414 1528 418 1532
rect 430 1528 434 1532
rect 158 1518 162 1522
rect 102 1488 106 1492
rect 102 1468 106 1472
rect 126 1478 130 1482
rect 46 1458 50 1462
rect 78 1458 82 1462
rect 62 1448 66 1452
rect 78 1448 82 1452
rect 94 1448 98 1452
rect 110 1448 114 1452
rect 142 1448 146 1452
rect 14 1378 18 1382
rect 70 1348 74 1352
rect 22 1328 26 1332
rect 70 1328 74 1332
rect 54 1308 58 1312
rect 14 1288 18 1292
rect 166 1488 170 1492
rect 246 1498 250 1502
rect 182 1478 186 1482
rect 238 1478 242 1482
rect 214 1468 218 1472
rect 230 1468 234 1472
rect 174 1448 178 1452
rect 494 1568 498 1572
rect 566 1558 570 1562
rect 510 1548 514 1552
rect 606 1518 610 1522
rect 438 1498 442 1502
rect 534 1498 538 1502
rect 294 1488 298 1492
rect 438 1488 442 1492
rect 518 1488 522 1492
rect 278 1478 282 1482
rect 502 1478 506 1482
rect 438 1468 442 1472
rect 166 1368 170 1372
rect 150 1358 154 1362
rect 158 1358 162 1362
rect 174 1358 178 1362
rect 102 1348 106 1352
rect 118 1348 122 1352
rect 150 1348 154 1352
rect 166 1348 170 1352
rect 134 1338 138 1342
rect 206 1348 210 1352
rect 102 1328 106 1332
rect 46 1288 50 1292
rect 70 1288 74 1292
rect 62 1268 66 1272
rect 70 1258 74 1262
rect 86 1258 90 1262
rect 54 1248 58 1252
rect 6 1168 10 1172
rect 62 1138 66 1142
rect 46 1098 50 1102
rect 30 1078 34 1082
rect 38 1078 42 1082
rect 54 1078 58 1082
rect 14 1068 18 1072
rect 46 1068 50 1072
rect 118 1308 122 1312
rect 198 1308 202 1312
rect 126 1268 130 1272
rect 182 1268 186 1272
rect 166 1258 170 1262
rect 182 1258 186 1262
rect 182 1228 186 1232
rect 166 1168 170 1172
rect 110 1138 114 1142
rect 118 1128 122 1132
rect 134 1118 138 1122
rect 110 1088 114 1092
rect 222 1298 226 1302
rect 214 1248 218 1252
rect 262 1388 266 1392
rect 286 1378 290 1382
rect 254 1368 258 1372
rect 270 1368 274 1372
rect 238 1348 242 1352
rect 270 1348 274 1352
rect 310 1378 314 1382
rect 294 1358 298 1362
rect 294 1348 298 1352
rect 318 1328 322 1332
rect 262 1308 266 1312
rect 246 1298 250 1302
rect 238 1288 242 1292
rect 358 1438 362 1442
rect 406 1438 410 1442
rect 390 1408 394 1412
rect 342 1388 346 1392
rect 334 1358 338 1362
rect 262 1278 266 1282
rect 286 1278 290 1282
rect 302 1278 306 1282
rect 326 1278 330 1282
rect 246 1268 250 1272
rect 302 1268 306 1272
rect 310 1268 314 1272
rect 270 1248 274 1252
rect 238 1238 242 1242
rect 206 1148 210 1152
rect 174 1128 178 1132
rect 238 1148 242 1152
rect 270 1138 274 1142
rect 214 1128 218 1132
rect 262 1128 266 1132
rect 302 1178 306 1182
rect 294 1158 298 1162
rect 318 1228 322 1232
rect 366 1348 370 1352
rect 510 1458 514 1462
rect 646 1558 650 1562
rect 630 1548 634 1552
rect 678 1678 682 1682
rect 726 1678 730 1682
rect 630 1478 634 1482
rect 718 1658 722 1662
rect 726 1648 730 1652
rect 686 1638 690 1642
rect 710 1618 714 1622
rect 734 1638 738 1642
rect 750 1618 754 1622
rect 894 1758 898 1762
rect 934 1758 938 1762
rect 838 1748 842 1752
rect 910 1748 914 1752
rect 918 1748 922 1752
rect 918 1738 922 1742
rect 886 1678 890 1682
rect 806 1658 810 1662
rect 822 1658 826 1662
rect 846 1638 850 1642
rect 894 1668 898 1672
rect 910 1648 914 1652
rect 886 1618 890 1622
rect 742 1538 746 1542
rect 782 1538 786 1542
rect 750 1528 754 1532
rect 774 1528 778 1532
rect 702 1518 706 1522
rect 678 1488 682 1492
rect 726 1488 730 1492
rect 670 1478 674 1482
rect 574 1468 578 1472
rect 630 1468 634 1472
rect 558 1458 562 1462
rect 542 1448 546 1452
rect 462 1438 466 1442
rect 550 1438 554 1442
rect 622 1438 626 1442
rect 578 1403 582 1407
rect 585 1403 589 1407
rect 422 1358 426 1362
rect 342 1278 346 1282
rect 350 1278 354 1282
rect 390 1328 394 1332
rect 390 1308 394 1312
rect 382 1288 386 1292
rect 422 1288 426 1292
rect 358 1268 362 1272
rect 374 1268 378 1272
rect 422 1268 426 1272
rect 342 1258 346 1262
rect 390 1248 394 1252
rect 414 1238 418 1242
rect 350 1228 354 1232
rect 502 1368 506 1372
rect 558 1358 562 1362
rect 518 1348 522 1352
rect 574 1348 578 1352
rect 438 1278 442 1282
rect 486 1328 490 1332
rect 510 1328 514 1332
rect 526 1328 530 1332
rect 494 1288 498 1292
rect 470 1248 474 1252
rect 486 1238 490 1242
rect 430 1218 434 1222
rect 462 1218 466 1222
rect 350 1168 354 1172
rect 422 1168 426 1172
rect 334 1158 338 1162
rect 310 1148 314 1152
rect 286 1138 290 1142
rect 278 1118 282 1122
rect 182 1088 186 1092
rect 38 1058 42 1062
rect 62 1058 66 1062
rect 14 958 18 962
rect 6 938 10 942
rect 6 868 10 872
rect 38 1048 42 1052
rect 62 1048 66 1052
rect 86 1068 90 1072
rect 110 1068 114 1072
rect 94 1058 98 1062
rect 158 1058 162 1062
rect 214 1058 218 1062
rect 222 1058 226 1062
rect 198 1048 202 1052
rect 222 1048 226 1052
rect 78 1038 82 1042
rect 126 1038 130 1042
rect 134 1038 138 1042
rect 110 958 114 962
rect 118 948 122 952
rect 142 948 146 952
rect 246 1038 250 1042
rect 238 1028 242 1032
rect 302 1088 306 1092
rect 302 1068 306 1072
rect 390 1158 394 1162
rect 342 1138 346 1142
rect 358 1138 362 1142
rect 470 1138 474 1142
rect 366 1108 370 1112
rect 422 1088 426 1092
rect 582 1318 586 1322
rect 526 1278 530 1282
rect 534 1278 538 1282
rect 542 1258 546 1262
rect 558 1258 562 1262
rect 574 1258 578 1262
rect 622 1288 626 1292
rect 694 1458 698 1462
rect 774 1468 778 1472
rect 726 1448 730 1452
rect 742 1438 746 1442
rect 750 1398 754 1402
rect 662 1348 666 1352
rect 678 1348 682 1352
rect 630 1278 634 1282
rect 646 1268 650 1272
rect 662 1268 666 1272
rect 726 1288 730 1292
rect 694 1238 698 1242
rect 654 1228 658 1232
rect 606 1218 610 1222
rect 578 1203 582 1207
rect 585 1203 589 1207
rect 750 1278 754 1282
rect 822 1478 826 1482
rect 870 1548 874 1552
rect 894 1548 898 1552
rect 862 1538 866 1542
rect 910 1538 914 1542
rect 854 1488 858 1492
rect 870 1478 874 1482
rect 838 1458 842 1462
rect 870 1458 874 1462
rect 886 1458 890 1462
rect 838 1448 842 1452
rect 854 1448 858 1452
rect 1062 1748 1066 1752
rect 1070 1748 1074 1752
rect 1142 1748 1146 1752
rect 1014 1738 1018 1742
rect 990 1728 994 1732
rect 1198 1738 1202 1742
rect 1206 1738 1210 1742
rect 1078 1718 1082 1722
rect 1118 1718 1122 1722
rect 1118 1708 1122 1712
rect 1166 1708 1170 1712
rect 1082 1703 1086 1707
rect 1089 1703 1093 1707
rect 1062 1688 1066 1692
rect 1150 1688 1154 1692
rect 1206 1718 1210 1722
rect 1214 1698 1218 1702
rect 1078 1678 1082 1682
rect 1206 1678 1210 1682
rect 1294 1748 1298 1752
rect 1542 1748 1546 1752
rect 1254 1688 1258 1692
rect 974 1668 978 1672
rect 1014 1668 1018 1672
rect 1038 1668 1042 1672
rect 982 1658 986 1662
rect 998 1648 1002 1652
rect 990 1628 994 1632
rect 998 1558 1002 1562
rect 926 1548 930 1552
rect 942 1548 946 1552
rect 1102 1659 1106 1663
rect 1022 1638 1026 1642
rect 1190 1638 1194 1642
rect 1206 1618 1210 1622
rect 1270 1738 1274 1742
rect 1294 1718 1298 1722
rect 1334 1718 1338 1722
rect 1398 1718 1402 1722
rect 1406 1718 1410 1722
rect 1310 1688 1314 1692
rect 1334 1678 1338 1682
rect 1342 1678 1346 1682
rect 1278 1668 1282 1672
rect 1262 1628 1266 1632
rect 1014 1568 1018 1572
rect 1038 1558 1042 1562
rect 1174 1558 1178 1562
rect 1326 1658 1330 1662
rect 1326 1618 1330 1622
rect 1414 1658 1418 1662
rect 1366 1638 1370 1642
rect 1382 1638 1386 1642
rect 1342 1628 1346 1632
rect 1358 1558 1362 1562
rect 1070 1548 1074 1552
rect 1094 1548 1098 1552
rect 1334 1548 1338 1552
rect 1358 1548 1362 1552
rect 1366 1548 1370 1552
rect 950 1528 954 1532
rect 998 1528 1002 1532
rect 1006 1528 1010 1532
rect 1030 1528 1034 1532
rect 1046 1528 1050 1532
rect 1078 1528 1082 1532
rect 934 1488 938 1492
rect 942 1488 946 1492
rect 982 1518 986 1522
rect 950 1468 954 1472
rect 958 1458 962 1462
rect 886 1438 890 1442
rect 902 1438 906 1442
rect 870 1418 874 1422
rect 862 1388 866 1392
rect 838 1378 842 1382
rect 878 1378 882 1382
rect 790 1338 794 1342
rect 846 1338 850 1342
rect 790 1278 794 1282
rect 750 1268 754 1272
rect 766 1258 770 1262
rect 742 1188 746 1192
rect 502 1168 506 1172
rect 558 1168 562 1172
rect 702 1168 706 1172
rect 734 1168 738 1172
rect 750 1168 754 1172
rect 542 1148 546 1152
rect 598 1148 602 1152
rect 630 1138 634 1142
rect 638 1128 642 1132
rect 598 1118 602 1122
rect 630 1118 634 1122
rect 638 1108 642 1112
rect 638 1098 642 1102
rect 662 1098 666 1102
rect 526 1088 530 1092
rect 558 1088 562 1092
rect 598 1088 602 1092
rect 374 1078 378 1082
rect 454 1078 458 1082
rect 486 1078 490 1082
rect 518 1078 522 1082
rect 422 1068 426 1072
rect 454 1068 458 1072
rect 350 1058 354 1062
rect 414 1058 418 1062
rect 334 1038 338 1042
rect 358 1038 362 1042
rect 318 1028 322 1032
rect 230 958 234 962
rect 286 958 290 962
rect 246 948 250 952
rect 654 1088 658 1092
rect 550 1068 554 1072
rect 582 1068 586 1072
rect 478 1058 482 1062
rect 366 968 370 972
rect 430 958 434 962
rect 470 958 474 962
rect 406 948 410 952
rect 94 938 98 942
rect 246 938 250 942
rect 262 938 266 942
rect 358 938 362 942
rect 366 938 370 942
rect 470 938 474 942
rect 78 928 82 932
rect 62 918 66 922
rect 30 868 34 872
rect 14 848 18 852
rect 86 918 90 922
rect 46 848 50 852
rect 134 928 138 932
rect 134 888 138 892
rect 30 818 34 822
rect 62 818 66 822
rect 78 778 82 782
rect 54 768 58 772
rect 6 758 10 762
rect 230 928 234 932
rect 190 888 194 892
rect 270 888 274 892
rect 214 878 218 882
rect 510 1048 514 1052
rect 534 1048 538 1052
rect 486 948 490 952
rect 510 948 514 952
rect 438 928 442 932
rect 478 928 482 932
rect 678 1078 682 1082
rect 550 1038 554 1042
rect 614 1038 618 1042
rect 686 1038 690 1042
rect 582 1018 586 1022
rect 578 1003 582 1007
rect 585 1003 589 1007
rect 638 988 642 992
rect 662 978 666 982
rect 614 958 618 962
rect 502 938 506 942
rect 526 938 530 942
rect 534 938 538 942
rect 350 918 354 922
rect 382 918 386 922
rect 422 918 426 922
rect 446 918 450 922
rect 462 918 466 922
rect 302 898 306 902
rect 654 947 658 951
rect 550 928 554 932
rect 598 928 602 932
rect 542 918 546 922
rect 478 888 482 892
rect 534 888 538 892
rect 518 878 522 882
rect 326 868 330 872
rect 446 868 450 872
rect 494 868 498 872
rect 182 858 186 862
rect 262 858 266 862
rect 158 848 162 852
rect 270 848 274 852
rect 358 848 362 852
rect 110 818 114 822
rect 102 778 106 782
rect 94 758 98 762
rect 174 778 178 782
rect 174 768 178 772
rect 270 768 274 772
rect 302 768 306 772
rect 310 768 314 772
rect 134 758 138 762
rect 166 758 170 762
rect 206 758 210 762
rect 230 758 234 762
rect 254 758 258 762
rect 46 748 50 752
rect 62 748 66 752
rect 102 748 106 752
rect 110 748 114 752
rect 158 748 162 752
rect 182 748 186 752
rect 278 748 282 752
rect 22 738 26 742
rect 502 838 506 842
rect 478 828 482 832
rect 462 788 466 792
rect 446 768 450 772
rect 174 738 178 742
rect 270 738 274 742
rect 422 738 426 742
rect 142 728 146 732
rect 222 728 226 732
rect 246 728 250 732
rect 142 718 146 722
rect 222 718 226 722
rect 238 718 242 722
rect 174 708 178 712
rect 230 708 234 712
rect 182 688 186 692
rect 246 688 250 692
rect 6 668 10 672
rect 70 668 74 672
rect 94 668 98 672
rect 150 668 154 672
rect 182 668 186 672
rect 38 658 42 662
rect 46 658 50 662
rect 22 648 26 652
rect 38 568 42 572
rect 6 528 10 532
rect 62 528 66 532
rect 30 488 34 492
rect 86 658 90 662
rect 78 648 82 652
rect 94 648 98 652
rect 118 638 122 642
rect 86 628 90 632
rect 110 558 114 562
rect 158 648 162 652
rect 198 658 202 662
rect 198 648 202 652
rect 190 638 194 642
rect 134 558 138 562
rect 110 548 114 552
rect 70 468 74 472
rect 30 368 34 372
rect 6 348 10 352
rect 70 458 74 462
rect 86 488 90 492
rect 150 518 154 522
rect 166 548 170 552
rect 174 548 178 552
rect 182 528 186 532
rect 142 478 146 482
rect 206 518 210 522
rect 278 728 282 732
rect 318 718 322 722
rect 334 718 338 722
rect 382 718 386 722
rect 374 708 378 712
rect 310 698 314 702
rect 270 688 274 692
rect 294 688 298 692
rect 454 748 458 752
rect 470 748 474 752
rect 446 738 450 742
rect 462 728 466 732
rect 430 708 434 712
rect 430 688 434 692
rect 286 678 290 682
rect 366 678 370 682
rect 390 678 394 682
rect 414 678 418 682
rect 310 668 314 672
rect 222 658 226 662
rect 254 658 258 662
rect 286 658 290 662
rect 262 648 266 652
rect 294 578 298 582
rect 222 548 226 552
rect 302 568 306 572
rect 318 638 322 642
rect 342 668 346 672
rect 422 668 426 672
rect 358 658 362 662
rect 382 658 386 662
rect 358 648 362 652
rect 422 648 426 652
rect 454 678 458 682
rect 446 648 450 652
rect 454 648 458 652
rect 398 638 402 642
rect 438 638 442 642
rect 334 588 338 592
rect 438 588 442 592
rect 326 548 330 552
rect 382 548 386 552
rect 398 548 402 552
rect 254 518 258 522
rect 246 498 250 502
rect 102 458 106 462
rect 174 458 178 462
rect 94 448 98 452
rect 150 448 154 452
rect 374 538 378 542
rect 350 528 354 532
rect 318 518 322 522
rect 294 478 298 482
rect 302 478 306 482
rect 382 528 386 532
rect 390 528 394 532
rect 406 498 410 502
rect 422 498 426 502
rect 438 488 442 492
rect 366 478 370 482
rect 374 478 378 482
rect 278 468 282 472
rect 198 458 202 462
rect 238 458 242 462
rect 246 458 250 462
rect 286 458 290 462
rect 318 458 322 462
rect 134 358 138 362
rect 126 348 130 352
rect 150 348 154 352
rect 62 338 66 342
rect 142 338 146 342
rect 166 338 170 342
rect 86 298 90 302
rect 6 278 10 282
rect 278 368 282 372
rect 198 358 202 362
rect 270 358 274 362
rect 182 348 186 352
rect 270 348 274 352
rect 198 338 202 342
rect 182 328 186 332
rect 142 318 146 322
rect 134 308 138 312
rect 174 308 178 312
rect 150 288 154 292
rect 38 268 42 272
rect 70 268 74 272
rect 94 268 98 272
rect 62 258 66 262
rect 110 258 114 262
rect 118 258 122 262
rect 238 338 242 342
rect 246 338 250 342
rect 318 438 322 442
rect 302 358 306 362
rect 374 358 378 362
rect 510 758 514 762
rect 526 788 530 792
rect 494 738 498 742
rect 478 728 482 732
rect 494 718 498 722
rect 478 688 482 692
rect 478 668 482 672
rect 518 718 522 722
rect 574 898 578 902
rect 574 888 578 892
rect 558 868 562 872
rect 542 848 546 852
rect 574 868 578 872
rect 758 1148 762 1152
rect 774 1098 778 1102
rect 798 1258 802 1262
rect 814 1248 818 1252
rect 822 1218 826 1222
rect 814 1118 818 1122
rect 782 1078 786 1082
rect 926 1348 930 1352
rect 950 1328 954 1332
rect 838 1258 842 1262
rect 830 1158 834 1162
rect 830 1108 834 1112
rect 934 1268 938 1272
rect 998 1488 1002 1492
rect 998 1468 1002 1472
rect 974 1448 978 1452
rect 1062 1518 1066 1522
rect 1086 1518 1090 1522
rect 1046 1478 1050 1482
rect 1046 1458 1050 1462
rect 1082 1503 1086 1507
rect 1089 1503 1093 1507
rect 1094 1478 1098 1482
rect 1102 1468 1106 1472
rect 1070 1458 1074 1462
rect 1038 1448 1042 1452
rect 1078 1378 1082 1382
rect 1006 1358 1010 1362
rect 1030 1358 1034 1362
rect 990 1338 994 1342
rect 982 1328 986 1332
rect 1038 1328 1042 1332
rect 1006 1318 1010 1322
rect 1038 1318 1042 1322
rect 998 1278 1002 1282
rect 990 1266 994 1270
rect 1006 1268 1010 1272
rect 1054 1308 1058 1312
rect 1118 1528 1122 1532
rect 1198 1528 1202 1532
rect 1118 1498 1122 1502
rect 1150 1498 1154 1502
rect 1118 1488 1122 1492
rect 1126 1478 1130 1482
rect 1206 1478 1210 1482
rect 1222 1478 1226 1482
rect 1190 1468 1194 1472
rect 1198 1468 1202 1472
rect 1110 1368 1114 1372
rect 1150 1458 1154 1462
rect 1174 1458 1178 1462
rect 1126 1448 1130 1452
rect 1166 1438 1170 1442
rect 1126 1358 1130 1362
rect 1118 1348 1122 1352
rect 1070 1328 1074 1332
rect 1082 1303 1086 1307
rect 1089 1303 1093 1307
rect 1118 1328 1122 1332
rect 1182 1428 1186 1432
rect 1350 1538 1354 1542
rect 1294 1528 1298 1532
rect 1270 1508 1274 1512
rect 1334 1518 1338 1522
rect 1398 1628 1402 1632
rect 1470 1718 1474 1722
rect 1478 1658 1482 1662
rect 1422 1618 1426 1622
rect 1406 1558 1410 1562
rect 1374 1538 1378 1542
rect 1366 1518 1370 1522
rect 1446 1547 1450 1551
rect 1422 1538 1426 1542
rect 1398 1508 1402 1512
rect 1350 1468 1354 1472
rect 1382 1468 1386 1472
rect 1278 1448 1282 1452
rect 1286 1428 1290 1432
rect 1470 1528 1474 1532
rect 1602 1803 1606 1807
rect 1609 1803 1613 1807
rect 1734 1798 1738 1802
rect 1782 1798 1786 1802
rect 2022 1778 2026 1782
rect 2158 1778 2162 1782
rect 2502 1778 2506 1782
rect 1838 1768 1842 1772
rect 1870 1768 1874 1772
rect 2054 1768 2058 1772
rect 2222 1768 2226 1772
rect 2086 1758 2090 1762
rect 2382 1758 2386 1762
rect 1654 1748 1658 1752
rect 1662 1748 1666 1752
rect 1838 1748 1842 1752
rect 1606 1738 1610 1742
rect 1670 1738 1674 1742
rect 1646 1728 1650 1732
rect 1534 1688 1538 1692
rect 1542 1688 1546 1692
rect 1534 1668 1538 1672
rect 1518 1658 1522 1662
rect 1510 1568 1514 1572
rect 1502 1558 1506 1562
rect 1582 1668 1586 1672
rect 1598 1658 1602 1662
rect 1582 1648 1586 1652
rect 1550 1558 1554 1562
rect 1602 1603 1606 1607
rect 1609 1603 1613 1607
rect 1598 1568 1602 1572
rect 1718 1738 1722 1742
rect 1750 1728 1754 1732
rect 1774 1728 1778 1732
rect 1718 1688 1722 1692
rect 1806 1688 1810 1692
rect 1734 1678 1738 1682
rect 1750 1668 1754 1672
rect 1702 1658 1706 1662
rect 1678 1648 1682 1652
rect 1822 1648 1826 1652
rect 1718 1568 1722 1572
rect 1654 1558 1658 1562
rect 1726 1558 1730 1562
rect 1798 1558 1802 1562
rect 1822 1558 1826 1562
rect 1686 1548 1690 1552
rect 1734 1548 1738 1552
rect 1526 1538 1530 1542
rect 1582 1538 1586 1542
rect 1710 1538 1714 1542
rect 1518 1528 1522 1532
rect 1438 1468 1442 1472
rect 1534 1468 1538 1472
rect 1694 1528 1698 1532
rect 1766 1538 1770 1542
rect 1782 1538 1786 1542
rect 1734 1518 1738 1522
rect 1766 1518 1770 1522
rect 1798 1518 1802 1522
rect 1750 1508 1754 1512
rect 1710 1478 1714 1482
rect 1726 1478 1730 1482
rect 1406 1458 1410 1462
rect 1430 1458 1434 1462
rect 1446 1458 1450 1462
rect 1526 1458 1530 1462
rect 1662 1458 1666 1462
rect 1734 1458 1738 1462
rect 1230 1388 1234 1392
rect 1318 1388 1322 1392
rect 1182 1378 1186 1382
rect 1206 1368 1210 1372
rect 1182 1328 1186 1332
rect 1198 1328 1202 1332
rect 1142 1318 1146 1322
rect 1182 1318 1186 1322
rect 1062 1288 1066 1292
rect 1118 1288 1122 1292
rect 1134 1288 1138 1292
rect 1054 1278 1058 1282
rect 1142 1278 1146 1282
rect 1158 1278 1162 1282
rect 974 1248 978 1252
rect 1014 1248 1018 1252
rect 966 1228 970 1232
rect 846 1218 850 1222
rect 918 1218 922 1222
rect 1054 1208 1058 1212
rect 1014 1178 1018 1182
rect 1134 1268 1138 1272
rect 1110 1258 1114 1262
rect 1238 1348 1242 1352
rect 1246 1288 1250 1292
rect 1206 1278 1210 1282
rect 1238 1278 1242 1282
rect 1198 1268 1202 1272
rect 1278 1318 1282 1322
rect 1286 1288 1290 1292
rect 1302 1278 1306 1282
rect 1270 1268 1274 1272
rect 1190 1258 1194 1262
rect 1254 1258 1258 1262
rect 1142 1248 1146 1252
rect 1174 1248 1178 1252
rect 1158 1238 1162 1242
rect 1134 1228 1138 1232
rect 1166 1228 1170 1232
rect 1214 1198 1218 1202
rect 1262 1238 1266 1242
rect 1062 1168 1066 1172
rect 854 1158 858 1162
rect 902 1158 906 1162
rect 1062 1158 1066 1162
rect 1086 1158 1090 1162
rect 886 1148 890 1152
rect 926 1147 930 1151
rect 998 1148 1002 1152
rect 1126 1148 1130 1152
rect 1174 1148 1178 1152
rect 934 1138 938 1142
rect 870 1128 874 1132
rect 878 1128 882 1132
rect 902 1118 906 1122
rect 846 1108 850 1112
rect 902 1108 906 1112
rect 870 1098 874 1102
rect 870 1088 874 1092
rect 838 1078 842 1082
rect 830 1068 834 1072
rect 774 1058 778 1062
rect 742 1048 746 1052
rect 806 1048 810 1052
rect 822 1048 826 1052
rect 1022 1138 1026 1142
rect 1054 1138 1058 1142
rect 1078 1138 1082 1142
rect 1166 1138 1170 1142
rect 982 1128 986 1132
rect 1102 1128 1106 1132
rect 1134 1128 1138 1132
rect 990 1118 994 1122
rect 998 1118 1002 1122
rect 1006 1108 1010 1112
rect 1014 1098 1018 1102
rect 950 1078 954 1082
rect 1006 1078 1010 1082
rect 886 1068 890 1072
rect 894 1048 898 1052
rect 910 1048 914 1052
rect 846 1038 850 1042
rect 862 1038 866 1042
rect 838 1008 842 1012
rect 750 988 754 992
rect 742 968 746 972
rect 726 958 730 962
rect 726 948 730 952
rect 678 878 682 882
rect 710 878 714 882
rect 598 858 602 862
rect 582 848 586 852
rect 566 828 570 832
rect 630 848 634 852
rect 774 978 778 982
rect 814 968 818 972
rect 846 968 850 972
rect 870 958 874 962
rect 790 938 794 942
rect 814 928 818 932
rect 766 898 770 902
rect 758 888 762 892
rect 750 878 754 882
rect 734 868 738 872
rect 766 858 770 862
rect 750 848 754 852
rect 654 838 658 842
rect 726 838 730 842
rect 622 818 626 822
rect 578 803 582 807
rect 585 803 589 807
rect 574 788 578 792
rect 558 768 562 772
rect 606 768 610 772
rect 542 738 546 742
rect 558 708 562 712
rect 550 678 554 682
rect 534 668 538 672
rect 742 818 746 822
rect 726 768 730 772
rect 654 758 658 762
rect 718 758 722 762
rect 654 747 658 751
rect 694 748 698 752
rect 726 748 730 752
rect 622 708 626 712
rect 566 698 570 702
rect 598 668 602 672
rect 614 668 618 672
rect 510 658 514 662
rect 606 658 610 662
rect 598 638 602 642
rect 486 618 490 622
rect 578 603 582 607
rect 585 603 589 607
rect 542 588 546 592
rect 526 568 530 572
rect 494 558 498 562
rect 510 548 514 552
rect 534 538 538 542
rect 470 488 474 492
rect 494 468 498 472
rect 526 468 530 472
rect 494 358 498 362
rect 542 488 546 492
rect 574 508 578 512
rect 574 488 578 492
rect 646 648 650 652
rect 718 738 722 742
rect 694 728 698 732
rect 678 708 682 712
rect 702 718 706 722
rect 662 668 666 672
rect 694 668 698 672
rect 686 658 690 662
rect 638 638 642 642
rect 630 608 634 612
rect 654 588 658 592
rect 662 568 666 572
rect 694 568 698 572
rect 846 928 850 932
rect 958 1068 962 1072
rect 974 1068 978 1072
rect 990 1068 994 1072
rect 1082 1103 1086 1107
rect 1089 1103 1093 1107
rect 1070 1098 1074 1102
rect 1110 1088 1114 1092
rect 1030 1078 1034 1082
rect 1054 1078 1058 1082
rect 1038 1068 1042 1072
rect 1070 1068 1074 1072
rect 1078 1068 1082 1072
rect 1150 1118 1154 1122
rect 1134 1058 1138 1062
rect 1158 1058 1162 1062
rect 958 1048 962 1052
rect 974 1048 978 1052
rect 1118 1048 1122 1052
rect 1078 1038 1082 1042
rect 1246 1128 1250 1132
rect 1262 1138 1266 1142
rect 1206 1088 1210 1092
rect 1254 1088 1258 1092
rect 1286 1248 1290 1252
rect 1286 1228 1290 1232
rect 1358 1398 1362 1402
rect 1438 1398 1442 1402
rect 1374 1388 1378 1392
rect 1598 1448 1602 1452
rect 1598 1418 1602 1422
rect 1638 1418 1642 1422
rect 1602 1403 1606 1407
rect 1609 1403 1613 1407
rect 1350 1348 1354 1352
rect 1422 1348 1426 1352
rect 1342 1318 1346 1322
rect 1582 1348 1586 1352
rect 1614 1338 1618 1342
rect 1566 1318 1570 1322
rect 1590 1318 1594 1322
rect 1758 1418 1762 1422
rect 1782 1508 1786 1512
rect 1822 1518 1826 1522
rect 1814 1498 1818 1502
rect 1806 1488 1810 1492
rect 1806 1478 1810 1482
rect 1790 1468 1794 1472
rect 1822 1488 1826 1492
rect 1774 1438 1778 1442
rect 1766 1398 1770 1402
rect 1854 1738 1858 1742
rect 1838 1728 1842 1732
rect 1910 1718 1914 1722
rect 2198 1748 2202 1752
rect 2230 1748 2234 1752
rect 2246 1748 2250 1752
rect 2278 1748 2282 1752
rect 1990 1738 1994 1742
rect 2006 1738 2010 1742
rect 2174 1738 2178 1742
rect 2190 1738 2194 1742
rect 2054 1728 2058 1732
rect 2038 1718 2042 1722
rect 1934 1698 1938 1702
rect 1838 1658 1842 1662
rect 1910 1658 1914 1662
rect 2030 1708 2034 1712
rect 1846 1648 1850 1652
rect 1982 1648 1986 1652
rect 1990 1648 1994 1652
rect 2070 1708 2074 1712
rect 2062 1698 2066 1702
rect 2106 1703 2110 1707
rect 2113 1703 2117 1707
rect 2142 1698 2146 1702
rect 2086 1688 2090 1692
rect 2070 1678 2074 1682
rect 1878 1638 1882 1642
rect 2038 1638 2042 1642
rect 1934 1608 1938 1612
rect 1910 1568 1914 1572
rect 1838 1558 1842 1562
rect 1958 1578 1962 1582
rect 1998 1568 2002 1572
rect 1918 1548 1922 1552
rect 1934 1548 1938 1552
rect 1990 1548 1994 1552
rect 1846 1528 1850 1532
rect 1838 1488 1842 1492
rect 1814 1458 1818 1462
rect 1830 1458 1834 1462
rect 1790 1448 1794 1452
rect 1758 1388 1762 1392
rect 1782 1368 1786 1372
rect 1694 1358 1698 1362
rect 1766 1358 1770 1362
rect 1678 1338 1682 1342
rect 1662 1328 1666 1332
rect 1614 1288 1618 1292
rect 1478 1278 1482 1282
rect 1502 1278 1506 1282
rect 1526 1278 1530 1282
rect 1534 1278 1538 1282
rect 1582 1278 1586 1282
rect 1590 1278 1594 1282
rect 1334 1268 1338 1272
rect 1406 1268 1410 1272
rect 1470 1268 1474 1272
rect 1382 1258 1386 1262
rect 1390 1248 1394 1252
rect 1326 1198 1330 1202
rect 1286 1168 1290 1172
rect 1302 1168 1306 1172
rect 1310 1168 1314 1172
rect 1342 1168 1346 1172
rect 1422 1238 1426 1242
rect 1454 1258 1458 1262
rect 1470 1258 1474 1262
rect 1526 1258 1530 1262
rect 1510 1248 1514 1252
rect 1398 1228 1402 1232
rect 1446 1228 1450 1232
rect 1486 1228 1490 1232
rect 1414 1198 1418 1202
rect 1446 1198 1450 1202
rect 1358 1158 1362 1162
rect 1302 1138 1306 1142
rect 1318 1138 1322 1142
rect 1350 1148 1354 1152
rect 1526 1178 1530 1182
rect 1518 1168 1522 1172
rect 1494 1158 1498 1162
rect 1502 1148 1506 1152
rect 1582 1248 1586 1252
rect 1566 1238 1570 1242
rect 1602 1203 1606 1207
rect 1609 1203 1613 1207
rect 1590 1188 1594 1192
rect 1598 1188 1602 1192
rect 1550 1178 1554 1182
rect 1534 1158 1538 1162
rect 1342 1138 1346 1142
rect 1358 1138 1362 1142
rect 1406 1138 1410 1142
rect 1446 1138 1450 1142
rect 1494 1138 1498 1142
rect 1326 1128 1330 1132
rect 1366 1128 1370 1132
rect 1398 1128 1402 1132
rect 1414 1128 1418 1132
rect 1470 1128 1474 1132
rect 1342 1088 1346 1092
rect 1302 1078 1306 1082
rect 1374 1078 1378 1082
rect 1182 1068 1186 1072
rect 1190 1068 1194 1072
rect 1238 1068 1242 1072
rect 1246 1068 1250 1072
rect 1222 1058 1226 1062
rect 1198 1048 1202 1052
rect 1166 1038 1170 1042
rect 1150 1028 1154 1032
rect 942 1018 946 1022
rect 1086 1018 1090 1022
rect 1182 1018 1186 1022
rect 886 938 890 942
rect 934 938 938 942
rect 918 908 922 912
rect 862 898 866 902
rect 878 898 882 902
rect 886 898 890 902
rect 814 888 818 892
rect 822 888 826 892
rect 934 888 938 892
rect 846 878 850 882
rect 1022 1008 1026 1012
rect 982 998 986 1002
rect 982 978 986 982
rect 1006 978 1010 982
rect 950 958 954 962
rect 974 958 978 962
rect 1014 948 1018 952
rect 998 938 1002 942
rect 758 768 762 772
rect 798 768 802 772
rect 742 728 746 732
rect 734 708 738 712
rect 718 698 722 702
rect 766 748 770 752
rect 782 748 786 752
rect 966 928 970 932
rect 982 928 986 932
rect 1006 898 1010 902
rect 966 878 970 882
rect 990 868 994 872
rect 950 768 954 772
rect 894 748 898 752
rect 838 728 842 732
rect 758 718 762 722
rect 790 708 794 712
rect 838 708 842 712
rect 950 748 954 752
rect 974 748 978 752
rect 902 738 906 742
rect 918 738 922 742
rect 750 688 754 692
rect 758 688 762 692
rect 718 638 722 642
rect 718 628 722 632
rect 750 628 754 632
rect 718 608 722 612
rect 630 547 634 551
rect 678 548 682 552
rect 686 548 690 552
rect 622 538 626 542
rect 670 538 674 542
rect 614 518 618 522
rect 694 518 698 522
rect 662 498 666 502
rect 558 478 562 482
rect 694 478 698 482
rect 702 478 706 482
rect 630 468 634 472
rect 654 468 658 472
rect 630 458 634 462
rect 646 458 650 462
rect 694 458 698 462
rect 558 418 562 422
rect 578 403 582 407
rect 585 403 589 407
rect 694 448 698 452
rect 638 428 642 432
rect 670 428 674 432
rect 566 388 570 392
rect 558 358 562 362
rect 454 348 458 352
rect 470 348 474 352
rect 502 348 506 352
rect 622 358 626 362
rect 662 358 666 362
rect 310 338 314 342
rect 414 338 418 342
rect 446 338 450 342
rect 214 318 218 322
rect 238 318 242 322
rect 286 308 290 312
rect 206 288 210 292
rect 222 288 226 292
rect 182 278 186 282
rect 214 278 218 282
rect 406 308 410 312
rect 166 268 170 272
rect 254 268 258 272
rect 294 268 298 272
rect 366 268 370 272
rect 438 268 442 272
rect 278 258 282 262
rect 310 258 314 262
rect 438 258 442 262
rect 174 248 178 252
rect 198 248 202 252
rect 246 248 250 252
rect 294 248 298 252
rect 358 228 362 232
rect 390 228 394 232
rect 470 258 474 262
rect 454 248 458 252
rect 462 218 466 222
rect 398 158 402 162
rect 30 148 34 152
rect 94 148 98 152
rect 158 148 162 152
rect 230 148 234 152
rect 262 148 266 152
rect 310 148 314 152
rect 342 148 346 152
rect 438 148 442 152
rect 14 118 18 122
rect 22 118 26 122
rect 6 78 10 82
rect 46 128 50 132
rect 54 88 58 92
rect 86 88 90 92
rect 126 88 130 92
rect 158 88 162 92
rect 38 58 42 62
rect 94 58 98 62
rect 142 58 146 62
rect 486 228 490 232
rect 470 148 474 152
rect 638 348 642 352
rect 662 278 666 282
rect 734 548 738 552
rect 718 508 722 512
rect 798 668 802 672
rect 782 628 786 632
rect 894 698 898 702
rect 846 688 850 692
rect 854 668 858 672
rect 822 658 826 662
rect 950 738 954 742
rect 942 718 946 722
rect 934 678 938 682
rect 886 658 890 662
rect 902 658 906 662
rect 894 648 898 652
rect 926 648 930 652
rect 822 638 826 642
rect 886 638 890 642
rect 910 638 914 642
rect 846 628 850 632
rect 806 588 810 592
rect 958 728 962 732
rect 966 728 970 732
rect 1038 978 1042 982
rect 1110 948 1114 952
rect 1062 938 1066 942
rect 1094 938 1098 942
rect 1030 898 1034 902
rect 1054 908 1058 912
rect 1082 903 1086 907
rect 1089 903 1093 907
rect 1134 938 1138 942
rect 1174 938 1178 942
rect 1078 888 1082 892
rect 1046 878 1050 882
rect 1022 868 1026 872
rect 1086 868 1090 872
rect 1126 868 1130 872
rect 1366 1068 1370 1072
rect 1294 1058 1298 1062
rect 1278 1038 1282 1042
rect 1246 1028 1250 1032
rect 1446 1118 1450 1122
rect 1430 1098 1434 1102
rect 1430 1078 1434 1082
rect 1390 1059 1394 1063
rect 1438 1058 1442 1062
rect 1246 948 1250 952
rect 1206 938 1210 942
rect 1206 898 1210 902
rect 1142 888 1146 892
rect 1022 858 1026 862
rect 1118 858 1122 862
rect 1150 858 1154 862
rect 1006 848 1010 852
rect 1014 798 1018 802
rect 1006 738 1010 742
rect 982 708 986 712
rect 966 688 970 692
rect 990 698 994 702
rect 1038 738 1042 742
rect 1022 728 1026 732
rect 1014 668 1018 672
rect 982 658 986 662
rect 998 658 1002 662
rect 950 608 954 612
rect 902 588 906 592
rect 774 548 778 552
rect 798 558 802 562
rect 790 538 794 542
rect 814 528 818 532
rect 790 498 794 502
rect 750 468 754 472
rect 726 458 730 462
rect 750 458 754 462
rect 758 448 762 452
rect 702 348 706 352
rect 678 288 682 292
rect 518 258 522 262
rect 542 258 546 262
rect 686 278 690 282
rect 606 268 610 272
rect 654 268 658 272
rect 558 238 562 242
rect 510 218 514 222
rect 534 168 538 172
rect 638 228 642 232
rect 578 203 582 207
rect 585 203 589 207
rect 662 238 666 242
rect 822 488 826 492
rect 830 478 834 482
rect 782 468 786 472
rect 822 448 826 452
rect 990 618 994 622
rect 982 598 986 602
rect 990 558 994 562
rect 910 548 914 552
rect 1286 918 1290 922
rect 1318 918 1322 922
rect 1262 898 1266 902
rect 1302 888 1306 892
rect 1270 878 1274 882
rect 1270 868 1274 872
rect 1302 858 1306 862
rect 1166 848 1170 852
rect 1238 848 1242 852
rect 1150 828 1154 832
rect 1174 828 1178 832
rect 1086 758 1090 762
rect 1446 1048 1450 1052
rect 1470 1088 1474 1092
rect 1486 1108 1490 1112
rect 1478 1078 1482 1082
rect 1470 1068 1474 1072
rect 1422 968 1426 972
rect 1454 968 1458 972
rect 1462 968 1466 972
rect 1398 958 1402 962
rect 1406 948 1410 952
rect 1430 948 1434 952
rect 1398 938 1402 942
rect 1382 928 1386 932
rect 1374 828 1378 832
rect 1318 818 1322 822
rect 1358 818 1362 822
rect 1422 928 1426 932
rect 1438 928 1442 932
rect 1414 838 1418 842
rect 1502 1128 1506 1132
rect 1550 1128 1554 1132
rect 1534 1098 1538 1102
rect 1558 1098 1562 1102
rect 1582 1078 1586 1082
rect 1502 1058 1506 1062
rect 1550 1048 1554 1052
rect 1630 1138 1634 1142
rect 1638 1128 1642 1132
rect 1630 1088 1634 1092
rect 1630 1068 1634 1072
rect 1622 1058 1626 1062
rect 1602 1003 1606 1007
rect 1609 1003 1613 1007
rect 1614 978 1618 982
rect 1590 958 1594 962
rect 1582 948 1586 952
rect 1526 938 1530 942
rect 1462 888 1466 892
rect 1454 878 1458 882
rect 1110 748 1114 752
rect 1182 748 1186 752
rect 1198 748 1202 752
rect 1070 718 1074 722
rect 1158 718 1162 722
rect 1082 703 1086 707
rect 1089 703 1093 707
rect 1078 688 1082 692
rect 1118 668 1122 672
rect 1174 698 1178 702
rect 1366 748 1370 752
rect 1214 738 1218 742
rect 1246 738 1250 742
rect 1294 718 1298 722
rect 1206 708 1210 712
rect 1254 708 1258 712
rect 1230 698 1234 702
rect 1190 668 1194 672
rect 1054 658 1058 662
rect 1126 658 1130 662
rect 1046 648 1050 652
rect 1078 648 1082 652
rect 1054 638 1058 642
rect 1102 588 1106 592
rect 1142 648 1146 652
rect 1182 648 1186 652
rect 1174 628 1178 632
rect 1166 618 1170 622
rect 1086 578 1090 582
rect 1126 578 1130 582
rect 1030 568 1034 572
rect 1062 568 1066 572
rect 1030 558 1034 562
rect 1006 548 1010 552
rect 1022 548 1026 552
rect 934 518 938 522
rect 894 508 898 512
rect 878 488 882 492
rect 918 488 922 492
rect 894 478 898 482
rect 902 478 906 482
rect 838 458 842 462
rect 830 428 834 432
rect 822 398 826 402
rect 774 388 778 392
rect 782 368 786 372
rect 766 348 770 352
rect 926 478 930 482
rect 910 468 914 472
rect 942 508 946 512
rect 966 488 970 492
rect 1014 488 1018 492
rect 958 478 962 482
rect 990 478 994 482
rect 918 458 922 462
rect 934 458 938 462
rect 870 448 874 452
rect 958 448 962 452
rect 830 378 834 382
rect 862 378 866 382
rect 982 368 986 372
rect 854 358 858 362
rect 1030 468 1034 472
rect 822 348 826 352
rect 950 348 954 352
rect 990 348 994 352
rect 1014 348 1018 352
rect 1054 468 1058 472
rect 1054 448 1058 452
rect 1054 428 1058 432
rect 1046 388 1050 392
rect 726 318 730 322
rect 766 318 770 322
rect 726 288 730 292
rect 702 258 706 262
rect 710 258 714 262
rect 758 248 762 252
rect 718 238 722 242
rect 686 218 690 222
rect 678 178 682 182
rect 630 168 634 172
rect 590 158 594 162
rect 654 158 658 162
rect 694 168 698 172
rect 718 158 722 162
rect 638 148 642 152
rect 678 148 682 152
rect 702 148 706 152
rect 502 138 506 142
rect 606 138 610 142
rect 494 128 498 132
rect 398 118 402 122
rect 414 118 418 122
rect 470 118 474 122
rect 502 118 506 122
rect 526 118 530 122
rect 470 98 474 102
rect 262 88 266 92
rect 278 88 282 92
rect 438 88 442 92
rect 246 78 250 82
rect 342 78 346 82
rect 406 78 410 82
rect 502 78 506 82
rect 566 128 570 132
rect 582 98 586 102
rect 558 88 562 92
rect 526 68 530 72
rect 222 58 226 62
rect 382 58 386 62
rect 390 58 394 62
rect 630 138 634 142
rect 654 138 658 142
rect 686 138 690 142
rect 718 138 722 142
rect 678 128 682 132
rect 934 328 938 332
rect 950 318 954 322
rect 910 308 914 312
rect 838 288 842 292
rect 846 288 850 292
rect 926 278 930 282
rect 974 328 978 332
rect 990 328 994 332
rect 990 318 994 322
rect 982 308 986 312
rect 1038 328 1042 332
rect 1022 318 1026 322
rect 1038 318 1042 322
rect 1014 288 1018 292
rect 974 278 978 282
rect 1150 547 1154 551
rect 1126 538 1130 542
rect 1082 503 1086 507
rect 1089 503 1093 507
rect 1086 478 1090 482
rect 1086 448 1090 452
rect 1062 358 1066 362
rect 1110 458 1114 462
rect 1110 448 1114 452
rect 1206 658 1210 662
rect 1222 588 1226 592
rect 1254 678 1258 682
rect 1278 678 1282 682
rect 1238 668 1242 672
rect 1270 668 1274 672
rect 1270 658 1274 662
rect 1238 638 1242 642
rect 1270 638 1274 642
rect 1230 578 1234 582
rect 1278 608 1282 612
rect 1206 568 1210 572
rect 1238 568 1242 572
rect 1278 568 1282 572
rect 1230 558 1234 562
rect 1350 708 1354 712
rect 1390 718 1394 722
rect 1350 688 1354 692
rect 1382 688 1386 692
rect 1334 668 1338 672
rect 1294 638 1298 642
rect 1238 548 1242 552
rect 1254 548 1258 552
rect 1286 548 1290 552
rect 1198 538 1202 542
rect 1214 538 1218 542
rect 1270 538 1274 542
rect 1278 538 1282 542
rect 1278 528 1282 532
rect 1222 488 1226 492
rect 1190 478 1194 482
rect 1238 478 1242 482
rect 1270 478 1274 482
rect 1198 468 1202 472
rect 1214 438 1218 442
rect 1230 428 1234 432
rect 1278 468 1282 472
rect 1262 458 1266 462
rect 1302 618 1306 622
rect 1446 748 1450 752
rect 1638 1048 1642 1052
rect 1654 1118 1658 1122
rect 1806 1438 1810 1442
rect 1750 1348 1754 1352
rect 1758 1338 1762 1342
rect 1766 1328 1770 1332
rect 1830 1348 1834 1352
rect 1830 1338 1834 1342
rect 1806 1278 1810 1282
rect 1774 1268 1778 1272
rect 1742 1258 1746 1262
rect 1750 1248 1754 1252
rect 1686 1188 1690 1192
rect 1678 1158 1682 1162
rect 1734 1178 1738 1182
rect 1694 1148 1698 1152
rect 1742 1118 1746 1122
rect 1734 1108 1738 1112
rect 1710 1098 1714 1102
rect 1726 1088 1730 1092
rect 1710 1078 1714 1082
rect 1662 1068 1666 1072
rect 1670 1068 1674 1072
rect 1702 1068 1706 1072
rect 1654 1058 1658 1062
rect 1694 1058 1698 1062
rect 1718 1068 1722 1072
rect 1678 1048 1682 1052
rect 1710 1048 1714 1052
rect 1646 968 1650 972
rect 1638 948 1642 952
rect 1694 958 1698 962
rect 1742 1078 1746 1082
rect 1790 1258 1794 1262
rect 1782 1228 1786 1232
rect 1830 1268 1834 1272
rect 1838 1178 1842 1182
rect 1814 1168 1818 1172
rect 1822 1158 1826 1162
rect 1790 1148 1794 1152
rect 1806 1148 1810 1152
rect 1798 1138 1802 1142
rect 1838 1138 1842 1142
rect 1782 1128 1786 1132
rect 1766 1098 1770 1102
rect 1782 1098 1786 1102
rect 1774 1088 1778 1092
rect 1774 1068 1778 1072
rect 1838 1098 1842 1102
rect 1790 1088 1794 1092
rect 1830 1068 1834 1072
rect 1782 1058 1786 1062
rect 1750 1048 1754 1052
rect 1758 1038 1762 1042
rect 1822 1058 1826 1062
rect 1814 1048 1818 1052
rect 1822 1048 1826 1052
rect 1774 978 1778 982
rect 1750 968 1754 972
rect 1686 948 1690 952
rect 1718 948 1722 952
rect 1662 938 1666 942
rect 1550 928 1554 932
rect 1574 928 1578 932
rect 1622 928 1626 932
rect 1646 928 1650 932
rect 1598 888 1602 892
rect 1558 878 1562 882
rect 1590 878 1594 882
rect 1526 868 1530 872
rect 1526 838 1530 842
rect 1654 888 1658 892
rect 1622 878 1626 882
rect 1646 878 1650 882
rect 1614 868 1618 872
rect 1646 868 1650 872
rect 1606 858 1610 862
rect 1590 848 1594 852
rect 1602 803 1606 807
rect 1609 803 1613 807
rect 1614 758 1618 762
rect 1558 748 1562 752
rect 1606 748 1610 752
rect 1622 748 1626 752
rect 1638 748 1642 752
rect 1470 738 1474 742
rect 1510 738 1514 742
rect 1574 738 1578 742
rect 1438 728 1442 732
rect 1438 708 1442 712
rect 1406 698 1410 702
rect 1398 688 1402 692
rect 1446 688 1450 692
rect 1406 668 1410 672
rect 1446 668 1450 672
rect 1398 658 1402 662
rect 1454 658 1458 662
rect 1350 618 1354 622
rect 1318 598 1322 602
rect 1478 648 1482 652
rect 1422 588 1426 592
rect 1438 588 1442 592
rect 1454 578 1458 582
rect 1446 568 1450 572
rect 1478 568 1482 572
rect 1302 558 1306 562
rect 1462 558 1466 562
rect 1486 558 1490 562
rect 1294 528 1298 532
rect 1326 548 1330 552
rect 1342 548 1346 552
rect 1382 547 1386 551
rect 1438 548 1442 552
rect 1334 538 1338 542
rect 1406 538 1410 542
rect 1318 528 1322 532
rect 1334 528 1338 532
rect 1510 688 1514 692
rect 1566 698 1570 702
rect 1526 668 1530 672
rect 1550 668 1554 672
rect 1510 658 1514 662
rect 1558 648 1562 652
rect 1510 638 1514 642
rect 1542 558 1546 562
rect 1302 468 1306 472
rect 1406 468 1410 472
rect 1502 468 1506 472
rect 1286 458 1290 462
rect 1310 458 1314 462
rect 1254 448 1258 452
rect 1278 448 1282 452
rect 1302 448 1306 452
rect 1334 448 1338 452
rect 1350 448 1354 452
rect 1438 448 1442 452
rect 1246 428 1250 432
rect 1150 388 1154 392
rect 1238 388 1242 392
rect 1190 378 1194 382
rect 1206 358 1210 362
rect 1246 358 1250 362
rect 1190 348 1194 352
rect 1166 328 1170 332
rect 1102 318 1106 322
rect 1054 308 1058 312
rect 1046 278 1050 282
rect 998 268 1002 272
rect 1054 268 1058 272
rect 950 258 954 262
rect 782 248 786 252
rect 862 248 866 252
rect 894 248 898 252
rect 942 248 946 252
rect 934 238 938 242
rect 782 228 786 232
rect 918 228 922 232
rect 854 218 858 222
rect 894 208 898 212
rect 982 228 986 232
rect 1014 248 1018 252
rect 974 218 978 222
rect 1006 218 1010 222
rect 838 168 842 172
rect 822 158 826 162
rect 782 138 786 142
rect 750 118 754 122
rect 646 98 650 102
rect 638 88 642 92
rect 606 78 610 82
rect 670 88 674 92
rect 742 88 746 92
rect 750 78 754 82
rect 694 68 698 72
rect 806 128 810 132
rect 798 78 802 82
rect 774 68 778 72
rect 782 68 786 72
rect 870 158 874 162
rect 910 158 914 162
rect 926 148 930 152
rect 942 148 946 152
rect 950 148 954 152
rect 846 138 850 142
rect 846 128 850 132
rect 838 78 842 82
rect 822 68 826 72
rect 638 58 642 62
rect 702 58 706 62
rect 766 58 770 62
rect 814 58 818 62
rect 886 138 890 142
rect 902 128 906 132
rect 926 128 930 132
rect 942 128 946 132
rect 886 118 890 122
rect 870 108 874 112
rect 862 98 866 102
rect 894 98 898 102
rect 910 88 914 92
rect 942 88 946 92
rect 918 78 922 82
rect 854 68 858 72
rect 934 68 938 72
rect 862 58 866 62
rect 894 58 898 62
rect 942 58 946 62
rect 998 138 1002 142
rect 1022 138 1026 142
rect 982 128 986 132
rect 1014 128 1018 132
rect 982 108 986 112
rect 1082 303 1086 307
rect 1089 303 1093 307
rect 1222 348 1226 352
rect 1190 338 1194 342
rect 1214 338 1218 342
rect 1222 328 1226 332
rect 1246 338 1250 342
rect 1174 288 1178 292
rect 1222 288 1226 292
rect 1078 278 1082 282
rect 1086 278 1090 282
rect 1110 278 1114 282
rect 1230 278 1234 282
rect 1110 268 1114 272
rect 1070 258 1074 262
rect 1062 248 1066 252
rect 1150 248 1154 252
rect 1182 248 1186 252
rect 1118 238 1122 242
rect 1190 218 1194 222
rect 1102 158 1106 162
rect 1182 158 1186 162
rect 1118 148 1122 152
rect 1158 148 1162 152
rect 1110 138 1114 142
rect 1158 138 1162 142
rect 1054 128 1058 132
rect 1222 148 1226 152
rect 1230 138 1234 142
rect 1254 308 1258 312
rect 1262 288 1266 292
rect 1670 878 1674 882
rect 1670 758 1674 762
rect 1694 938 1698 942
rect 1694 918 1698 922
rect 1774 938 1778 942
rect 1726 928 1730 932
rect 1726 898 1730 902
rect 1830 948 1834 952
rect 1854 1488 1858 1492
rect 1862 1488 1866 1492
rect 1862 1468 1866 1472
rect 1862 1418 1866 1422
rect 1854 1348 1858 1352
rect 1902 1538 1906 1542
rect 1894 1518 1898 1522
rect 1878 1498 1882 1502
rect 1886 1458 1890 1462
rect 1878 1448 1882 1452
rect 1894 1448 1898 1452
rect 1870 1398 1874 1402
rect 1982 1538 1986 1542
rect 1990 1538 1994 1542
rect 2046 1538 2050 1542
rect 1982 1528 1986 1532
rect 1918 1518 1922 1522
rect 1934 1508 1938 1512
rect 1910 1468 1914 1472
rect 1982 1488 1986 1492
rect 1918 1458 1922 1462
rect 1958 1458 1962 1462
rect 1910 1438 1914 1442
rect 1878 1348 1882 1352
rect 1902 1348 1906 1352
rect 1854 1258 1858 1262
rect 1854 1248 1858 1252
rect 1854 1118 1858 1122
rect 1846 1088 1850 1092
rect 1894 1268 1898 1272
rect 1942 1448 1946 1452
rect 1926 1428 1930 1432
rect 2318 1747 2322 1751
rect 2398 1748 2402 1752
rect 2430 1748 2434 1752
rect 2542 1758 2546 1762
rect 2662 1758 2666 1762
rect 2222 1738 2226 1742
rect 2238 1738 2242 1742
rect 2254 1738 2258 1742
rect 2390 1738 2394 1742
rect 2406 1738 2410 1742
rect 2430 1738 2434 1742
rect 2470 1738 2474 1742
rect 2486 1738 2490 1742
rect 2270 1728 2274 1732
rect 2190 1718 2194 1722
rect 2206 1718 2210 1722
rect 2222 1718 2226 1722
rect 2246 1718 2250 1722
rect 2182 1688 2186 1692
rect 2102 1668 2106 1672
rect 2166 1668 2170 1672
rect 2086 1658 2090 1662
rect 2142 1658 2146 1662
rect 2158 1648 2162 1652
rect 2206 1698 2210 1702
rect 2230 1688 2234 1692
rect 2270 1688 2274 1692
rect 2422 1728 2426 1732
rect 2454 1728 2458 1732
rect 2390 1718 2394 1722
rect 2430 1718 2434 1722
rect 2462 1718 2466 1722
rect 2494 1728 2498 1732
rect 2502 1728 2506 1732
rect 2358 1688 2362 1692
rect 2390 1688 2394 1692
rect 2406 1688 2410 1692
rect 2454 1688 2458 1692
rect 2470 1688 2474 1692
rect 2478 1688 2482 1692
rect 2294 1678 2298 1682
rect 2270 1668 2274 1672
rect 2286 1668 2290 1672
rect 2318 1668 2322 1672
rect 2366 1668 2370 1672
rect 2406 1668 2410 1672
rect 2446 1668 2450 1672
rect 2198 1628 2202 1632
rect 2190 1618 2194 1622
rect 2198 1618 2202 1622
rect 2102 1608 2106 1612
rect 2118 1578 2122 1582
rect 2174 1568 2178 1572
rect 2358 1658 2362 1662
rect 2230 1648 2234 1652
rect 2278 1648 2282 1652
rect 2302 1648 2306 1652
rect 2310 1648 2314 1652
rect 2246 1618 2250 1622
rect 2294 1618 2298 1622
rect 2310 1618 2314 1622
rect 2294 1608 2298 1612
rect 2230 1598 2234 1602
rect 2222 1588 2226 1592
rect 2222 1568 2226 1572
rect 2158 1558 2162 1562
rect 2198 1558 2202 1562
rect 2142 1548 2146 1552
rect 2054 1528 2058 1532
rect 2070 1528 2074 1532
rect 2134 1528 2138 1532
rect 2106 1503 2110 1507
rect 2113 1503 2117 1507
rect 2190 1548 2194 1552
rect 2214 1548 2218 1552
rect 2182 1538 2186 1542
rect 2214 1538 2218 1542
rect 2342 1648 2346 1652
rect 2374 1648 2378 1652
rect 2398 1648 2402 1652
rect 2358 1638 2362 1642
rect 2382 1638 2386 1642
rect 2350 1578 2354 1582
rect 2278 1548 2282 1552
rect 2158 1528 2162 1532
rect 2182 1498 2186 1502
rect 2246 1498 2250 1502
rect 2142 1488 2146 1492
rect 2038 1478 2042 1482
rect 2086 1478 2090 1482
rect 2118 1478 2122 1482
rect 2126 1468 2130 1472
rect 2142 1468 2146 1472
rect 2086 1458 2090 1462
rect 2230 1488 2234 1492
rect 2294 1528 2298 1532
rect 2326 1528 2330 1532
rect 2270 1518 2274 1522
rect 2262 1488 2266 1492
rect 2254 1468 2258 1472
rect 2206 1458 2210 1462
rect 2214 1458 2218 1462
rect 2238 1458 2242 1462
rect 2166 1448 2170 1452
rect 2166 1438 2170 1442
rect 2102 1428 2106 1432
rect 2142 1418 2146 1422
rect 2014 1408 2018 1412
rect 2022 1398 2026 1402
rect 2078 1388 2082 1392
rect 1950 1378 1954 1382
rect 2014 1378 2018 1382
rect 1942 1368 1946 1372
rect 1990 1368 1994 1372
rect 1998 1368 2002 1372
rect 2062 1368 2066 1372
rect 2102 1368 2106 1372
rect 1958 1358 1962 1362
rect 2038 1358 2042 1362
rect 1966 1348 1970 1352
rect 1982 1348 1986 1352
rect 2030 1348 2034 1352
rect 1926 1338 1930 1342
rect 1942 1338 1946 1342
rect 1974 1338 1978 1342
rect 1910 1308 1914 1312
rect 1918 1308 1922 1312
rect 1942 1308 1946 1312
rect 1934 1288 1938 1292
rect 1918 1278 1922 1282
rect 1950 1278 1954 1282
rect 1934 1258 1938 1262
rect 2062 1348 2066 1352
rect 2014 1328 2018 1332
rect 1974 1258 1978 1262
rect 1894 1238 1898 1242
rect 1926 1238 1930 1242
rect 2022 1248 2026 1252
rect 1910 1168 1914 1172
rect 1918 1158 1922 1162
rect 1942 1158 1946 1162
rect 1918 1128 1922 1132
rect 1934 1128 1938 1132
rect 1894 1118 1898 1122
rect 1870 1108 1874 1112
rect 1910 1088 1914 1092
rect 1926 1078 1930 1082
rect 1958 1148 1962 1152
rect 2006 1148 2010 1152
rect 1910 1068 1914 1072
rect 1846 1058 1850 1062
rect 1814 928 1818 932
rect 1798 908 1802 912
rect 1838 908 1842 912
rect 1758 898 1762 902
rect 1718 878 1722 882
rect 1702 858 1706 862
rect 1830 888 1834 892
rect 1814 878 1818 882
rect 1822 878 1826 882
rect 1934 1048 1938 1052
rect 1878 1038 1882 1042
rect 1862 978 1866 982
rect 1918 978 1922 982
rect 1854 968 1858 972
rect 1870 968 1874 972
rect 1902 948 1906 952
rect 1862 928 1866 932
rect 1854 908 1858 912
rect 1894 938 1898 942
rect 1886 908 1890 912
rect 1870 898 1874 902
rect 1878 888 1882 892
rect 1902 888 1906 892
rect 1934 898 1938 902
rect 1958 1058 1962 1062
rect 1958 1048 1962 1052
rect 2078 1328 2082 1332
rect 2086 1328 2090 1332
rect 2190 1378 2194 1382
rect 2238 1448 2242 1452
rect 2286 1488 2290 1492
rect 2302 1488 2306 1492
rect 2294 1468 2298 1472
rect 2318 1458 2322 1462
rect 2334 1458 2338 1462
rect 2278 1448 2282 1452
rect 2286 1448 2290 1452
rect 2270 1438 2274 1442
rect 2278 1438 2282 1442
rect 2198 1368 2202 1372
rect 2286 1368 2290 1372
rect 2174 1348 2178 1352
rect 2198 1348 2202 1352
rect 2158 1338 2162 1342
rect 2118 1328 2122 1332
rect 2134 1328 2138 1332
rect 2150 1328 2154 1332
rect 2106 1303 2110 1307
rect 2113 1303 2117 1307
rect 2078 1278 2082 1282
rect 2086 1268 2090 1272
rect 2086 1258 2090 1262
rect 2070 1238 2074 1242
rect 2142 1278 2146 1282
rect 2110 1268 2114 1272
rect 2190 1328 2194 1332
rect 2182 1308 2186 1312
rect 2166 1278 2170 1282
rect 2126 1258 2130 1262
rect 2158 1258 2162 1262
rect 2246 1348 2250 1352
rect 2262 1338 2266 1342
rect 2222 1328 2226 1332
rect 2254 1318 2258 1322
rect 2238 1278 2242 1282
rect 2286 1328 2290 1332
rect 2270 1268 2274 1272
rect 2286 1268 2290 1272
rect 2230 1258 2234 1262
rect 2254 1258 2258 1262
rect 2278 1258 2282 1262
rect 2142 1248 2146 1252
rect 2246 1248 2250 1252
rect 2262 1248 2266 1252
rect 2166 1238 2170 1242
rect 2198 1238 2202 1242
rect 2222 1238 2226 1242
rect 2134 1218 2138 1222
rect 2102 1208 2106 1212
rect 2238 1208 2242 1212
rect 2222 1168 2226 1172
rect 2046 1158 2050 1162
rect 2078 1148 2082 1152
rect 2118 1148 2122 1152
rect 2038 1128 2042 1132
rect 2046 1118 2050 1122
rect 1974 1108 1978 1112
rect 1998 1108 2002 1112
rect 2014 1088 2018 1092
rect 2022 1078 2026 1082
rect 2030 1078 2034 1082
rect 2038 1078 2042 1082
rect 2054 1078 2058 1082
rect 2006 1048 2010 1052
rect 2046 1068 2050 1072
rect 2070 1098 2074 1102
rect 2094 1118 2098 1122
rect 2102 1118 2106 1122
rect 2106 1103 2110 1107
rect 2113 1103 2117 1107
rect 2086 1088 2090 1092
rect 2070 1068 2074 1072
rect 2062 1058 2066 1062
rect 2006 988 2010 992
rect 2038 988 2042 992
rect 2182 1148 2186 1152
rect 2246 1148 2250 1152
rect 2254 1148 2258 1152
rect 2158 1138 2162 1142
rect 2214 1138 2218 1142
rect 2230 1138 2234 1142
rect 2182 1128 2186 1132
rect 2206 1128 2210 1132
rect 2222 1108 2226 1112
rect 2214 1088 2218 1092
rect 2366 1558 2370 1562
rect 2494 1668 2498 1672
rect 2550 1748 2554 1752
rect 2590 1738 2594 1742
rect 2558 1728 2562 1732
rect 2526 1708 2530 1712
rect 2534 1688 2538 1692
rect 2558 1688 2562 1692
rect 2654 1728 2658 1732
rect 2670 1728 2674 1732
rect 2606 1718 2610 1722
rect 2574 1678 2578 1682
rect 2454 1658 2458 1662
rect 2470 1658 2474 1662
rect 2478 1658 2482 1662
rect 2414 1648 2418 1652
rect 2414 1638 2418 1642
rect 2438 1618 2442 1622
rect 2462 1618 2466 1622
rect 2518 1608 2522 1612
rect 2478 1578 2482 1582
rect 2462 1548 2466 1552
rect 2390 1508 2394 1512
rect 2358 1498 2362 1502
rect 2390 1498 2394 1502
rect 2398 1468 2402 1472
rect 2494 1568 2498 1572
rect 2550 1638 2554 1642
rect 2574 1658 2578 1662
rect 2638 1698 2642 1702
rect 2670 1688 2674 1692
rect 2590 1638 2594 1642
rect 2558 1598 2562 1602
rect 2590 1588 2594 1592
rect 2534 1558 2538 1562
rect 2542 1558 2546 1562
rect 2558 1558 2562 1562
rect 2574 1558 2578 1562
rect 2502 1548 2506 1552
rect 2542 1548 2546 1552
rect 2430 1528 2434 1532
rect 2422 1498 2426 1502
rect 2446 1498 2450 1502
rect 2526 1528 2530 1532
rect 2502 1518 2506 1522
rect 2510 1518 2514 1522
rect 2502 1508 2506 1512
rect 2518 1508 2522 1512
rect 2494 1498 2498 1502
rect 2486 1488 2490 1492
rect 2430 1468 2434 1472
rect 2446 1468 2450 1472
rect 2390 1458 2394 1462
rect 2406 1458 2410 1462
rect 2422 1458 2426 1462
rect 2302 1448 2306 1452
rect 2342 1448 2346 1452
rect 2374 1438 2378 1442
rect 2374 1378 2378 1382
rect 2334 1368 2338 1372
rect 2350 1368 2354 1372
rect 2326 1358 2330 1362
rect 2358 1348 2362 1352
rect 2406 1448 2410 1452
rect 2430 1448 2434 1452
rect 2462 1438 2466 1442
rect 2446 1428 2450 1432
rect 2422 1408 2426 1412
rect 2414 1388 2418 1392
rect 2422 1388 2426 1392
rect 2414 1368 2418 1372
rect 2406 1358 2410 1362
rect 2326 1338 2330 1342
rect 2310 1328 2314 1332
rect 2374 1328 2378 1332
rect 2302 1268 2306 1272
rect 2294 1178 2298 1182
rect 2390 1328 2394 1332
rect 2382 1318 2386 1322
rect 2318 1298 2322 1302
rect 2326 1288 2330 1292
rect 2350 1288 2354 1292
rect 2358 1278 2362 1282
rect 2334 1268 2338 1272
rect 2342 1208 2346 1212
rect 2382 1268 2386 1272
rect 2366 1258 2370 1262
rect 2382 1248 2386 1252
rect 2358 1238 2362 1242
rect 2398 1308 2402 1312
rect 2398 1258 2402 1262
rect 2406 1238 2410 1242
rect 2382 1228 2386 1232
rect 2390 1228 2394 1232
rect 2350 1168 2354 1172
rect 2294 1158 2298 1162
rect 2310 1158 2314 1162
rect 2366 1158 2370 1162
rect 2302 1148 2306 1152
rect 2358 1148 2362 1152
rect 2286 1138 2290 1142
rect 2310 1138 2314 1142
rect 2350 1138 2354 1142
rect 2262 1128 2266 1132
rect 2238 1088 2242 1092
rect 2158 1078 2162 1082
rect 2166 1078 2170 1082
rect 2094 1068 2098 1072
rect 2182 1068 2186 1072
rect 2246 1068 2250 1072
rect 2270 1068 2274 1072
rect 2118 1058 2122 1062
rect 2158 1058 2162 1062
rect 2206 1058 2210 1062
rect 2222 1058 2226 1062
rect 2174 1048 2178 1052
rect 2070 1038 2074 1042
rect 2230 1038 2234 1042
rect 2206 988 2210 992
rect 2054 968 2058 972
rect 2062 968 2066 972
rect 2110 968 2114 972
rect 2046 958 2050 962
rect 2094 958 2098 962
rect 2070 948 2074 952
rect 1950 918 1954 922
rect 2006 938 2010 942
rect 2014 928 2018 932
rect 2022 928 2026 932
rect 1966 908 1970 912
rect 2006 898 2010 902
rect 1974 878 1978 882
rect 1982 878 1986 882
rect 1990 878 1994 882
rect 1846 868 1850 872
rect 1854 868 1858 872
rect 1918 868 1922 872
rect 1942 868 1946 872
rect 1814 858 1818 862
rect 2022 868 2026 872
rect 1950 858 1954 862
rect 1798 848 1802 852
rect 1846 848 1850 852
rect 1958 848 1962 852
rect 1798 798 1802 802
rect 1686 748 1690 752
rect 1646 738 1650 742
rect 1734 738 1738 742
rect 1662 728 1666 732
rect 1710 728 1714 732
rect 1590 618 1594 622
rect 1602 603 1606 607
rect 1609 603 1613 607
rect 1590 588 1594 592
rect 1630 598 1634 602
rect 1622 548 1626 552
rect 1566 528 1570 532
rect 1582 528 1586 532
rect 1574 498 1578 502
rect 1598 498 1602 502
rect 1534 438 1538 442
rect 1454 368 1458 372
rect 1390 358 1394 362
rect 1398 358 1402 362
rect 1382 348 1386 352
rect 1294 338 1298 342
rect 1318 308 1322 312
rect 1302 298 1306 302
rect 1294 288 1298 292
rect 1254 258 1258 262
rect 1286 258 1290 262
rect 1310 288 1314 292
rect 1574 358 1578 362
rect 1558 348 1562 352
rect 1342 338 1346 342
rect 1406 338 1410 342
rect 1518 338 1522 342
rect 1542 338 1546 342
rect 1326 298 1330 302
rect 1334 288 1338 292
rect 1318 268 1322 272
rect 1366 328 1370 332
rect 1390 328 1394 332
rect 1414 328 1418 332
rect 1358 308 1362 312
rect 1630 418 1634 422
rect 1602 403 1606 407
rect 1609 403 1613 407
rect 1654 678 1658 682
rect 1654 588 1658 592
rect 1694 708 1698 712
rect 1814 768 1818 772
rect 1830 768 1834 772
rect 1942 838 1946 842
rect 1958 838 1962 842
rect 1990 838 1994 842
rect 1998 838 2002 842
rect 1950 818 1954 822
rect 1886 808 1890 812
rect 1990 808 1994 812
rect 1854 768 1858 772
rect 1910 768 1914 772
rect 1942 768 1946 772
rect 1814 748 1818 752
rect 1846 748 1850 752
rect 1782 738 1786 742
rect 1790 728 1794 732
rect 1750 718 1754 722
rect 1758 718 1762 722
rect 1774 718 1778 722
rect 1734 678 1738 682
rect 1766 678 1770 682
rect 1758 668 1762 672
rect 1678 588 1682 592
rect 1670 548 1674 552
rect 1662 538 1666 542
rect 1702 538 1706 542
rect 1702 508 1706 512
rect 1790 668 1794 672
rect 1846 738 1850 742
rect 1862 738 1866 742
rect 1894 738 1898 742
rect 1822 708 1826 712
rect 1918 748 1922 752
rect 1934 748 1938 752
rect 2014 768 2018 772
rect 1998 748 2002 752
rect 1958 738 1962 742
rect 1870 728 1874 732
rect 1838 668 1842 672
rect 1862 668 1866 672
rect 1910 698 1914 702
rect 2062 938 2066 942
rect 2094 938 2098 942
rect 2158 948 2162 952
rect 2238 978 2242 982
rect 2318 1108 2322 1112
rect 2294 1088 2298 1092
rect 2302 1088 2306 1092
rect 2342 1098 2346 1102
rect 2318 1078 2322 1082
rect 2342 1078 2346 1082
rect 2414 1148 2418 1152
rect 2390 1128 2394 1132
rect 2614 1578 2618 1582
rect 2590 1538 2594 1542
rect 2606 1528 2610 1532
rect 2678 1608 2682 1612
rect 2646 1558 2650 1562
rect 2694 1558 2698 1562
rect 2622 1518 2626 1522
rect 2646 1538 2650 1542
rect 2686 1538 2690 1542
rect 2542 1498 2546 1502
rect 2614 1498 2618 1502
rect 2638 1498 2642 1502
rect 2510 1488 2514 1492
rect 2534 1488 2538 1492
rect 2574 1478 2578 1482
rect 2582 1478 2586 1482
rect 2534 1468 2538 1472
rect 2542 1468 2546 1472
rect 2590 1468 2594 1472
rect 2638 1488 2642 1492
rect 2630 1468 2634 1472
rect 2646 1468 2650 1472
rect 2526 1458 2530 1462
rect 2582 1458 2586 1462
rect 2614 1458 2618 1462
rect 2654 1458 2658 1462
rect 2510 1448 2514 1452
rect 2518 1448 2522 1452
rect 2550 1448 2554 1452
rect 2566 1398 2570 1402
rect 2550 1378 2554 1382
rect 2470 1368 2474 1372
rect 2478 1368 2482 1372
rect 2494 1368 2498 1372
rect 2462 1358 2466 1362
rect 2510 1358 2514 1362
rect 2614 1418 2618 1422
rect 2622 1398 2626 1402
rect 2662 1388 2666 1392
rect 2590 1378 2594 1382
rect 2582 1358 2586 1362
rect 2606 1358 2610 1362
rect 2662 1358 2666 1362
rect 2462 1348 2466 1352
rect 2486 1348 2490 1352
rect 2502 1348 2506 1352
rect 2518 1348 2522 1352
rect 2534 1348 2538 1352
rect 2478 1338 2482 1342
rect 2462 1328 2466 1332
rect 2454 1318 2458 1322
rect 2430 1288 2434 1292
rect 2470 1278 2474 1282
rect 2454 1258 2458 1262
rect 2430 1238 2434 1242
rect 2438 1238 2442 1242
rect 2430 1198 2434 1202
rect 2566 1338 2570 1342
rect 2542 1328 2546 1332
rect 2502 1318 2506 1322
rect 2526 1318 2530 1322
rect 2550 1308 2554 1312
rect 2534 1288 2538 1292
rect 2598 1348 2602 1352
rect 2622 1338 2626 1342
rect 2662 1338 2666 1342
rect 2590 1328 2594 1332
rect 2606 1328 2610 1332
rect 2630 1328 2634 1332
rect 2646 1328 2650 1332
rect 2574 1308 2578 1312
rect 2574 1298 2578 1302
rect 2622 1298 2626 1302
rect 2558 1288 2562 1292
rect 2598 1288 2602 1292
rect 2630 1278 2634 1282
rect 2494 1268 2498 1272
rect 2494 1258 2498 1262
rect 2582 1248 2586 1252
rect 2510 1228 2514 1232
rect 2622 1268 2626 1272
rect 2646 1268 2650 1272
rect 2590 1208 2594 1212
rect 2486 1198 2490 1202
rect 2686 1488 2690 1492
rect 2702 1488 2706 1492
rect 2686 1478 2690 1482
rect 2686 1458 2690 1462
rect 2678 1338 2682 1342
rect 2702 1268 2706 1272
rect 2662 1258 2666 1262
rect 2550 1188 2554 1192
rect 2526 1178 2530 1182
rect 2470 1158 2474 1162
rect 2462 1148 2466 1152
rect 2486 1148 2490 1152
rect 2478 1138 2482 1142
rect 2510 1138 2514 1142
rect 2534 1158 2538 1162
rect 2542 1158 2546 1162
rect 2558 1168 2562 1172
rect 2582 1158 2586 1162
rect 2670 1158 2674 1162
rect 2630 1148 2634 1152
rect 2702 1148 2706 1152
rect 2582 1138 2586 1142
rect 2598 1138 2602 1142
rect 2622 1138 2626 1142
rect 2662 1138 2666 1142
rect 2454 1128 2458 1132
rect 2502 1128 2506 1132
rect 2566 1128 2570 1132
rect 2310 1058 2314 1062
rect 2302 998 2306 1002
rect 2254 958 2258 962
rect 2278 958 2282 962
rect 2222 948 2226 952
rect 2134 928 2138 932
rect 2150 918 2154 922
rect 2106 903 2110 907
rect 2113 903 2117 907
rect 2150 898 2154 902
rect 2062 878 2066 882
rect 2070 868 2074 872
rect 2078 858 2082 862
rect 2126 858 2130 862
rect 2054 848 2058 852
rect 2086 848 2090 852
rect 2046 838 2050 842
rect 2038 828 2042 832
rect 2046 798 2050 802
rect 2086 808 2090 812
rect 2054 768 2058 772
rect 2078 758 2082 762
rect 2054 748 2058 752
rect 2022 738 2026 742
rect 2062 738 2066 742
rect 2078 738 2082 742
rect 2030 728 2034 732
rect 2046 728 2050 732
rect 1958 708 1962 712
rect 2022 718 2026 722
rect 2038 708 2042 712
rect 2022 698 2026 702
rect 1942 688 1946 692
rect 1902 668 1906 672
rect 1918 668 1922 672
rect 1934 668 1938 672
rect 1806 658 1810 662
rect 1758 568 1762 572
rect 1806 568 1810 572
rect 1726 558 1730 562
rect 1790 558 1794 562
rect 1862 658 1866 662
rect 1886 658 1890 662
rect 1918 658 1922 662
rect 1926 598 1930 602
rect 1990 658 1994 662
rect 2062 698 2066 702
rect 2054 688 2058 692
rect 2094 758 2098 762
rect 2134 747 2138 751
rect 2182 918 2186 922
rect 2198 878 2202 882
rect 2310 968 2314 972
rect 2334 1058 2338 1062
rect 2350 1058 2354 1062
rect 2398 1038 2402 1042
rect 2422 1118 2426 1122
rect 2470 1118 2474 1122
rect 2430 1108 2434 1112
rect 2438 1108 2442 1112
rect 2462 1108 2466 1112
rect 2358 958 2362 962
rect 2406 958 2410 962
rect 2486 1088 2490 1092
rect 2470 1058 2474 1062
rect 2478 1058 2482 1062
rect 2438 1008 2442 1012
rect 2470 998 2474 1002
rect 2462 968 2466 972
rect 2398 948 2402 952
rect 2414 948 2418 952
rect 2334 938 2338 942
rect 2350 938 2354 942
rect 2374 938 2378 942
rect 2390 938 2394 942
rect 2214 868 2218 872
rect 2230 868 2234 872
rect 2182 858 2186 862
rect 2198 828 2202 832
rect 2182 818 2186 822
rect 2174 738 2178 742
rect 2110 728 2114 732
rect 2158 728 2162 732
rect 2094 718 2098 722
rect 2086 688 2090 692
rect 2106 703 2110 707
rect 2113 703 2117 707
rect 2366 928 2370 932
rect 2382 928 2386 932
rect 2310 918 2314 922
rect 2262 888 2266 892
rect 2254 878 2258 882
rect 2246 868 2250 872
rect 2294 898 2298 902
rect 2318 908 2322 912
rect 2374 908 2378 912
rect 2494 1028 2498 1032
rect 2502 968 2506 972
rect 2494 958 2498 962
rect 2486 938 2490 942
rect 2414 928 2418 932
rect 2270 878 2274 882
rect 2318 878 2322 882
rect 2366 878 2370 882
rect 2430 898 2434 902
rect 2430 888 2434 892
rect 2454 888 2458 892
rect 2462 878 2466 882
rect 2278 868 2282 872
rect 2342 858 2346 862
rect 2390 858 2394 862
rect 2318 848 2322 852
rect 2342 838 2346 842
rect 2222 768 2226 772
rect 2238 768 2242 772
rect 2198 718 2202 722
rect 2206 718 2210 722
rect 2198 698 2202 702
rect 2198 678 2202 682
rect 2262 748 2266 752
rect 2230 738 2234 742
rect 2270 738 2274 742
rect 2238 708 2242 712
rect 2446 858 2450 862
rect 2422 788 2426 792
rect 2454 838 2458 842
rect 2446 778 2450 782
rect 2382 758 2386 762
rect 2406 758 2410 762
rect 2438 758 2442 762
rect 2294 748 2298 752
rect 2326 748 2330 752
rect 2342 748 2346 752
rect 2366 748 2370 752
rect 2302 738 2306 742
rect 2374 738 2378 742
rect 2598 1108 2602 1112
rect 2558 1098 2562 1102
rect 2526 1088 2530 1092
rect 2606 1078 2610 1082
rect 2638 1078 2642 1082
rect 2702 1078 2706 1082
rect 2614 1068 2618 1072
rect 2662 1068 2666 1072
rect 2558 1058 2562 1062
rect 2646 1058 2650 1062
rect 2606 1048 2610 1052
rect 2550 1038 2554 1042
rect 2630 1038 2634 1042
rect 2670 1038 2674 1042
rect 2582 1018 2586 1022
rect 2558 988 2562 992
rect 2646 968 2650 972
rect 2558 958 2562 962
rect 2510 908 2514 912
rect 2510 888 2514 892
rect 2622 938 2626 942
rect 2550 928 2554 932
rect 2590 918 2594 922
rect 2654 908 2658 912
rect 2606 888 2610 892
rect 2638 888 2642 892
rect 2686 898 2690 902
rect 2558 868 2562 872
rect 2534 858 2538 862
rect 2566 858 2570 862
rect 2582 858 2586 862
rect 2518 848 2522 852
rect 2486 798 2490 802
rect 2542 828 2546 832
rect 2526 788 2530 792
rect 2478 768 2482 772
rect 2550 758 2554 762
rect 2390 748 2394 752
rect 2398 738 2402 742
rect 2406 738 2410 742
rect 2518 738 2522 742
rect 2294 718 2298 722
rect 2390 718 2394 722
rect 2286 708 2290 712
rect 2342 708 2346 712
rect 2374 698 2378 702
rect 2246 688 2250 692
rect 2270 688 2274 692
rect 2326 688 2330 692
rect 2142 668 2146 672
rect 2230 668 2234 672
rect 2118 658 2122 662
rect 2134 658 2138 662
rect 2158 658 2162 662
rect 1942 588 1946 592
rect 1830 568 1834 572
rect 1910 568 1914 572
rect 1862 558 1866 562
rect 1774 548 1778 552
rect 1782 548 1786 552
rect 1814 548 1818 552
rect 2334 668 2338 672
rect 2358 668 2362 672
rect 2198 658 2202 662
rect 2118 638 2122 642
rect 2150 638 2154 642
rect 1734 538 1738 542
rect 1742 538 1746 542
rect 1758 528 1762 532
rect 1734 518 1738 522
rect 1766 518 1770 522
rect 1718 478 1722 482
rect 1718 459 1722 463
rect 2062 548 2066 552
rect 2102 548 2106 552
rect 1806 538 1810 542
rect 1814 538 1818 542
rect 1806 518 1810 522
rect 1758 488 1762 492
rect 2054 538 2058 542
rect 1878 508 1882 512
rect 1894 508 1898 512
rect 1958 508 1962 512
rect 1982 508 1986 512
rect 1998 508 2002 512
rect 1870 478 1874 482
rect 1942 478 1946 482
rect 1742 458 1746 462
rect 1894 448 1898 452
rect 1926 448 1930 452
rect 1742 438 1746 442
rect 1646 368 1650 372
rect 1590 348 1594 352
rect 1566 318 1570 322
rect 1526 308 1530 312
rect 1454 298 1458 302
rect 1390 278 1394 282
rect 1350 268 1354 272
rect 1406 268 1410 272
rect 1534 288 1538 292
rect 1494 278 1498 282
rect 1510 278 1514 282
rect 1574 278 1578 282
rect 1526 268 1530 272
rect 1366 258 1370 262
rect 1518 258 1522 262
rect 1758 418 1762 422
rect 1734 358 1738 362
rect 2054 518 2058 522
rect 2182 548 2186 552
rect 2286 658 2290 662
rect 2294 658 2298 662
rect 2294 618 2298 622
rect 2310 618 2314 622
rect 2374 658 2378 662
rect 2366 648 2370 652
rect 2358 638 2362 642
rect 2358 618 2362 622
rect 2350 588 2354 592
rect 2286 548 2290 552
rect 2310 548 2314 552
rect 2166 538 2170 542
rect 2118 528 2122 532
rect 2190 518 2194 522
rect 2070 508 2074 512
rect 2106 503 2110 507
rect 2113 503 2117 507
rect 2430 728 2434 732
rect 2406 718 2410 722
rect 2430 718 2434 722
rect 2486 718 2490 722
rect 2438 698 2442 702
rect 2422 678 2426 682
rect 2494 678 2498 682
rect 2454 668 2458 672
rect 2478 668 2482 672
rect 2414 658 2418 662
rect 2486 658 2490 662
rect 2486 628 2490 632
rect 2446 618 2450 622
rect 2398 588 2402 592
rect 2406 568 2410 572
rect 2430 568 2434 572
rect 2510 668 2514 672
rect 2566 848 2570 852
rect 2622 828 2626 832
rect 2566 798 2570 802
rect 2574 778 2578 782
rect 2598 778 2602 782
rect 2590 758 2594 762
rect 2606 768 2610 772
rect 2686 788 2690 792
rect 2654 758 2658 762
rect 2670 758 2674 762
rect 2638 748 2642 752
rect 2662 748 2666 752
rect 2638 738 2642 742
rect 2558 728 2562 732
rect 2590 728 2594 732
rect 2630 728 2634 732
rect 2670 718 2674 722
rect 2654 708 2658 712
rect 2678 708 2682 712
rect 2566 688 2570 692
rect 2550 678 2554 682
rect 2574 678 2578 682
rect 2630 668 2634 672
rect 2502 648 2506 652
rect 2526 648 2530 652
rect 2518 638 2522 642
rect 2622 588 2626 592
rect 2614 568 2618 572
rect 2598 558 2602 562
rect 2606 548 2610 552
rect 2622 548 2626 552
rect 2446 538 2450 542
rect 2390 528 2394 532
rect 2302 518 2306 522
rect 2294 508 2298 512
rect 2278 488 2282 492
rect 2334 488 2338 492
rect 2062 478 2066 482
rect 1990 468 1994 472
rect 2014 468 2018 472
rect 2126 468 2130 472
rect 2030 458 2034 462
rect 2094 458 2098 462
rect 2150 458 2154 462
rect 1814 358 1818 362
rect 1878 358 1882 362
rect 1894 358 1898 362
rect 1918 358 1922 362
rect 1718 348 1722 352
rect 1742 348 1746 352
rect 1774 348 1778 352
rect 1798 348 1802 352
rect 1638 338 1642 342
rect 1670 338 1674 342
rect 1686 338 1690 342
rect 1886 338 1890 342
rect 1918 338 1922 342
rect 1774 328 1778 332
rect 1918 328 1922 332
rect 1934 328 1938 332
rect 1614 318 1618 322
rect 1702 318 1706 322
rect 1302 248 1306 252
rect 1358 248 1362 252
rect 1470 248 1474 252
rect 1534 248 1538 252
rect 1566 248 1570 252
rect 1382 238 1386 242
rect 1430 218 1434 222
rect 1310 158 1314 162
rect 1374 158 1378 162
rect 1382 148 1386 152
rect 1574 158 1578 162
rect 1478 148 1482 152
rect 1550 148 1554 152
rect 1374 138 1378 142
rect 1470 138 1474 142
rect 1486 138 1490 142
rect 1134 128 1138 132
rect 1190 128 1194 132
rect 1230 128 1234 132
rect 1246 128 1250 132
rect 1366 128 1370 132
rect 1550 128 1554 132
rect 1110 118 1114 122
rect 1046 108 1050 112
rect 1082 103 1086 107
rect 1089 103 1093 107
rect 1174 118 1178 122
rect 1206 118 1210 122
rect 1102 98 1106 102
rect 1126 98 1130 102
rect 1166 98 1170 102
rect 1054 88 1058 92
rect 1110 88 1114 92
rect 982 78 986 82
rect 1006 78 1010 82
rect 1030 78 1034 82
rect 1038 78 1042 82
rect 966 68 970 72
rect 982 68 986 72
rect 998 68 1002 72
rect 1022 68 1026 72
rect 1246 98 1250 102
rect 1158 88 1162 92
rect 1166 78 1170 82
rect 1214 78 1218 82
rect 1230 78 1234 82
rect 1054 68 1058 72
rect 1110 68 1114 72
rect 1014 58 1018 62
rect 1030 58 1034 62
rect 1174 58 1178 62
rect 1182 58 1186 62
rect 1206 58 1210 62
rect 30 48 34 52
rect 86 48 90 52
rect 150 48 154 52
rect 278 48 282 52
rect 438 48 442 52
rect 830 48 834 52
rect 870 48 874 52
rect 958 48 962 52
rect 1134 48 1138 52
rect 1166 48 1170 52
rect 1326 118 1330 122
rect 1254 88 1258 92
rect 1302 88 1306 92
rect 1342 88 1346 92
rect 1254 78 1258 82
rect 1414 118 1418 122
rect 1398 88 1402 92
rect 1318 78 1322 82
rect 1350 78 1354 82
rect 1366 78 1370 82
rect 1310 68 1314 72
rect 1374 68 1378 72
rect 1438 108 1442 112
rect 1510 98 1514 102
rect 1534 98 1538 102
rect 1630 298 1634 302
rect 1662 298 1666 302
rect 1750 298 1754 302
rect 1654 278 1658 282
rect 1862 308 1866 312
rect 1782 298 1786 302
rect 1678 278 1682 282
rect 1822 278 1826 282
rect 1718 268 1722 272
rect 1638 258 1642 262
rect 1614 218 1618 222
rect 1602 203 1606 207
rect 1609 203 1613 207
rect 1670 248 1674 252
rect 1822 258 1826 262
rect 1814 248 1818 252
rect 1790 238 1794 242
rect 1694 158 1698 162
rect 1766 158 1770 162
rect 2022 388 2026 392
rect 1974 368 1978 372
rect 2254 458 2258 462
rect 2174 388 2178 392
rect 2046 358 2050 362
rect 2062 358 2066 362
rect 2118 358 2122 362
rect 2038 348 2042 352
rect 2062 348 2066 352
rect 2086 348 2090 352
rect 2006 338 2010 342
rect 2102 328 2106 332
rect 2190 328 2194 332
rect 2054 318 2058 322
rect 1942 278 1946 282
rect 2326 448 2330 452
rect 2318 388 2322 392
rect 2510 528 2514 532
rect 2574 538 2578 542
rect 2582 538 2586 542
rect 2598 538 2602 542
rect 2606 528 2610 532
rect 2438 518 2442 522
rect 2518 518 2522 522
rect 2550 518 2554 522
rect 2454 478 2458 482
rect 2430 468 2434 472
rect 2358 448 2362 452
rect 2390 448 2394 452
rect 2422 448 2426 452
rect 2334 368 2338 372
rect 2294 358 2298 362
rect 2342 348 2346 352
rect 2246 338 2250 342
rect 2318 338 2322 342
rect 2230 328 2234 332
rect 2310 328 2314 332
rect 2158 308 2162 312
rect 2198 308 2202 312
rect 2106 303 2110 307
rect 2113 303 2117 307
rect 2046 288 2050 292
rect 1902 268 1906 272
rect 1926 268 1930 272
rect 2014 268 2018 272
rect 1878 158 1882 162
rect 1734 148 1738 152
rect 1830 148 1834 152
rect 1886 148 1890 152
rect 1630 138 1634 142
rect 1798 138 1802 142
rect 1622 128 1626 132
rect 1694 128 1698 132
rect 1590 98 1594 102
rect 1542 88 1546 92
rect 1526 78 1530 82
rect 1646 98 1650 102
rect 1702 88 1706 92
rect 1702 58 1706 62
rect 1222 48 1226 52
rect 1270 48 1274 52
rect 1358 48 1362 52
rect 1382 48 1386 52
rect 1422 48 1426 52
rect 222 38 226 42
rect 1542 38 1546 42
rect 526 8 530 12
rect 550 8 554 12
rect 838 8 842 12
rect 578 3 582 7
rect 585 3 589 7
rect 1602 3 1606 7
rect 1609 3 1613 7
rect 1846 138 1850 142
rect 1758 98 1762 102
rect 1814 98 1818 102
rect 1718 88 1722 92
rect 1846 78 1850 82
rect 1774 58 1778 62
rect 1878 108 1882 112
rect 1902 108 1906 112
rect 1910 98 1914 102
rect 2078 278 2082 282
rect 2102 278 2106 282
rect 2174 278 2178 282
rect 2086 268 2090 272
rect 2006 258 2010 262
rect 1982 158 1986 162
rect 2006 158 2010 162
rect 1926 148 1930 152
rect 1998 148 2002 152
rect 1950 138 1954 142
rect 1966 138 1970 142
rect 1950 128 1954 132
rect 1894 88 1898 92
rect 1942 78 1946 82
rect 1982 78 1986 82
rect 1910 68 1914 72
rect 1982 68 1986 72
rect 2070 238 2074 242
rect 2070 188 2074 192
rect 2054 168 2058 172
rect 2094 248 2098 252
rect 2118 248 2122 252
rect 2198 268 2202 272
rect 2142 238 2146 242
rect 2110 228 2114 232
rect 2214 258 2218 262
rect 2166 238 2170 242
rect 2150 178 2154 182
rect 2182 178 2186 182
rect 2094 168 2098 172
rect 2062 148 2066 152
rect 2078 148 2082 152
rect 2110 148 2114 152
rect 2038 138 2042 142
rect 2054 138 2058 142
rect 2102 128 2106 132
rect 2182 148 2186 152
rect 2142 138 2146 142
rect 2134 118 2138 122
rect 2106 103 2110 107
rect 2113 103 2117 107
rect 2054 98 2058 102
rect 2358 328 2362 332
rect 2254 318 2258 322
rect 2366 308 2370 312
rect 2398 368 2402 372
rect 2598 508 2602 512
rect 2550 488 2554 492
rect 2558 488 2562 492
rect 2502 478 2506 482
rect 2510 478 2514 482
rect 2534 468 2538 472
rect 2486 458 2490 462
rect 2510 458 2514 462
rect 2502 448 2506 452
rect 2526 448 2530 452
rect 2534 448 2538 452
rect 2502 428 2506 432
rect 2462 358 2466 362
rect 2470 348 2474 352
rect 2382 298 2386 302
rect 2422 338 2426 342
rect 2422 318 2426 322
rect 2462 338 2466 342
rect 2446 328 2450 332
rect 2406 298 2410 302
rect 2430 298 2434 302
rect 2334 288 2338 292
rect 2390 288 2394 292
rect 2294 278 2298 282
rect 2310 278 2314 282
rect 2326 278 2330 282
rect 2374 278 2378 282
rect 2270 268 2274 272
rect 2294 268 2298 272
rect 2262 258 2266 262
rect 2278 258 2282 262
rect 2246 188 2250 192
rect 2230 168 2234 172
rect 2230 148 2234 152
rect 2238 148 2242 152
rect 2198 138 2202 142
rect 2166 128 2170 132
rect 2246 128 2250 132
rect 2158 108 2162 112
rect 2214 98 2218 102
rect 2182 88 2186 92
rect 2222 78 2226 82
rect 2238 78 2242 82
rect 2038 68 2042 72
rect 2134 68 2138 72
rect 2374 258 2378 262
rect 2374 248 2378 252
rect 2382 248 2386 252
rect 2278 168 2282 172
rect 2310 168 2314 172
rect 2270 138 2274 142
rect 2286 138 2290 142
rect 2294 128 2298 132
rect 2342 228 2346 232
rect 2446 288 2450 292
rect 2486 278 2490 282
rect 2566 478 2570 482
rect 2542 378 2546 382
rect 2590 458 2594 462
rect 2558 448 2562 452
rect 2590 418 2594 422
rect 2558 398 2562 402
rect 2590 378 2594 382
rect 2582 358 2586 362
rect 2558 338 2562 342
rect 2566 308 2570 312
rect 2590 298 2594 302
rect 2542 288 2546 292
rect 2574 288 2578 292
rect 2662 668 2666 672
rect 2662 538 2666 542
rect 2670 528 2674 532
rect 2654 498 2658 502
rect 2678 498 2682 502
rect 2614 428 2618 432
rect 2614 398 2618 402
rect 2694 558 2698 562
rect 2694 478 2698 482
rect 2614 358 2618 362
rect 2678 358 2682 362
rect 2622 348 2626 352
rect 2606 338 2610 342
rect 2630 338 2634 342
rect 2638 318 2642 322
rect 2542 278 2546 282
rect 2574 278 2578 282
rect 2430 268 2434 272
rect 2550 268 2554 272
rect 2350 168 2354 172
rect 2406 168 2410 172
rect 2358 148 2362 152
rect 2398 148 2402 152
rect 2374 128 2378 132
rect 2342 108 2346 112
rect 2334 98 2338 102
rect 2270 88 2274 92
rect 2294 78 2298 82
rect 2278 68 2282 72
rect 2318 68 2322 72
rect 1958 58 1962 62
rect 2022 58 2026 62
rect 2158 58 2162 62
rect 2438 258 2442 262
rect 2462 258 2466 262
rect 2430 238 2434 242
rect 2446 238 2450 242
rect 2414 138 2418 142
rect 2422 128 2426 132
rect 2414 98 2418 102
rect 2414 88 2418 92
rect 2486 248 2490 252
rect 2518 248 2522 252
rect 2558 218 2562 222
rect 2614 258 2618 262
rect 2478 188 2482 192
rect 2502 188 2506 192
rect 2470 148 2474 152
rect 2486 148 2490 152
rect 2510 178 2514 182
rect 2518 158 2522 162
rect 2526 148 2530 152
rect 2590 148 2594 152
rect 2462 138 2466 142
rect 2566 138 2570 142
rect 2486 128 2490 132
rect 2454 68 2458 72
rect 2526 128 2530 132
rect 2550 118 2554 122
rect 2550 108 2554 112
rect 2534 98 2538 102
rect 2574 98 2578 102
rect 2574 88 2578 92
rect 2622 88 2626 92
rect 2510 78 2514 82
rect 2526 78 2530 82
rect 2566 78 2570 82
rect 2590 78 2594 82
rect 2502 68 2506 72
rect 2638 268 2642 272
rect 2638 158 2642 162
rect 2654 318 2658 322
rect 2702 468 2706 472
rect 2662 278 2666 282
rect 2678 118 2682 122
rect 2686 118 2690 122
rect 2638 78 2642 82
rect 2286 58 2290 62
rect 2334 58 2338 62
rect 2358 58 2362 62
rect 2398 58 2402 62
rect 2422 58 2426 62
rect 2518 58 2522 62
rect 2550 58 2554 62
rect 2558 58 2562 62
rect 2694 108 2698 112
rect 2686 88 2690 92
rect 1718 48 1722 52
rect 1862 48 1866 52
rect 1974 48 1978 52
rect 2006 48 2010 52
rect 2070 48 2074 52
rect 2462 48 2466 52
rect 2606 48 2610 52
rect 2614 48 2618 52
rect 2654 48 2658 52
<< metal3 >>
rect 576 1803 578 1807
rect 582 1803 585 1807
rect 590 1803 592 1807
rect 1600 1803 1602 1807
rect 1606 1803 1609 1807
rect 1614 1803 1616 1807
rect 450 1798 454 1801
rect 794 1798 838 1801
rect 1738 1798 1782 1801
rect 742 1792 745 1798
rect 742 1778 758 1781
rect 770 1778 782 1781
rect 2026 1778 2158 1781
rect 2162 1778 2502 1781
rect 742 1772 745 1778
rect 1842 1768 1870 1771
rect 18 1758 54 1761
rect 98 1758 102 1761
rect 898 1758 934 1761
rect 2054 1761 2057 1768
rect 2054 1758 2086 1761
rect 2222 1761 2225 1768
rect 2222 1758 2382 1761
rect 2546 1758 2662 1761
rect -26 1748 -22 1752
rect 582 1748 654 1751
rect 842 1748 910 1751
rect 922 1748 926 1751
rect 1066 1748 1070 1751
rect 1146 1748 1294 1751
rect 1546 1748 1654 1751
rect 1658 1748 1662 1751
rect 1842 1748 2190 1751
rect 2202 1748 2230 1751
rect 2242 1748 2246 1751
rect 2282 1748 2318 1751
rect 582 1742 585 1748
rect 2402 1748 2430 1751
rect 2554 1748 2593 1751
rect 2590 1742 2593 1748
rect 66 1738 86 1741
rect 266 1738 302 1741
rect 378 1738 398 1741
rect 402 1738 446 1741
rect 450 1738 502 1741
rect 922 1738 993 1741
rect 1018 1738 1198 1741
rect 1210 1738 1270 1741
rect 1610 1738 1670 1741
rect 1722 1738 1854 1741
rect 1994 1738 1998 1741
rect 2178 1738 2190 1741
rect 2226 1738 2230 1741
rect 2242 1738 2254 1741
rect 2394 1738 2406 1741
rect 2434 1738 2470 1741
rect 2474 1738 2486 1741
rect -26 1731 -22 1732
rect 6 1731 9 1738
rect -26 1728 54 1731
rect 158 1731 161 1738
rect 990 1732 993 1738
rect 2006 1732 2009 1738
rect 158 1728 214 1731
rect 218 1728 238 1731
rect 242 1728 246 1731
rect 386 1728 406 1731
rect 410 1728 454 1731
rect 1650 1728 1750 1731
rect 1778 1728 1838 1731
rect 2058 1728 2270 1731
rect 2426 1728 2454 1731
rect 2498 1728 2502 1731
rect 2538 1728 2558 1731
rect 2658 1728 2670 1731
rect 2734 1728 2738 1732
rect 138 1718 142 1721
rect 198 1718 206 1721
rect 210 1718 270 1721
rect 274 1718 302 1721
rect 498 1718 526 1721
rect 530 1718 622 1721
rect 1082 1718 1118 1721
rect 1210 1718 1294 1721
rect 1298 1718 1334 1721
rect 1402 1718 1406 1721
rect 1410 1718 1470 1721
rect 1750 1721 1753 1728
rect 1750 1718 1910 1721
rect 2042 1718 2158 1721
rect 2194 1718 2206 1721
rect 2226 1718 2246 1721
rect 2394 1718 2430 1721
rect 2454 1718 2462 1721
rect 2466 1718 2606 1721
rect 122 1708 142 1711
rect 1122 1708 1166 1711
rect 2034 1708 2070 1711
rect 2194 1708 2526 1711
rect 1080 1703 1082 1707
rect 1086 1703 1089 1707
rect 1094 1703 1096 1707
rect 2104 1703 2106 1707
rect 2110 1703 2113 1707
rect 2118 1703 2120 1707
rect -26 1698 -22 1702
rect 1938 1698 2062 1701
rect 2146 1698 2150 1701
rect 2162 1698 2206 1701
rect 2226 1698 2638 1701
rect 1066 1688 1150 1691
rect 1214 1691 1217 1698
rect 1214 1688 1254 1691
rect 1258 1688 1310 1691
rect 1538 1688 1542 1691
rect 1722 1688 1806 1691
rect 2010 1688 2086 1691
rect 2090 1688 2182 1691
rect 2234 1688 2270 1691
rect 2350 1688 2358 1691
rect 2362 1688 2390 1691
rect 2398 1688 2406 1691
rect 2410 1688 2446 1691
rect 2458 1688 2470 1691
rect 2482 1688 2534 1691
rect 2562 1688 2574 1691
rect 2674 1688 2702 1691
rect 2734 1691 2738 1692
rect 2706 1688 2738 1691
rect -26 1678 -22 1682
rect 322 1678 350 1681
rect 434 1678 470 1681
rect 474 1678 510 1681
rect 682 1678 726 1681
rect 730 1678 886 1681
rect 1210 1678 1334 1681
rect 1338 1678 1342 1681
rect 2074 1678 2294 1681
rect 2298 1678 2574 1681
rect 66 1668 110 1671
rect 202 1668 310 1671
rect 362 1668 422 1671
rect 450 1668 454 1671
rect 530 1668 550 1671
rect 570 1668 614 1671
rect 898 1668 974 1671
rect 1078 1671 1081 1678
rect 1042 1668 1081 1671
rect 1538 1668 1582 1671
rect 1734 1671 1737 1678
rect 1586 1668 1737 1671
rect 2106 1668 2166 1671
rect 2274 1668 2286 1671
rect 2322 1668 2326 1671
rect 2370 1668 2406 1671
rect 2410 1668 2446 1671
rect 2450 1668 2494 1671
rect 2734 1668 2738 1672
rect -26 1658 -22 1662
rect 58 1658 118 1661
rect 178 1658 190 1661
rect 242 1658 254 1661
rect 298 1658 326 1661
rect 506 1658 534 1661
rect 538 1658 582 1661
rect 722 1658 806 1661
rect 826 1658 926 1661
rect 930 1658 982 1661
rect 1014 1661 1017 1668
rect 1014 1659 1102 1661
rect 1278 1661 1281 1668
rect 1014 1658 1105 1659
rect 1278 1658 1326 1661
rect 1418 1658 1478 1661
rect 1522 1658 1598 1661
rect 1750 1661 1753 1668
rect 1706 1658 1753 1661
rect 1842 1658 1910 1661
rect 2090 1658 2142 1661
rect 2278 1658 2305 1661
rect 2362 1658 2454 1661
rect 2466 1658 2470 1661
rect 2482 1658 2574 1661
rect 2278 1652 2281 1658
rect 2302 1652 2305 1658
rect 386 1648 550 1651
rect 626 1648 726 1651
rect 914 1648 998 1651
rect 1586 1648 1678 1651
rect 1682 1648 1822 1651
rect 1850 1648 1982 1651
rect 1994 1648 2158 1651
rect 2162 1648 2230 1651
rect 2314 1648 2342 1651
rect 2366 1648 2374 1651
rect 2386 1648 2398 1651
rect 2410 1648 2414 1651
rect -26 1638 -22 1642
rect 134 1641 137 1648
rect 2382 1642 2385 1648
rect 106 1638 137 1641
rect 434 1638 478 1641
rect 618 1638 646 1641
rect 650 1638 686 1641
rect 690 1638 734 1641
rect 738 1638 846 1641
rect 850 1638 1022 1641
rect 1026 1638 1190 1641
rect 1194 1638 1366 1641
rect 1370 1638 1382 1641
rect 1882 1638 2038 1641
rect 2042 1638 2358 1641
rect 2418 1638 2550 1641
rect 2554 1638 2590 1641
rect 2734 1638 2738 1642
rect 994 1628 1262 1631
rect 1266 1628 1342 1631
rect 1346 1628 1398 1631
rect 2002 1628 2198 1631
rect 714 1618 750 1621
rect 890 1618 1206 1621
rect 1330 1618 1422 1621
rect 1906 1618 2190 1621
rect 2202 1618 2246 1621
rect 2250 1618 2294 1621
rect 2298 1618 2310 1621
rect 2442 1618 2462 1621
rect 1938 1608 2102 1611
rect 2298 1608 2518 1611
rect 2522 1608 2662 1611
rect 2666 1608 2678 1611
rect 576 1603 578 1607
rect 582 1603 585 1607
rect 590 1603 592 1607
rect 1600 1603 1602 1607
rect 1606 1603 1609 1607
rect 1614 1603 1616 1607
rect 2234 1598 2558 1601
rect -26 1588 -22 1592
rect 138 1588 166 1591
rect 2226 1588 2334 1591
rect 2338 1588 2590 1591
rect 82 1578 142 1581
rect 266 1578 350 1581
rect 474 1578 502 1581
rect 1962 1578 2118 1581
rect 2122 1578 2350 1581
rect 2482 1578 2614 1581
rect -26 1568 -22 1572
rect 170 1568 206 1571
rect 298 1568 358 1571
rect 1358 1568 1510 1571
rect 1602 1568 1718 1571
rect 1914 1568 1998 1571
rect 2178 1568 2222 1571
rect 142 1562 145 1568
rect 42 1558 46 1561
rect 298 1558 334 1561
rect 354 1558 390 1561
rect 494 1561 497 1568
rect 494 1558 566 1561
rect 1014 1561 1017 1568
rect 1358 1562 1361 1568
rect 1002 1558 1017 1561
rect 1030 1558 1038 1561
rect 1042 1558 1174 1561
rect 1410 1558 1502 1561
rect 1506 1558 1550 1561
rect 1730 1558 1798 1561
rect 1826 1558 1838 1561
rect 1842 1558 2158 1561
rect 2162 1558 2198 1561
rect 2214 1558 2281 1561
rect -26 1551 -22 1552
rect -26 1548 30 1551
rect 34 1548 78 1551
rect 138 1548 142 1551
rect 218 1548 246 1551
rect 330 1548 366 1551
rect 370 1548 406 1551
rect 506 1548 510 1551
rect 646 1551 649 1558
rect 634 1548 649 1551
rect 874 1548 894 1551
rect 898 1548 926 1551
rect 930 1548 942 1551
rect 946 1548 1070 1551
rect 1074 1548 1094 1551
rect 1338 1548 1358 1551
rect 1362 1548 1366 1551
rect 1654 1551 1657 1558
rect 2214 1552 2217 1558
rect 2278 1552 2281 1558
rect 2494 1561 2497 1568
rect 2494 1558 2534 1561
rect 2546 1558 2558 1561
rect 2578 1558 2646 1561
rect 2650 1558 2694 1561
rect 1374 1548 1446 1551
rect 742 1542 745 1548
rect 1374 1542 1377 1548
rect 1654 1548 1686 1551
rect 1738 1548 1918 1551
rect 1994 1548 2049 1551
rect 2146 1548 2190 1551
rect 2366 1551 2369 1558
rect 2366 1548 2462 1551
rect 2506 1548 2542 1551
rect 194 1538 238 1541
rect 242 1538 278 1541
rect 306 1538 382 1541
rect 786 1538 862 1541
rect 914 1538 1350 1541
rect 1426 1538 1526 1541
rect 1530 1538 1582 1541
rect 1714 1538 1766 1541
rect 1786 1538 1798 1541
rect 1934 1541 1937 1548
rect 2046 1542 2049 1548
rect 1906 1538 1937 1541
rect 1986 1538 1990 1541
rect 2186 1538 2214 1541
rect 2594 1538 2646 1541
rect 2682 1538 2686 1541
rect 258 1528 390 1531
rect 418 1528 430 1531
rect 754 1528 774 1531
rect 954 1528 998 1531
rect 1010 1528 1030 1531
rect 1034 1528 1046 1531
rect 1082 1528 1118 1531
rect 1202 1528 1294 1531
rect 1298 1528 1470 1531
rect 1474 1528 1518 1531
rect 1698 1528 1846 1531
rect 1850 1528 1982 1531
rect 1986 1528 2054 1531
rect 2058 1528 2070 1531
rect 2138 1528 2158 1531
rect 2298 1528 2326 1531
rect 2418 1528 2430 1531
rect 2530 1528 2606 1531
rect 2510 1522 2513 1528
rect 34 1518 158 1521
rect 610 1518 702 1521
rect 986 1518 1062 1521
rect 1066 1518 1086 1521
rect 1338 1518 1366 1521
rect 1738 1518 1766 1521
rect 1802 1518 1822 1521
rect 1898 1518 1918 1521
rect 2274 1518 2502 1521
rect 2546 1518 2622 1521
rect -26 1508 -22 1512
rect 1274 1508 1398 1511
rect 1754 1508 1782 1511
rect 1786 1508 1934 1511
rect 1938 1508 1998 1511
rect 2386 1508 2390 1511
rect 2506 1508 2518 1511
rect 1080 1503 1082 1507
rect 1086 1503 1089 1507
rect 1094 1503 1096 1507
rect 2104 1503 2106 1507
rect 2110 1503 2113 1507
rect 2118 1503 2120 1507
rect 58 1498 246 1501
rect 442 1498 534 1501
rect 1122 1498 1150 1501
rect 1818 1498 1878 1501
rect 2186 1498 2246 1501
rect 2362 1498 2390 1501
rect 2394 1498 2422 1501
rect 2426 1498 2446 1501
rect 2450 1498 2494 1501
rect 2498 1498 2542 1501
rect 2618 1498 2638 1501
rect 10 1488 86 1491
rect 106 1488 166 1491
rect 510 1488 518 1491
rect 522 1488 678 1491
rect 730 1488 854 1491
rect 938 1488 942 1491
rect 1002 1488 1118 1491
rect 1810 1488 1822 1491
rect 1842 1488 1854 1491
rect 1986 1488 2142 1491
rect 2234 1488 2262 1491
rect 2266 1488 2286 1491
rect 2306 1488 2486 1491
rect 2514 1488 2534 1491
rect 2642 1488 2686 1491
rect 2690 1488 2697 1491
rect 294 1482 297 1488
rect 58 1478 126 1481
rect 186 1478 238 1481
rect 438 1481 441 1488
rect 438 1478 502 1481
rect 634 1478 670 1481
rect 1050 1478 1094 1481
rect 1130 1478 1206 1481
rect 1210 1478 1222 1481
rect 1714 1478 1726 1481
rect 1730 1478 1806 1481
rect 1862 1481 1865 1488
rect 1810 1478 1865 1481
rect 2042 1478 2086 1481
rect 2122 1478 2158 1481
rect 2162 1478 2574 1481
rect 2578 1478 2582 1481
rect 2702 1481 2705 1488
rect 2690 1478 2705 1481
rect 42 1468 102 1471
rect 278 1471 281 1478
rect 234 1468 281 1471
rect 442 1468 574 1471
rect 578 1468 630 1471
rect 822 1471 825 1478
rect 870 1471 873 1478
rect 822 1468 873 1471
rect 954 1468 998 1471
rect 1106 1468 1190 1471
rect 1194 1468 1198 1471
rect 1354 1468 1382 1471
rect 1386 1468 1438 1471
rect 1442 1468 1534 1471
rect 1794 1468 1857 1471
rect 1866 1468 1886 1471
rect 1914 1468 2121 1471
rect 2130 1468 2134 1471
rect 2146 1468 2254 1471
rect 2298 1468 2398 1471
rect 2426 1468 2430 1471
rect 2450 1468 2534 1471
rect 2546 1468 2590 1471
rect 2634 1468 2646 1471
rect -26 1458 -22 1462
rect 42 1458 46 1461
rect 214 1461 217 1468
rect 82 1458 217 1461
rect 514 1458 558 1461
rect 774 1461 777 1468
rect 698 1458 777 1461
rect 842 1458 870 1461
rect 890 1458 958 1461
rect 1050 1458 1070 1461
rect 1154 1458 1174 1461
rect 1410 1458 1414 1461
rect 1426 1458 1430 1461
rect 1438 1458 1446 1461
rect 1450 1458 1526 1461
rect 1666 1458 1734 1461
rect 1818 1458 1830 1461
rect 1854 1461 1857 1468
rect 1854 1458 1886 1461
rect 1922 1458 1945 1461
rect 1962 1458 2086 1461
rect 2118 1461 2121 1468
rect 2118 1458 2206 1461
rect 2218 1458 2238 1461
rect 2242 1458 2289 1461
rect 2322 1458 2334 1461
rect 2394 1458 2406 1461
rect 2426 1458 2510 1461
rect 2514 1458 2526 1461
rect 2586 1458 2614 1461
rect 2618 1458 2654 1461
rect 2658 1458 2686 1461
rect 1942 1452 1945 1458
rect 2286 1452 2289 1458
rect 66 1448 78 1451
rect 98 1448 110 1451
rect 146 1448 174 1451
rect 546 1448 726 1451
rect 858 1448 974 1451
rect 978 1448 1038 1451
rect 1130 1448 1278 1451
rect 1602 1448 1790 1451
rect 1882 1448 1894 1451
rect 1950 1448 2166 1451
rect 2170 1448 2238 1451
rect 2250 1448 2278 1451
rect 2306 1448 2342 1451
rect 2410 1448 2430 1451
rect 2522 1448 2550 1451
rect 362 1438 406 1441
rect 466 1438 550 1441
rect 554 1438 622 1441
rect 838 1441 841 1448
rect 746 1438 841 1441
rect 890 1438 902 1441
rect 906 1438 1166 1441
rect 1778 1438 1806 1441
rect 1810 1438 1902 1441
rect 1950 1441 1953 1448
rect 1914 1438 1953 1441
rect 2170 1438 2270 1441
rect 2282 1438 2374 1441
rect 2510 1441 2513 1448
rect 2466 1438 2513 1441
rect 1186 1428 1286 1431
rect 1930 1428 2102 1431
rect 874 1418 1598 1421
rect 1642 1418 1758 1421
rect 1866 1418 2006 1421
rect 2446 1421 2449 1428
rect 2146 1418 2449 1421
rect 2586 1418 2614 1421
rect 2018 1408 2422 1411
rect 390 1402 393 1408
rect 576 1403 578 1407
rect 582 1403 585 1407
rect 590 1403 592 1407
rect 1600 1403 1602 1407
rect 1606 1403 1609 1407
rect 1614 1403 1616 1407
rect 746 1398 750 1401
rect 1362 1398 1438 1401
rect 1762 1398 1766 1401
rect 1874 1398 2022 1401
rect 2570 1398 2622 1401
rect 266 1388 342 1391
rect 386 1388 502 1391
rect 506 1388 862 1391
rect 1234 1388 1318 1391
rect 1322 1388 1374 1391
rect 1762 1388 2006 1391
rect 2010 1388 2078 1391
rect 2190 1388 2246 1391
rect 2250 1388 2414 1391
rect 2426 1388 2662 1391
rect 2190 1382 2193 1388
rect 18 1378 286 1381
rect 290 1378 310 1381
rect 842 1378 878 1381
rect 1082 1378 1182 1381
rect 1954 1378 2014 1381
rect 2378 1378 2550 1381
rect 2554 1378 2582 1381
rect 170 1368 254 1371
rect 1114 1368 1206 1371
rect 1778 1368 1782 1371
rect 1786 1368 1942 1371
rect 1994 1368 1998 1371
rect 2106 1368 2198 1371
rect 2290 1368 2334 1371
rect 2354 1368 2414 1371
rect 2418 1368 2470 1371
rect 2474 1368 2478 1371
rect 2590 1371 2593 1378
rect 2498 1368 2593 1371
rect 270 1362 273 1368
rect 154 1358 158 1361
rect 162 1358 174 1361
rect 178 1358 190 1361
rect 298 1358 334 1361
rect 502 1361 505 1368
rect 502 1358 558 1361
rect 1010 1358 1030 1361
rect 1034 1358 1126 1361
rect 1698 1358 1766 1361
rect 1770 1358 1958 1361
rect 1962 1358 2038 1361
rect 2062 1361 2065 1368
rect 2286 1361 2289 1368
rect 2062 1358 2289 1361
rect 2330 1358 2406 1361
rect 2410 1358 2414 1361
rect 2454 1358 2462 1361
rect 2466 1358 2510 1361
rect 2586 1358 2606 1361
rect -26 1348 -22 1352
rect 74 1348 102 1351
rect 106 1348 118 1351
rect 130 1348 150 1351
rect 170 1348 206 1351
rect 242 1348 270 1351
rect 274 1348 294 1351
rect 358 1348 366 1351
rect 422 1351 425 1358
rect 2662 1352 2665 1358
rect 370 1348 425 1351
rect 578 1348 662 1351
rect 682 1348 793 1351
rect 930 1348 1118 1351
rect 1178 1348 1238 1351
rect 1354 1348 1422 1351
rect 1586 1348 1750 1351
rect 1834 1348 1854 1351
rect 1858 1348 1878 1351
rect 1906 1348 1966 1351
rect 1970 1348 1982 1351
rect 2066 1348 2174 1351
rect 2178 1348 2198 1351
rect 2202 1348 2246 1351
rect 2258 1348 2358 1351
rect 2362 1348 2422 1351
rect 2466 1348 2486 1351
rect 2506 1348 2518 1351
rect -26 1341 -23 1348
rect -26 1338 134 1341
rect 518 1341 521 1348
rect 486 1338 521 1341
rect 790 1342 793 1348
rect 850 1338 990 1341
rect 994 1338 1614 1341
rect 1618 1338 1678 1341
rect 1762 1338 1766 1341
rect 1810 1338 1830 1341
rect 1834 1338 1926 1341
rect 1946 1338 1974 1341
rect 2030 1341 2033 1348
rect 2030 1338 2086 1341
rect 2162 1338 2262 1341
rect 2306 1338 2326 1341
rect 2342 1338 2478 1341
rect 2534 1341 2537 1348
rect 2534 1338 2566 1341
rect 2598 1341 2601 1348
rect 2598 1338 2622 1341
rect 2666 1338 2678 1341
rect 2734 1338 2738 1342
rect 486 1332 489 1338
rect 2342 1332 2345 1338
rect 2462 1332 2465 1338
rect 26 1328 70 1331
rect 106 1328 318 1331
rect 394 1328 486 1331
rect 514 1328 526 1331
rect 954 1328 982 1331
rect 1042 1328 1070 1331
rect 1122 1328 1174 1331
rect 1186 1328 1198 1331
rect 1666 1328 1766 1331
rect 1770 1328 2014 1331
rect 2018 1328 2070 1331
rect 2074 1328 2078 1331
rect 2090 1328 2118 1331
rect 2154 1328 2190 1331
rect 2226 1328 2254 1331
rect 2290 1328 2310 1331
rect 2378 1328 2390 1331
rect 2526 1328 2542 1331
rect 2594 1328 2606 1331
rect 2626 1328 2630 1331
rect 2634 1328 2646 1331
rect 2650 1328 2702 1331
rect 394 1318 582 1321
rect 1010 1318 1038 1321
rect 1042 1318 1142 1321
rect 1146 1318 1182 1321
rect 1282 1318 1342 1321
rect 1570 1318 1590 1321
rect 2134 1321 2137 1328
rect 2526 1322 2529 1328
rect 2058 1318 2137 1321
rect 2258 1318 2382 1321
rect 2458 1318 2502 1321
rect 390 1312 393 1318
rect 58 1308 118 1311
rect 122 1308 126 1311
rect 202 1308 262 1311
rect 890 1308 1054 1311
rect 1914 1308 1918 1311
rect 1922 1308 1942 1311
rect 2186 1308 2302 1311
rect 2402 1308 2550 1311
rect 2554 1308 2574 1311
rect 1080 1303 1082 1307
rect 1086 1303 1089 1307
rect 1094 1303 1096 1307
rect 2104 1303 2106 1307
rect 2110 1303 2113 1307
rect 2118 1303 2120 1307
rect 2318 1302 2321 1308
rect 226 1298 246 1301
rect 2326 1298 2430 1301
rect 2578 1298 2622 1301
rect 2326 1292 2329 1298
rect -26 1288 -22 1292
rect 18 1288 46 1291
rect 50 1288 70 1291
rect 426 1288 494 1291
rect 498 1288 622 1291
rect 626 1288 726 1291
rect 1066 1288 1118 1291
rect 1250 1288 1286 1291
rect 1594 1288 1614 1291
rect 1938 1288 2326 1291
rect 2354 1288 2430 1291
rect 238 1281 241 1288
rect 238 1278 262 1281
rect 290 1278 302 1281
rect 330 1278 342 1281
rect 382 1281 385 1288
rect 1134 1282 1137 1288
rect 354 1278 385 1281
rect 442 1278 526 1281
rect 530 1278 534 1281
rect 634 1278 750 1281
rect 1002 1278 1054 1281
rect 1146 1278 1158 1281
rect 1210 1278 1238 1281
rect 1242 1278 1254 1281
rect 1482 1278 1502 1281
rect 1530 1278 1534 1281
rect 1586 1278 1590 1281
rect 1746 1278 1806 1281
rect 1810 1278 1918 1281
rect 1922 1278 1950 1281
rect 1954 1278 2078 1281
rect 2082 1278 2142 1281
rect 2170 1278 2174 1281
rect 2362 1278 2470 1281
rect 2534 1281 2537 1288
rect 2558 1281 2561 1288
rect 2534 1278 2561 1281
rect 2598 1281 2601 1288
rect 2598 1278 2630 1281
rect 66 1268 126 1271
rect 130 1268 182 1271
rect 186 1268 246 1271
rect 314 1268 358 1271
rect 362 1268 374 1271
rect 378 1268 422 1271
rect 790 1271 793 1278
rect 754 1268 793 1271
rect 838 1268 934 1271
rect 990 1270 1006 1271
rect 74 1258 86 1261
rect 186 1258 190 1261
rect 302 1261 305 1268
rect 302 1258 342 1261
rect 346 1258 542 1261
rect 562 1258 574 1261
rect 646 1261 649 1268
rect 662 1261 665 1268
rect 838 1262 841 1268
rect 994 1268 1006 1270
rect 1138 1268 1198 1271
rect 1262 1271 1265 1278
rect 1202 1268 1265 1271
rect 1302 1271 1305 1278
rect 2238 1272 2241 1278
rect 1274 1268 1305 1271
rect 1338 1268 1406 1271
rect 1466 1268 1470 1271
rect 1778 1268 1830 1271
rect 1834 1268 1894 1271
rect 1898 1268 2086 1271
rect 2090 1268 2110 1271
rect 2274 1268 2286 1271
rect 2306 1268 2334 1271
rect 2386 1268 2494 1271
rect 2626 1268 2646 1271
rect 2682 1268 2702 1271
rect 2734 1271 2738 1272
rect 2706 1268 2738 1271
rect 646 1258 665 1261
rect 770 1258 798 1261
rect 1114 1258 1190 1261
rect 1194 1258 1254 1261
rect 1386 1258 1454 1261
rect 1458 1258 1470 1261
rect 1474 1258 1526 1261
rect 1746 1258 1790 1261
rect 1794 1258 1854 1261
rect 1938 1258 1974 1261
rect 2022 1258 2054 1261
rect 2130 1258 2158 1261
rect 2162 1258 2230 1261
rect 2234 1258 2254 1261
rect 2282 1258 2366 1261
rect 2402 1258 2406 1261
rect 2410 1258 2454 1261
rect 2498 1258 2662 1261
rect -26 1251 -22 1252
rect -26 1248 54 1251
rect 166 1251 169 1258
rect 2022 1252 2025 1258
rect 166 1248 214 1251
rect 274 1248 390 1251
rect 414 1248 470 1251
rect 978 1248 1014 1251
rect 1138 1248 1142 1251
rect 1178 1248 1286 1251
rect 1290 1248 1390 1251
rect 1514 1248 1582 1251
rect 1754 1248 1854 1251
rect 2086 1251 2089 1258
rect 2086 1248 2142 1251
rect 2146 1248 2246 1251
rect 2250 1248 2262 1251
rect 2386 1248 2433 1251
rect 414 1242 417 1248
rect 242 1238 270 1241
rect 490 1238 694 1241
rect 814 1241 817 1248
rect 2430 1242 2433 1248
rect 2438 1248 2582 1251
rect 2734 1248 2738 1252
rect 2438 1242 2441 1248
rect 698 1238 817 1241
rect 1162 1238 1169 1241
rect 1218 1238 1262 1241
rect 1266 1238 1406 1241
rect 1410 1238 1422 1241
rect 1426 1238 1566 1241
rect 1898 1238 1926 1241
rect 2074 1238 2166 1241
rect 2202 1238 2214 1241
rect 2226 1238 2230 1241
rect 2354 1238 2358 1241
rect 1166 1232 1169 1238
rect 186 1228 318 1231
rect 354 1228 654 1231
rect 970 1228 974 1231
rect 978 1228 1134 1231
rect 1290 1228 1398 1231
rect 1402 1228 1446 1231
rect 1450 1228 1486 1231
rect 1786 1228 2174 1231
rect 2178 1228 2382 1231
rect 2386 1228 2390 1231
rect 2406 1231 2409 1238
rect 2406 1228 2510 1231
rect 434 1218 462 1221
rect 466 1218 606 1221
rect 826 1218 846 1221
rect 850 1218 918 1221
rect 2138 1218 2326 1221
rect 1058 1208 1214 1211
rect 2106 1208 2238 1211
rect 2346 1208 2590 1211
rect 576 1203 578 1207
rect 582 1203 585 1207
rect 590 1203 592 1207
rect 1600 1203 1602 1207
rect 1606 1203 1609 1207
rect 1614 1203 1616 1207
rect 954 1198 1214 1201
rect 1330 1198 1414 1201
rect 1418 1198 1446 1201
rect 2306 1198 2430 1201
rect 2482 1198 2486 1201
rect 746 1188 1590 1191
rect 1602 1188 1686 1191
rect 2434 1188 2550 1191
rect 1018 1178 1358 1181
rect 1362 1178 1526 1181
rect 1530 1178 1550 1181
rect 1738 1178 1838 1181
rect 1842 1178 2294 1181
rect 2298 1178 2526 1181
rect -26 1171 -22 1172
rect -26 1168 6 1171
rect 10 1168 166 1171
rect 302 1171 305 1178
rect 302 1168 350 1171
rect 426 1168 502 1171
rect 506 1168 558 1171
rect 562 1168 702 1171
rect 738 1168 750 1171
rect 1066 1168 1286 1171
rect 1306 1168 1310 1171
rect 1818 1168 1862 1171
rect 1914 1168 1942 1171
rect 1946 1168 2222 1171
rect 2226 1168 2350 1171
rect 2354 1168 2390 1171
rect 2410 1168 2558 1171
rect 298 1158 334 1161
rect 834 1158 854 1161
rect 858 1158 902 1161
rect 1066 1158 1086 1161
rect 1342 1161 1345 1168
rect 1342 1158 1358 1161
rect 1518 1161 1521 1168
rect 1498 1158 1534 1161
rect 1682 1158 1822 1161
rect 1826 1158 1918 1161
rect 1946 1158 2046 1161
rect 2182 1158 2294 1161
rect 2314 1158 2366 1161
rect 2426 1158 2470 1161
rect 2586 1158 2670 1161
rect -26 1148 -22 1152
rect 210 1148 238 1151
rect 390 1151 393 1158
rect 2182 1152 2185 1158
rect 342 1148 393 1151
rect 546 1148 598 1151
rect 754 1148 758 1151
rect 890 1148 926 1151
rect 310 1142 313 1148
rect 342 1142 345 1148
rect 1002 1148 1126 1151
rect 1130 1148 1174 1151
rect 1302 1148 1334 1151
rect 1354 1148 1502 1151
rect 1698 1148 1790 1151
rect 1810 1148 1814 1151
rect 2082 1148 2118 1151
rect 2306 1148 2358 1151
rect 2362 1148 2414 1151
rect 2418 1148 2462 1151
rect 2534 1151 2537 1158
rect 2490 1148 2537 1151
rect 2542 1151 2545 1158
rect 2542 1148 2630 1151
rect 2734 1151 2738 1152
rect 2706 1148 2738 1151
rect 1302 1142 1305 1148
rect 1958 1142 1961 1148
rect 2006 1142 2009 1148
rect 66 1138 110 1141
rect 214 1138 270 1141
rect 274 1138 286 1141
rect 362 1138 470 1141
rect 634 1138 934 1141
rect 938 1138 1022 1141
rect 1058 1138 1078 1141
rect 1082 1138 1166 1141
rect 1322 1138 1342 1141
rect 1362 1138 1366 1141
rect 1410 1138 1446 1141
rect 1498 1138 1630 1141
rect 1802 1138 1838 1141
rect 2074 1138 2158 1141
rect 2162 1138 2214 1141
rect 2246 1141 2249 1148
rect 2234 1138 2249 1141
rect 2254 1141 2257 1148
rect 2254 1138 2286 1141
rect 2306 1138 2310 1141
rect 2354 1138 2478 1141
rect 2506 1138 2510 1141
rect 2586 1138 2598 1141
rect 2626 1138 2662 1141
rect 174 1132 177 1138
rect 214 1132 217 1138
rect -26 1131 -22 1132
rect -26 1128 110 1131
rect 114 1128 118 1131
rect 266 1128 270 1131
rect 642 1128 870 1131
rect 882 1128 982 1131
rect 986 1128 993 1131
rect 1106 1128 1134 1131
rect 1262 1131 1265 1138
rect 1250 1128 1326 1131
rect 1338 1128 1366 1131
rect 1402 1128 1414 1131
rect 1474 1128 1502 1131
rect 1642 1128 1782 1131
rect 1922 1128 1934 1131
rect 2042 1128 2086 1131
rect 2090 1128 2182 1131
rect 2210 1128 2262 1131
rect 2266 1128 2390 1131
rect 2394 1128 2454 1131
rect 2458 1128 2502 1131
rect 2570 1128 2574 1131
rect 2734 1128 2738 1132
rect 138 1118 278 1121
rect 602 1118 630 1121
rect 818 1118 902 1121
rect 994 1118 998 1121
rect 1010 1118 1150 1121
rect 1550 1121 1553 1128
rect 1450 1118 1553 1121
rect 1658 1118 1742 1121
rect 1858 1118 1894 1121
rect 2050 1118 2094 1121
rect 2106 1118 2329 1121
rect 2426 1118 2470 1121
rect 370 1108 630 1111
rect 634 1108 638 1111
rect 834 1108 846 1111
rect 906 1108 1006 1111
rect 1490 1108 1734 1111
rect 1874 1108 1894 1111
rect 1978 1108 1998 1111
rect 2226 1108 2318 1111
rect 2326 1111 2329 1118
rect 2326 1108 2430 1111
rect 2466 1108 2534 1111
rect 2538 1108 2598 1111
rect 2602 1108 2614 1111
rect 2734 1108 2738 1112
rect 46 1102 49 1108
rect 1080 1103 1082 1107
rect 1086 1103 1089 1107
rect 1094 1103 1096 1107
rect 2104 1103 2106 1107
rect 2110 1103 2113 1107
rect 2118 1103 2120 1107
rect 2438 1102 2441 1108
rect 642 1098 662 1101
rect 666 1098 774 1101
rect 778 1098 870 1101
rect 1018 1098 1070 1101
rect 1386 1098 1430 1101
rect 1538 1098 1558 1101
rect 1562 1098 1710 1101
rect 1770 1098 1782 1101
rect 1842 1098 2006 1101
rect 2018 1098 2070 1101
rect 2126 1098 2342 1101
rect 2482 1098 2558 1101
rect 2562 1098 2737 1101
rect 30 1088 110 1091
rect 114 1088 182 1091
rect 414 1088 422 1091
rect 426 1088 526 1091
rect 530 1088 558 1091
rect 562 1088 598 1091
rect 602 1088 654 1091
rect 874 1088 1110 1091
rect 1114 1088 1206 1091
rect 1258 1088 1342 1091
rect 1346 1088 1470 1091
rect 1730 1088 1774 1091
rect 1794 1088 1846 1091
rect 1850 1088 1910 1091
rect 1914 1088 2006 1091
rect 2010 1088 2014 1091
rect 2126 1091 2129 1098
rect 2734 1092 2737 1098
rect 2090 1088 2129 1091
rect 2242 1088 2294 1091
rect 2490 1088 2526 1091
rect 2734 1088 2738 1092
rect 30 1082 33 1088
rect 42 1078 54 1081
rect 302 1081 305 1088
rect 302 1078 374 1081
rect 458 1078 486 1081
rect 522 1078 678 1081
rect 786 1078 838 1081
rect 954 1078 1006 1081
rect 1010 1078 1030 1081
rect 1058 1078 1193 1081
rect 1306 1078 1374 1081
rect 1434 1078 1478 1081
rect 1630 1081 1633 1088
rect 1586 1078 1633 1081
rect 1714 1078 1742 1081
rect 1930 1078 2014 1081
rect 2034 1078 2038 1081
rect 2042 1078 2054 1081
rect 2214 1081 2217 1088
rect 2170 1078 2217 1081
rect 2302 1081 2305 1088
rect 2302 1078 2318 1081
rect 2322 1078 2342 1081
rect 2610 1078 2638 1081
rect 2642 1078 2702 1081
rect 1190 1072 1193 1078
rect 1742 1072 1745 1078
rect 18 1068 46 1071
rect 90 1068 110 1071
rect 426 1068 454 1071
rect 542 1068 550 1071
rect 554 1068 582 1071
rect 834 1068 886 1071
rect 890 1068 902 1071
rect 962 1068 974 1071
rect 994 1068 1038 1071
rect 1042 1068 1070 1071
rect 1082 1068 1182 1071
rect 1242 1068 1246 1071
rect 1474 1068 1590 1071
rect 1634 1068 1662 1071
rect 1666 1068 1670 1071
rect 1706 1068 1718 1071
rect 1778 1068 1782 1071
rect 1826 1068 1830 1071
rect 2022 1071 2025 1078
rect 1914 1068 2046 1071
rect 2074 1068 2094 1071
rect 2158 1071 2161 1078
rect 2158 1068 2182 1071
rect 2250 1068 2270 1071
rect 2274 1068 2302 1071
rect 2618 1068 2662 1071
rect 2734 1068 2738 1072
rect 42 1058 46 1061
rect 54 1058 62 1061
rect 98 1058 102 1061
rect 218 1058 222 1061
rect 302 1061 305 1068
rect 302 1058 350 1061
rect 418 1058 478 1061
rect 742 1058 774 1061
rect 806 1058 1134 1061
rect 1162 1058 1222 1061
rect 1366 1061 1369 1068
rect 1298 1058 1369 1061
rect 2222 1062 2225 1068
rect 1394 1059 1438 1061
rect 1390 1058 1438 1059
rect 1506 1058 1622 1061
rect 1658 1058 1694 1061
rect 1698 1058 1702 1061
rect 1706 1058 1782 1061
rect 1826 1058 1846 1061
rect 1850 1058 1958 1061
rect 1962 1058 2062 1061
rect 2122 1058 2158 1061
rect 2162 1058 2185 1061
rect 2202 1058 2206 1061
rect 2314 1058 2318 1061
rect 2354 1058 2470 1061
rect 2562 1058 2646 1061
rect 54 1051 57 1058
rect 42 1048 57 1051
rect 158 1051 161 1058
rect 742 1052 745 1058
rect 806 1052 809 1058
rect 66 1048 161 1051
rect 202 1048 222 1051
rect 514 1048 534 1051
rect 826 1048 894 1051
rect 914 1048 958 1051
rect 978 1048 1006 1051
rect 1202 1048 1214 1051
rect 1418 1048 1446 1051
rect 1554 1048 1638 1051
rect 1682 1048 1710 1051
rect 1818 1048 1822 1051
rect 1826 1048 1833 1051
rect 1938 1048 1958 1051
rect 2010 1048 2174 1051
rect 2182 1051 2185 1058
rect 2334 1051 2337 1058
rect 2182 1048 2337 1051
rect 2478 1051 2481 1058
rect 2478 1048 2606 1051
rect 82 1038 126 1041
rect 138 1038 142 1041
rect 250 1038 334 1041
rect 338 1038 358 1041
rect 554 1038 614 1041
rect 618 1038 686 1041
rect 806 1041 809 1048
rect 690 1038 809 1041
rect 850 1038 862 1041
rect 1118 1041 1121 1048
rect 1082 1038 1121 1041
rect 1170 1038 1278 1041
rect 1750 1041 1753 1048
rect 1750 1038 1758 1041
rect 1882 1038 2070 1041
rect 2234 1038 2238 1041
rect 2242 1038 2398 1041
rect 2494 1038 2550 1041
rect 2634 1038 2670 1041
rect 2494 1032 2497 1038
rect 242 1028 318 1031
rect 1154 1028 1246 1031
rect 586 1018 942 1021
rect 1090 1018 1182 1021
rect 2482 1018 2582 1021
rect 2438 1012 2441 1018
rect 842 1008 1022 1011
rect 576 1003 578 1007
rect 582 1003 585 1007
rect 590 1003 592 1007
rect 1600 1003 1602 1007
rect 1606 1003 1609 1007
rect 1614 1003 1616 1007
rect 1898 998 2302 1001
rect 2306 998 2358 1001
rect 2362 998 2470 1001
rect 982 992 985 998
rect -26 988 -22 992
rect 642 988 750 991
rect 2010 988 2038 991
rect 2210 988 2494 991
rect 2498 988 2558 991
rect 666 978 774 981
rect 778 978 982 981
rect 986 978 1006 981
rect 1778 978 1822 981
rect 1826 978 1862 981
rect 1866 978 1918 981
rect 2242 978 2662 981
rect 2734 978 2738 982
rect 1038 972 1041 978
rect -26 971 -22 972
rect -26 968 6 971
rect 746 968 814 971
rect 818 968 846 971
rect 850 968 873 971
rect 1426 968 1454 971
rect 1458 968 1462 971
rect 1614 971 1617 978
rect 1614 968 1646 971
rect 1650 968 1750 971
rect 2058 968 2062 971
rect 2066 968 2110 971
rect 2394 968 2462 971
rect 2506 968 2646 971
rect 18 958 110 961
rect 234 958 286 961
rect 366 961 369 968
rect 870 962 873 968
rect 366 958 430 961
rect 474 958 502 961
rect 618 958 726 961
rect 1402 958 1406 961
rect 1594 958 1622 961
rect 1690 958 1694 961
rect 1854 961 1857 968
rect 1870 961 1873 968
rect 1854 958 1873 961
rect 2050 958 2094 961
rect 2098 958 2254 961
rect 2310 961 2313 968
rect 2282 958 2313 961
rect 2354 958 2358 961
rect 2410 958 2494 961
rect 2734 961 2738 962
rect 2562 958 2738 961
rect 950 952 953 958
rect -26 948 -22 952
rect 94 948 118 951
rect 122 948 142 951
rect 250 948 254 951
rect 410 948 486 951
rect 490 948 494 951
rect 514 948 654 951
rect 6 942 9 948
rect 94 942 97 948
rect 502 942 505 948
rect 730 948 750 951
rect 974 951 977 958
rect 974 948 1014 951
rect 1114 948 1177 951
rect 886 942 889 948
rect 1174 942 1177 948
rect 1206 948 1246 951
rect 1258 948 1406 951
rect 1410 948 1430 951
rect 1586 948 1638 951
rect 1690 948 1718 951
rect 1834 948 1902 951
rect 1906 948 2070 951
rect 2226 948 2398 951
rect 2402 948 2406 951
rect 2418 948 2534 951
rect 1206 942 1209 948
rect 2158 942 2161 948
rect 226 938 233 941
rect 250 938 262 941
rect 362 938 366 941
rect 530 938 534 941
rect 538 938 790 941
rect 1002 938 1062 941
rect 1098 938 1134 941
rect 1402 938 1441 941
rect 1530 938 1553 941
rect 1666 938 1694 941
rect 1778 938 1894 941
rect 2066 938 2094 941
rect 2338 938 2350 941
rect 2354 938 2374 941
rect 2394 938 2486 941
rect 2734 941 2738 942
rect 2626 938 2738 941
rect 230 932 233 938
rect -26 928 -22 932
rect 82 928 134 931
rect 470 931 473 938
rect 442 928 473 931
rect 482 928 550 931
rect 554 928 558 931
rect 602 928 606 931
rect 818 928 846 931
rect 934 931 937 938
rect 1382 932 1385 938
rect 1438 932 1441 938
rect 1550 932 1553 938
rect 2006 932 2009 938
rect 850 928 937 931
rect 970 928 982 931
rect 1426 928 1430 931
rect 1578 928 1622 931
rect 1626 928 1646 931
rect 1650 928 1726 931
rect 1730 928 1798 931
rect 1818 928 1862 931
rect 2026 928 2134 931
rect 2386 928 2414 931
rect 2546 928 2550 931
rect 350 922 353 928
rect 66 918 86 921
rect 386 918 422 921
rect 426 918 446 921
rect 450 918 462 921
rect 466 918 542 921
rect 1290 918 1318 921
rect 1690 918 1694 921
rect 2014 921 2017 928
rect 1954 918 2017 921
rect 2154 918 2182 921
rect 2366 921 2369 928
rect 2314 918 2369 921
rect 2386 918 2590 921
rect 2734 918 2738 922
rect -26 908 -22 912
rect 922 908 1054 911
rect 1802 908 1838 911
rect 1858 908 1886 911
rect 1970 908 2094 911
rect 2322 908 2374 911
rect 2514 908 2654 911
rect 1080 903 1082 907
rect 1086 903 1089 907
rect 1094 903 1096 907
rect 2104 903 2106 907
rect 2110 903 2113 907
rect 2118 903 2120 907
rect 578 898 766 901
rect 866 898 878 901
rect 1010 898 1030 901
rect 1210 898 1262 901
rect 1730 898 1758 901
rect 1874 898 1934 901
rect 1938 898 2006 901
rect 2154 898 2294 901
rect 2298 898 2430 901
rect 2594 898 2686 901
rect 302 892 305 898
rect 138 888 190 891
rect 482 888 534 891
rect 762 888 814 891
rect 886 891 889 898
rect 826 888 889 891
rect 938 888 1078 891
rect 1082 888 1142 891
rect 1466 888 1590 891
rect 1594 888 1598 891
rect 1658 888 1825 891
rect 270 882 273 888
rect 574 881 577 888
rect 522 878 577 881
rect 682 878 710 881
rect 714 878 750 881
rect 754 878 846 881
rect 850 878 966 881
rect 970 878 1046 881
rect 1302 881 1305 888
rect 1822 882 1825 888
rect 1882 888 1886 891
rect 1906 888 1910 891
rect 1982 888 2262 891
rect 2266 888 2430 891
rect 2458 888 2510 891
rect 2514 888 2518 891
rect 2530 888 2606 891
rect 2734 891 2738 892
rect 2642 888 2738 891
rect 1274 878 1305 881
rect 1458 878 1558 881
rect 1594 878 1622 881
rect 1650 878 1670 881
rect 1722 878 1814 881
rect 1830 881 1833 888
rect 1982 882 1985 888
rect 1830 878 1958 881
rect 1962 878 1974 881
rect 1994 878 2062 881
rect 2066 878 2150 881
rect 2202 878 2249 881
rect 2258 878 2270 881
rect 2370 878 2462 881
rect 2466 878 2678 881
rect 10 868 30 871
rect 214 871 217 878
rect 2246 872 2249 878
rect 214 868 326 871
rect 498 868 558 871
rect 562 868 574 871
rect 906 868 990 871
rect 1026 868 1086 871
rect 1618 868 1646 871
rect 1706 868 1846 871
rect 1858 868 1918 871
rect 1946 868 2022 871
rect 2066 868 2070 871
rect 2218 868 2230 871
rect 2258 868 2278 871
rect 2318 871 2321 878
rect 2318 868 2334 871
rect 2554 868 2558 871
rect 2582 868 2622 871
rect 2734 868 2738 872
rect 186 858 262 861
rect 446 861 449 868
rect 446 858 598 861
rect 734 861 737 868
rect 734 858 766 861
rect 1014 858 1022 861
rect 1026 858 1118 861
rect 1126 861 1129 868
rect 1126 858 1150 861
rect 1270 861 1273 868
rect 1270 858 1302 861
rect 1526 861 1529 868
rect 1702 862 1705 868
rect 2582 862 2585 868
rect 1526 858 1606 861
rect 1818 858 1950 861
rect 1954 858 1958 861
rect 2082 858 2126 861
rect 2186 858 2222 861
rect 2242 858 2342 861
rect 2394 858 2446 861
rect 2538 858 2566 861
rect 18 848 46 851
rect 114 848 158 851
rect 162 848 270 851
rect 274 848 350 851
rect 354 848 358 851
rect 546 848 582 851
rect 634 848 750 851
rect 1010 848 1166 851
rect 1170 848 1238 851
rect 1594 848 1798 851
rect 1850 848 1958 851
rect 1998 848 2049 851
rect 1998 842 2001 848
rect 2046 842 2049 848
rect 2082 848 2086 851
rect 2202 848 2318 851
rect 2454 848 2518 851
rect 2570 848 2574 851
rect 2054 842 2057 848
rect 2454 842 2457 848
rect 498 838 502 841
rect 658 838 726 841
rect 1418 838 1526 841
rect 1786 838 1942 841
rect 1962 838 1990 841
rect 2346 838 2350 841
rect 654 832 657 838
rect 482 828 566 831
rect 1154 828 1174 831
rect 1178 828 1374 831
rect 2042 828 2198 831
rect 2546 828 2622 831
rect -26 818 -22 822
rect 34 818 62 821
rect 66 818 110 821
rect 626 818 742 821
rect 1322 818 1358 821
rect 1362 818 1406 821
rect 1954 818 2182 821
rect 1890 808 1990 811
rect 1994 808 2086 811
rect 576 803 578 807
rect 582 803 585 807
rect 590 803 592 807
rect 1600 803 1602 807
rect 1606 803 1609 807
rect 1614 803 1616 807
rect 986 798 1014 801
rect 1802 798 2046 801
rect 2490 798 2566 801
rect 466 788 526 791
rect 562 788 574 791
rect 2426 788 2526 791
rect -26 778 -22 782
rect 82 778 86 781
rect 178 778 182 781
rect 2450 778 2574 781
rect 2686 781 2689 788
rect 2602 778 2689 781
rect 102 771 105 778
rect 302 772 305 778
rect 58 768 105 771
rect 130 768 174 771
rect 562 768 606 771
rect 610 768 726 771
rect 762 768 798 771
rect 802 768 950 771
rect 1818 768 1830 771
rect 1858 768 1910 771
rect 2058 768 2222 771
rect 2242 768 2294 771
rect 2482 768 2566 771
rect 2570 768 2606 771
rect -26 761 -22 762
rect -26 758 6 761
rect 10 758 94 761
rect 98 758 134 761
rect 170 758 206 761
rect 234 758 238 761
rect 242 758 254 761
rect 270 761 273 768
rect 310 761 313 768
rect 270 758 313 761
rect 446 761 449 768
rect 446 758 510 761
rect 658 758 718 761
rect 1594 758 1614 761
rect 1854 761 1857 768
rect 1674 758 1857 761
rect 1942 762 1945 768
rect 2014 761 2017 768
rect 2014 758 2078 761
rect 2098 758 2286 761
rect 2290 758 2382 761
rect 2386 758 2406 761
rect 2410 758 2438 761
rect 2442 758 2550 761
rect 2658 758 2670 761
rect 38 748 46 751
rect 50 748 54 751
rect 98 748 102 751
rect 114 748 158 751
rect 162 748 182 751
rect 282 748 286 751
rect 458 748 470 751
rect 62 741 65 748
rect 270 742 273 748
rect 494 742 497 748
rect 658 748 694 751
rect 730 748 766 751
rect 786 748 894 751
rect 898 748 950 751
rect 1086 751 1089 758
rect 2590 752 2593 758
rect 978 748 1089 751
rect 1114 748 1182 751
rect 1202 748 1217 751
rect 1214 742 1217 748
rect 1246 748 1366 751
rect 1562 748 1606 751
rect 1610 748 1622 751
rect 1626 748 1638 751
rect 1690 748 1814 751
rect 1850 748 1918 751
rect 1962 748 1998 751
rect 2058 748 2134 751
rect 1246 742 1249 748
rect 26 738 65 741
rect 178 738 246 741
rect 426 738 446 741
rect 546 738 702 741
rect 722 738 902 741
rect 906 738 918 741
rect 954 738 1006 741
rect 1366 741 1369 748
rect 1446 741 1449 748
rect 1366 738 1449 741
rect 1474 738 1510 741
rect 1514 738 1574 741
rect 1650 738 1734 741
rect 1850 738 1862 741
rect 1890 738 1894 741
rect 1934 741 1937 748
rect 2266 748 2294 751
rect 2330 748 2342 751
rect 2370 748 2390 751
rect 2394 748 2401 751
rect 2642 748 2662 751
rect 2734 751 2738 752
rect 2666 748 2738 751
rect 1934 738 1958 741
rect 2026 738 2062 741
rect 2074 738 2078 741
rect 2098 738 2113 741
rect 2178 738 2230 741
rect 2274 738 2302 741
rect 2378 738 2398 741
rect 2402 738 2406 741
rect 2522 738 2638 741
rect 1022 732 1025 738
rect 1038 732 1041 738
rect 146 728 222 731
rect 226 728 246 731
rect 266 728 278 731
rect 466 728 478 731
rect 602 728 694 731
rect 746 728 838 731
rect 962 728 966 731
rect 1050 728 1438 731
rect 1442 728 1662 731
rect 1782 731 1785 738
rect 2110 732 2113 738
rect 1714 728 1785 731
rect 1794 728 1798 731
rect 2034 728 2046 731
rect 2162 728 2278 731
rect 2282 728 2430 731
rect 2562 728 2590 731
rect 2634 728 2638 731
rect -26 718 -22 722
rect 138 718 142 721
rect 226 718 230 721
rect 242 718 318 721
rect 338 718 382 721
rect 498 718 518 721
rect 706 718 758 721
rect 890 718 942 721
rect 946 718 1070 721
rect 1074 718 1158 721
rect 1298 718 1390 721
rect 1754 718 1758 721
rect 1870 721 1873 728
rect 1778 718 1873 721
rect 2026 718 2094 721
rect 2202 718 2206 721
rect 2218 718 2294 721
rect 2306 718 2390 721
rect 2410 718 2430 721
rect 2442 718 2486 721
rect 2674 718 2686 721
rect 174 712 177 718
rect 790 712 793 718
rect 226 708 230 711
rect 378 708 430 711
rect 562 708 622 711
rect 626 708 678 711
rect 682 708 734 711
rect 842 708 982 711
rect 1210 708 1254 711
rect 1354 708 1438 711
rect 1626 708 1694 711
rect 1826 708 1958 711
rect 2042 708 2054 711
rect 2242 708 2270 711
rect 2290 708 2342 711
rect 2658 708 2678 711
rect 310 702 313 708
rect 1080 703 1082 707
rect 1086 703 1089 707
rect 1094 703 1096 707
rect 2104 703 2106 707
rect 2110 703 2113 707
rect 2118 703 2120 707
rect 570 698 718 701
rect 898 698 990 701
rect 1178 698 1230 701
rect 1410 698 1566 701
rect 1914 698 2022 701
rect 2066 698 2097 701
rect 2202 698 2374 701
rect 2378 698 2438 701
rect 258 688 270 691
rect 274 688 294 691
rect 434 688 478 691
rect 754 688 758 691
rect 762 688 846 691
rect 850 688 966 691
rect 1082 688 1350 691
rect 1354 688 1382 691
rect 1402 688 1446 691
rect 1450 688 1510 691
rect 1946 688 2046 691
rect 2058 688 2086 691
rect 2094 691 2097 698
rect 2094 688 2246 691
rect 2274 688 2326 691
rect 2570 688 2737 691
rect 182 682 185 688
rect 246 681 249 688
rect 2734 682 2737 688
rect 234 678 249 681
rect 394 678 414 681
rect 418 678 454 681
rect 458 678 550 681
rect 554 678 934 681
rect 938 678 1254 681
rect 1258 678 1278 681
rect 1354 678 1654 681
rect 1738 678 1766 681
rect 2010 678 2198 681
rect 2202 678 2422 681
rect 2426 678 2494 681
rect 2554 678 2574 681
rect 2734 678 2738 682
rect -26 671 -22 672
rect -26 668 6 671
rect 10 668 70 671
rect 90 668 94 671
rect 154 668 182 671
rect 286 671 289 678
rect 286 668 310 671
rect 366 671 369 678
rect 346 668 369 671
rect 426 668 478 671
rect 538 668 598 671
rect 618 668 662 671
rect 698 668 798 671
rect 802 668 854 671
rect 858 668 1014 671
rect 1122 668 1190 671
rect 1242 668 1270 671
rect 1274 668 1334 671
rect 1338 668 1406 671
rect 1410 668 1446 671
rect 1530 668 1550 671
rect 1762 668 1790 671
rect 1794 668 1838 671
rect 1866 668 1902 671
rect 1922 668 1934 671
rect 1938 668 2142 671
rect 2154 668 2230 671
rect 2338 668 2358 671
rect 2386 668 2454 671
rect 2462 668 2478 671
rect 2574 671 2577 678
rect 2574 668 2630 671
rect 222 662 225 668
rect 50 658 86 661
rect 202 658 206 661
rect 258 658 286 661
rect 362 658 382 661
rect 386 658 510 661
rect 514 658 606 661
rect 610 658 686 661
rect 690 658 790 661
rect 794 658 822 661
rect 890 658 902 661
rect 978 658 982 661
rect 1002 658 1054 661
rect 1058 658 1126 661
rect 1182 658 1206 661
rect 1274 658 1398 661
rect 1402 658 1454 661
rect 1514 658 1561 661
rect 1810 658 1862 661
rect 1866 658 1886 661
rect 1890 658 1918 661
rect 1994 658 2118 661
rect 2138 658 2158 661
rect 2162 658 2198 661
rect 2378 658 2382 661
rect 2462 661 2465 668
rect 2418 658 2465 661
rect 2482 658 2486 661
rect 2510 661 2513 668
rect 2662 662 2665 668
rect 2510 658 2662 661
rect -26 648 -22 652
rect 38 651 41 658
rect 1182 652 1185 658
rect 1558 652 1561 658
rect 2286 652 2289 658
rect 2294 652 2297 658
rect 26 648 41 651
rect 82 648 94 651
rect 98 648 158 651
rect 202 648 262 651
rect 362 648 422 651
rect 450 648 454 651
rect 650 648 654 651
rect 658 648 894 651
rect 1050 648 1078 651
rect 2370 648 2502 651
rect 2506 648 2526 651
rect 318 642 321 648
rect 122 638 190 641
rect 402 638 438 641
rect 602 638 638 641
rect 714 638 718 641
rect 826 638 886 641
rect 926 641 929 648
rect 914 638 929 641
rect 1142 641 1145 648
rect 1142 638 1238 641
rect 1242 638 1270 641
rect 1478 641 1481 648
rect 1298 638 1510 641
rect 2122 638 2150 641
rect 2362 638 2518 641
rect 86 632 89 638
rect 710 628 718 631
rect 722 628 750 631
rect 786 628 846 631
rect 1054 631 1057 638
rect 1054 628 1110 631
rect 1114 628 1174 631
rect 2446 628 2486 631
rect 2446 622 2449 628
rect 490 618 990 621
rect 1170 618 1302 621
rect 1354 618 1422 621
rect 1426 618 1590 621
rect 2298 618 2310 621
rect 2314 618 2358 621
rect 2734 618 2738 622
rect 634 608 718 611
rect 954 608 1278 611
rect 576 603 578 607
rect 582 603 585 607
rect 590 603 592 607
rect 1600 603 1602 607
rect 1606 603 1609 607
rect 1614 603 1616 607
rect 986 598 1318 601
rect 1634 598 1814 601
rect 338 588 438 591
rect 442 588 494 591
rect 498 588 542 591
rect 658 588 806 591
rect 810 588 902 591
rect 1106 588 1222 591
rect 1426 588 1438 591
rect 1594 588 1654 591
rect 1658 588 1678 591
rect 1926 591 1929 598
rect 1926 588 1942 591
rect 2354 588 2398 591
rect 2734 591 2738 592
rect 2626 588 2738 591
rect 298 578 1046 581
rect 1090 578 1126 581
rect 1234 578 1454 581
rect 666 568 694 571
rect 1034 568 1062 571
rect 1210 568 1238 571
rect 1282 568 1326 571
rect 1450 568 1478 571
rect 1762 568 1806 571
rect 1834 568 1910 571
rect 2410 568 2430 571
rect 2734 568 2738 572
rect 38 561 41 568
rect 38 558 110 561
rect 302 561 305 568
rect 210 558 305 561
rect 526 561 529 568
rect 498 558 529 561
rect 994 558 1030 561
rect 1234 558 1302 561
rect 1306 558 1462 561
rect 1466 558 1486 561
rect 1490 558 1542 561
rect 1730 558 1790 561
rect 2614 561 2617 568
rect 2602 558 2617 561
rect 134 551 137 558
rect 114 548 137 551
rect 170 548 174 551
rect 178 548 222 551
rect 386 548 398 551
rect 326 542 329 548
rect 370 538 374 541
rect 510 541 513 548
rect 634 548 678 551
rect 690 548 734 551
rect 738 548 745 551
rect 798 551 801 558
rect 778 548 801 551
rect 1010 548 1022 551
rect 510 538 534 541
rect 538 538 622 541
rect 674 538 790 541
rect 910 541 913 548
rect 1154 548 1201 551
rect 1198 542 1201 548
rect 1214 548 1238 551
rect 1258 548 1286 551
rect 1290 548 1302 551
rect 1318 548 1326 551
rect 1346 548 1382 551
rect 1214 542 1217 548
rect 910 538 1126 541
rect 1274 538 1278 541
rect 1318 541 1321 548
rect 1406 548 1438 551
rect 1442 548 1622 551
rect 1674 548 1774 551
rect 1778 548 1782 551
rect 1862 551 1865 558
rect 1818 548 1865 551
rect 2050 548 2062 551
rect 2186 548 2286 551
rect 2290 548 2310 551
rect 2338 548 2606 551
rect 2618 548 2622 551
rect 2694 551 2697 558
rect 2734 551 2738 552
rect 2626 548 2738 551
rect 1406 542 1409 548
rect 1282 538 1321 541
rect 1330 538 1334 541
rect 1666 538 1702 541
rect 1738 538 1742 541
rect 1810 538 1814 541
rect 2046 538 2054 541
rect 2102 541 2105 548
rect 2058 538 2105 541
rect 2170 538 2446 541
rect 2450 538 2574 541
rect 2602 538 2662 541
rect -26 528 -22 532
rect 10 528 62 531
rect 150 528 182 531
rect 354 528 382 531
rect 818 528 822 531
rect 826 528 937 531
rect 1250 528 1278 531
rect 1282 528 1294 531
rect 1322 528 1334 531
rect 1570 528 1582 531
rect 1762 528 1766 531
rect 2054 528 2118 531
rect 2394 528 2441 531
rect 2582 531 2585 538
rect 2514 528 2585 531
rect 2610 528 2670 531
rect 150 522 153 528
rect 210 518 254 521
rect 390 521 393 528
rect 934 522 937 528
rect 2054 522 2057 528
rect 2438 522 2441 528
rect 322 518 393 521
rect 618 518 694 521
rect 1738 518 1766 521
rect 1770 518 1806 521
rect 2194 518 2302 521
rect 2522 518 2550 521
rect -26 508 -22 512
rect 578 508 694 511
rect 698 508 718 511
rect 898 508 942 511
rect 1706 508 1878 511
rect 1898 508 1958 511
rect 1962 508 1982 511
rect 2002 508 2070 511
rect 2274 508 2294 511
rect 2554 508 2598 511
rect 1080 503 1082 507
rect 1086 503 1089 507
rect 1094 503 1096 507
rect 2104 503 2106 507
rect 2110 503 2113 507
rect 2118 503 2120 507
rect -26 498 246 501
rect 410 498 422 501
rect 666 498 718 501
rect 794 498 921 501
rect 1578 498 1598 501
rect 2658 498 2678 501
rect 2734 498 2738 502
rect -26 492 -23 498
rect 918 492 921 498
rect 2278 492 2281 498
rect -26 488 -22 492
rect 34 488 86 491
rect 442 488 470 491
rect 474 488 542 491
rect 578 488 638 491
rect 826 488 878 491
rect 922 488 966 491
rect 970 488 1014 491
rect 1218 488 1222 491
rect 2282 488 2334 491
rect 2510 488 2550 491
rect 2562 488 2638 491
rect 298 478 302 481
rect 370 478 374 481
rect 574 481 577 488
rect 562 478 577 481
rect 698 478 702 481
rect 834 478 894 481
rect 906 478 926 481
rect 962 478 990 481
rect 994 478 1086 481
rect 1090 478 1190 481
rect 1242 478 1270 481
rect 1758 481 1761 488
rect 2510 482 2513 488
rect 1722 478 1870 481
rect 1874 478 1942 481
rect 1946 478 2062 481
rect 2458 478 2502 481
rect 2538 478 2566 481
rect 2570 478 2694 481
rect 142 472 145 478
rect -26 468 -22 472
rect 74 468 142 471
rect 294 471 297 478
rect 282 468 297 471
rect 634 468 654 471
rect 754 468 782 471
rect 786 468 910 471
rect 914 468 1030 471
rect 1034 468 1054 471
rect 1282 468 1302 471
rect 1410 468 1478 471
rect 1482 468 1502 471
rect 1994 468 2014 471
rect 2434 468 2534 471
rect 2734 471 2738 472
rect 2706 468 2738 471
rect 74 458 102 461
rect 178 458 198 461
rect 242 458 246 461
rect 250 458 286 461
rect 290 458 318 461
rect 494 461 497 468
rect 526 461 529 468
rect 494 458 529 461
rect 634 458 646 461
rect 650 458 694 461
rect 698 458 726 461
rect 754 458 825 461
rect 842 458 918 461
rect 938 458 1110 461
rect 1198 461 1201 468
rect 1198 458 1262 461
rect 1290 458 1310 461
rect 1334 458 1441 461
rect 1722 459 1742 461
rect 1718 458 1742 459
rect 2014 461 2017 468
rect 1894 458 1929 461
rect 2014 458 2030 461
rect 2126 461 2129 468
rect 2486 462 2489 468
rect 2098 458 2129 461
rect 2154 458 2254 461
rect 2258 458 2425 461
rect 2514 458 2590 461
rect 822 452 825 458
rect 1334 452 1337 458
rect 1438 452 1441 458
rect 1894 452 1897 458
rect 1926 452 1929 458
rect 2326 452 2329 458
rect 2422 452 2425 458
rect 98 448 150 451
rect 698 448 758 451
rect 874 448 958 451
rect 1058 448 1086 451
rect 1258 448 1278 451
rect 1298 448 1302 451
rect 2362 448 2390 451
rect 2426 448 2502 451
rect 2538 448 2558 451
rect 2734 448 2738 452
rect 318 442 321 448
rect 1110 442 1113 448
rect 1350 441 1353 448
rect 2526 442 2529 448
rect 1218 438 1353 441
rect 1538 438 1742 441
rect 642 428 670 431
rect 674 428 830 431
rect 1058 428 1230 431
rect 1234 428 1246 431
rect 2506 428 2614 431
rect 562 418 1574 421
rect 1578 418 1630 421
rect 1634 418 1758 421
rect 2594 418 2598 421
rect 576 403 578 407
rect 582 403 585 407
rect 590 403 592 407
rect 822 402 825 408
rect 1600 403 1602 407
rect 1606 403 1609 407
rect 1614 403 1616 407
rect 2562 398 2614 401
rect 570 388 774 391
rect 1050 388 1062 391
rect 1066 388 1150 391
rect 1154 388 1238 391
rect 2026 388 2174 391
rect 2322 388 2334 391
rect 834 378 862 381
rect 866 378 1110 381
rect 1194 378 1198 381
rect 2546 378 2590 381
rect 34 368 278 371
rect 786 368 982 371
rect 1390 368 1454 371
rect 1650 368 1974 371
rect 2338 368 2398 371
rect 1390 362 1393 368
rect -26 361 -22 362
rect -26 358 134 361
rect 202 358 270 361
rect 306 358 374 361
rect 498 358 558 361
rect 626 358 662 361
rect 1066 358 1206 361
rect 1234 358 1246 361
rect 1250 358 1294 361
rect 1410 358 1574 361
rect 1578 358 1734 361
rect 1882 358 1894 361
rect 1898 358 1918 361
rect 2050 358 2062 361
rect 2298 358 2462 361
rect 2466 358 2542 361
rect 2546 358 2582 361
rect 2618 358 2678 361
rect 130 348 150 351
rect 162 348 182 351
rect 274 348 326 351
rect 458 348 470 351
rect 506 348 638 351
rect 642 348 702 351
rect 706 348 766 351
rect 854 351 857 358
rect 826 348 857 351
rect 954 348 990 351
rect 1018 348 1190 351
rect 1214 348 1222 351
rect 1226 348 1297 351
rect 1398 351 1401 358
rect 1814 352 1817 358
rect 1386 348 1401 351
rect 1562 348 1590 351
rect 1594 348 1641 351
rect 6 341 9 348
rect 310 342 313 348
rect 1294 342 1297 348
rect 1638 342 1641 348
rect 1670 348 1718 351
rect 1746 348 1774 351
rect 1910 348 2038 351
rect 2042 348 2062 351
rect 2118 351 2121 358
rect 2090 348 2121 351
rect 2346 348 2462 351
rect 2466 348 2470 351
rect 2474 348 2622 351
rect 1670 342 1673 348
rect 6 338 62 341
rect 146 338 150 341
rect 170 338 198 341
rect 242 338 246 341
rect 418 338 446 341
rect 1194 338 1214 341
rect 1242 338 1246 341
rect 1346 338 1406 341
rect 1410 338 1518 341
rect 1522 338 1542 341
rect 1798 341 1801 348
rect 1690 338 1801 341
rect 1910 341 1913 348
rect 2246 342 2249 348
rect 1890 338 1918 341
rect 2010 338 2105 341
rect 990 332 993 338
rect 2102 332 2105 338
rect 2190 338 2206 341
rect 2322 338 2361 341
rect 2190 332 2193 338
rect 2358 332 2361 338
rect 2466 338 2558 341
rect 2610 338 2630 341
rect 2422 332 2425 338
rect 186 328 241 331
rect 938 328 974 331
rect 1042 328 1166 331
rect 1226 328 1366 331
rect 1394 328 1414 331
rect 1418 328 1422 331
rect 1770 328 1774 331
rect 1922 328 1934 331
rect 2234 328 2310 331
rect 2442 328 2446 331
rect 238 322 241 328
rect 146 318 214 321
rect 730 318 766 321
rect 770 318 950 321
rect 994 318 1022 321
rect 1042 318 1102 321
rect 1282 318 1566 321
rect 1618 318 1702 321
rect 2058 318 2246 321
rect 2258 318 2422 321
rect 2602 318 2638 321
rect 2642 318 2654 321
rect 138 308 174 311
rect 178 308 286 311
rect 290 308 406 311
rect 914 308 982 311
rect 986 308 1054 311
rect 1258 308 1318 311
rect 1322 308 1358 311
rect 1362 308 1526 311
rect 1858 308 1862 311
rect 2162 308 2198 311
rect 2210 308 2366 311
rect 2378 308 2566 311
rect 1080 303 1082 307
rect 1086 303 1089 307
rect 1094 303 1096 307
rect 2104 303 2106 307
rect 2110 303 2113 307
rect 2118 303 2120 307
rect -26 298 -22 302
rect 90 298 206 301
rect 1306 298 1326 301
rect 1330 298 1454 301
rect 1634 298 1662 301
rect 1666 298 1750 301
rect 1754 298 1782 301
rect 2410 298 2430 301
rect 2522 298 2590 301
rect 2382 292 2385 298
rect 210 288 222 291
rect 682 288 726 291
rect 842 288 846 291
rect 1018 288 1174 291
rect 1218 288 1222 291
rect 1266 288 1294 291
rect 1314 288 1334 291
rect 1538 288 1681 291
rect 2050 288 2334 291
rect 2394 288 2446 291
rect 2546 288 2574 291
rect -26 281 -22 282
rect -26 278 6 281
rect 150 281 153 288
rect 1678 282 1681 288
rect 150 278 182 281
rect 218 278 222 281
rect 666 278 686 281
rect 690 278 926 281
rect 978 278 1046 281
rect 1050 278 1078 281
rect 1090 278 1110 281
rect 1194 278 1230 281
rect 1234 278 1390 281
rect 1514 278 1574 281
rect 1578 278 1654 281
rect 1826 278 1942 281
rect 2082 278 2102 281
rect 2286 278 2294 281
rect 2298 278 2310 281
rect 2330 278 2374 281
rect 2490 278 2542 281
rect 2578 278 2662 281
rect 42 268 70 271
rect 98 268 166 271
rect 258 268 294 271
rect 370 268 438 271
rect 658 268 998 271
rect 1058 268 1110 271
rect 1322 268 1350 271
rect 1354 268 1406 271
rect 1494 271 1497 278
rect 1494 268 1526 271
rect 1530 268 1537 271
rect 1722 268 1902 271
rect 1930 268 2014 271
rect 2174 271 2177 278
rect 2090 268 2177 271
rect 2202 268 2270 271
rect 2274 268 2294 271
rect 2486 271 2489 278
rect 2434 268 2489 271
rect 2554 268 2617 271
rect 66 258 110 261
rect 114 258 118 261
rect 282 258 310 261
rect 442 258 457 261
rect 474 258 518 261
rect 606 261 609 268
rect 2374 262 2377 268
rect 2614 262 2617 268
rect 2734 268 2738 272
rect 2638 262 2641 268
rect 546 258 609 261
rect 706 258 710 261
rect 714 258 950 261
rect 954 258 1070 261
rect 1074 258 1254 261
rect 1282 258 1286 261
rect 1370 258 1518 261
rect 1534 258 1569 261
rect 1642 258 1822 261
rect 2010 258 2214 261
rect 2218 258 2262 261
rect 2266 258 2278 261
rect 2442 258 2462 261
rect 2486 258 2521 261
rect 454 252 457 258
rect 1534 252 1537 258
rect 1566 252 1569 258
rect 2486 252 2489 258
rect 2518 252 2521 258
rect 178 248 198 251
rect 250 248 294 251
rect 718 248 758 251
rect 786 248 862 251
rect 898 248 937 251
rect 946 248 1014 251
rect 1066 248 1102 251
rect 1118 248 1150 251
rect 1186 248 1302 251
rect 1362 248 1366 251
rect 1382 248 1470 251
rect 1674 248 1814 251
rect 2098 248 2118 251
rect 2366 248 2374 251
rect 2378 248 2382 251
rect 2734 248 2738 252
rect 718 242 721 248
rect 934 242 937 248
rect 1118 242 1121 248
rect 1382 242 1385 248
rect 562 238 662 241
rect 1794 238 2070 241
rect 2146 238 2166 241
rect 2170 238 2422 241
rect 2426 238 2430 241
rect 2442 238 2446 241
rect 362 228 390 231
rect 394 228 486 231
rect 490 228 638 231
rect 642 228 782 231
rect 922 228 982 231
rect 2114 228 2342 231
rect 466 218 510 221
rect 514 218 686 221
rect 858 218 974 221
rect 978 218 1006 221
rect 1194 218 1430 221
rect 1434 218 1614 221
rect 2562 218 2574 221
rect 898 208 990 211
rect 576 203 578 207
rect 582 203 585 207
rect 590 203 592 207
rect 1600 203 1602 207
rect 1606 203 1609 207
rect 1614 203 1616 207
rect 2074 188 2246 191
rect 2250 188 2382 191
rect 2386 188 2478 191
rect 2482 188 2502 191
rect 2154 178 2182 181
rect 678 172 681 178
rect -26 168 -22 172
rect 538 168 630 171
rect 842 168 1478 171
rect 2058 168 2070 171
rect 2098 168 2230 171
rect 2282 168 2310 171
rect 2314 168 2350 171
rect 2510 171 2513 178
rect 2410 168 2513 171
rect 594 158 641 161
rect 694 161 697 168
rect 658 158 697 161
rect 722 158 822 161
rect 874 158 910 161
rect 1106 158 1134 161
rect 1314 158 1374 161
rect 1698 158 1766 161
rect 1882 158 1982 161
rect 2010 158 2518 161
rect 2526 158 2638 161
rect -26 148 -22 152
rect 34 148 94 151
rect 162 148 230 151
rect 398 151 401 158
rect 638 152 641 158
rect 346 148 401 151
rect 442 148 470 151
rect 682 148 702 151
rect 722 148 849 151
rect 922 148 926 151
rect 946 148 950 151
rect 1122 148 1158 151
rect 1182 151 1185 158
rect 1574 152 1577 158
rect 2526 152 2529 158
rect 1182 148 1222 151
rect 1234 148 1382 151
rect 1482 148 1550 151
rect 1738 148 1830 151
rect 1890 148 1926 151
rect 2002 148 2062 151
rect 2082 148 2110 151
rect 2186 148 2201 151
rect 2234 148 2238 151
rect 2338 148 2358 151
rect 2402 148 2462 151
rect 2466 148 2470 151
rect 262 141 265 148
rect 310 141 313 148
rect 846 142 849 148
rect 1230 142 1233 148
rect 2198 142 2201 148
rect 262 138 313 141
rect 506 138 606 141
rect 634 138 654 141
rect 658 138 670 141
rect 690 138 718 141
rect 722 138 782 141
rect 890 138 894 141
rect 1002 138 1022 141
rect 1026 138 1110 141
rect 1162 138 1230 141
rect 1378 138 1470 141
rect 1482 138 1486 141
rect 1490 138 1630 141
rect 1802 138 1846 141
rect 1954 138 1966 141
rect 2042 138 2054 141
rect 2058 138 2142 141
rect 2274 138 2286 141
rect 2290 138 2414 141
rect 2418 138 2462 141
rect 2486 141 2489 148
rect 2590 142 2593 148
rect 2466 138 2489 141
rect 678 132 681 138
rect 2526 132 2529 138
rect 2566 132 2569 138
rect -26 128 -22 132
rect 498 128 566 131
rect 682 128 806 131
rect 810 128 846 131
rect 906 128 926 131
rect 946 128 950 131
rect 986 128 1006 131
rect 1010 128 1014 131
rect 1026 128 1054 131
rect 1138 128 1190 131
rect 1202 128 1230 131
rect 1250 128 1366 131
rect 1554 128 1622 131
rect 1626 128 1694 131
rect 2074 128 2102 131
rect 2106 128 2166 131
rect 2250 128 2294 131
rect 2298 128 2374 131
rect 2378 128 2422 131
rect 2426 128 2486 131
rect 18 118 22 121
rect 46 121 49 128
rect 26 118 49 121
rect 402 118 414 121
rect 418 118 470 121
rect 506 118 526 121
rect 754 118 886 121
rect 890 118 1105 121
rect 1114 118 1174 121
rect 1210 118 1238 121
rect 1250 118 1326 121
rect 1346 118 1414 121
rect 1950 121 1953 128
rect 1950 118 2134 121
rect 2554 118 2678 121
rect 2682 118 2686 121
rect 874 108 982 111
rect 1050 108 1054 111
rect 1102 111 1105 118
rect 1102 108 1438 111
rect 1882 108 1902 111
rect 2162 108 2342 111
rect 2346 108 2550 111
rect 2634 108 2694 111
rect 1080 103 1082 107
rect 1086 103 1089 107
rect 1094 103 1096 107
rect 2104 103 2106 107
rect 2110 103 2113 107
rect 2118 103 2120 107
rect -26 98 -22 102
rect 474 98 582 101
rect 586 98 646 101
rect 866 98 894 101
rect 1106 98 1126 101
rect 1170 98 1246 101
rect 1250 98 1401 101
rect 1514 98 1534 101
rect 1538 98 1590 101
rect 1594 98 1646 101
rect 1650 98 1758 101
rect 1818 98 1910 101
rect 1914 98 2054 101
rect 2218 98 2321 101
rect 2338 98 2414 101
rect 2538 98 2574 101
rect 1398 92 1401 98
rect 58 88 86 91
rect 130 88 158 91
rect 162 88 262 91
rect 266 88 278 91
rect 282 88 438 91
rect 562 88 638 91
rect 674 88 734 91
rect 746 88 910 91
rect 914 88 942 91
rect 1058 88 1062 91
rect 1066 88 1110 91
rect 1162 88 1254 91
rect 1258 88 1302 91
rect 1306 88 1342 91
rect 1402 88 1542 91
rect 1706 88 1718 91
rect 1898 88 2182 91
rect 2186 88 2270 91
rect 2318 91 2321 98
rect 2318 88 2414 91
rect 2578 88 2622 91
rect 2686 82 2689 88
rect 250 78 342 81
rect 410 78 502 81
rect 610 78 750 81
rect 802 78 838 81
rect 986 78 1006 81
rect 1034 78 1038 81
rect 1042 78 1166 81
rect 1178 78 1214 81
rect 1226 78 1230 81
rect 1314 78 1318 81
rect 1354 78 1366 81
rect 1370 78 1526 81
rect 1850 78 1942 81
rect 1986 78 2222 81
rect 2242 78 2294 81
rect 2514 78 2526 81
rect 2570 78 2590 81
rect 2734 78 2738 82
rect -26 71 -22 72
rect 6 71 9 78
rect -26 68 9 71
rect 530 68 694 71
rect 698 68 702 71
rect 738 68 774 71
rect 786 68 806 71
rect 826 68 854 71
rect 918 71 921 78
rect 898 68 921 71
rect 938 68 966 71
rect 986 68 990 71
rect 1002 68 1022 71
rect 1042 68 1054 71
rect 1254 71 1257 78
rect 1114 68 1257 71
rect 1314 68 1374 71
rect 1986 68 2038 71
rect 2042 68 2134 71
rect 2282 68 2318 71
rect 2322 68 2454 71
rect 2638 71 2641 78
rect 2506 68 2641 71
rect 382 62 385 68
rect 42 58 94 61
rect 98 58 142 61
rect 146 58 222 61
rect 226 58 382 61
rect 394 58 441 61
rect 642 58 702 61
rect 770 58 814 61
rect 866 58 894 61
rect 898 58 942 61
rect 1018 58 1030 61
rect 1034 58 1174 61
rect 1186 58 1206 61
rect 1210 58 1702 61
rect 1718 58 1774 61
rect 1910 61 1913 68
rect 1910 58 1958 61
rect 2026 58 2073 61
rect 2162 58 2286 61
rect 2338 58 2358 61
rect 2426 58 2518 61
rect 2554 58 2558 61
rect 438 52 441 58
rect 1718 52 1721 58
rect 2070 52 2073 58
rect -26 51 -22 52
rect -26 48 30 51
rect 90 48 150 51
rect 222 48 278 51
rect 834 48 870 51
rect 962 48 1134 51
rect 1170 48 1222 51
rect 1266 48 1270 51
rect 1362 48 1382 51
rect 1426 48 1545 51
rect 1866 48 1974 51
rect 1978 48 2006 51
rect 2398 51 2401 58
rect 2398 48 2462 51
rect 2610 48 2614 51
rect 2618 48 2654 51
rect 222 42 225 48
rect 1542 42 1545 48
rect -26 28 -22 32
rect 2734 28 2738 32
rect 838 12 841 18
rect 530 8 550 11
rect 576 3 578 7
rect 582 3 585 7
rect 590 3 592 7
rect 1600 3 1602 7
rect 1606 3 1609 7
rect 1614 3 1616 7
<< m4contact >>
rect 578 1803 582 1807
rect 586 1803 589 1807
rect 589 1803 590 1807
rect 1602 1803 1606 1807
rect 1610 1803 1613 1807
rect 1613 1803 1614 1807
rect 446 1798 450 1802
rect 742 1788 746 1792
rect 926 1748 930 1752
rect 2190 1748 2194 1752
rect 2238 1748 2242 1752
rect 1998 1738 2002 1742
rect 2230 1738 2234 1742
rect 2006 1728 2010 1732
rect 2534 1728 2538 1732
rect 142 1718 146 1722
rect 2158 1718 2162 1722
rect 2190 1708 2194 1712
rect 1082 1703 1086 1707
rect 1090 1703 1093 1707
rect 1093 1703 1094 1707
rect 2106 1703 2110 1707
rect 2114 1703 2117 1707
rect 2117 1703 2118 1707
rect 2150 1698 2154 1702
rect 2158 1698 2162 1702
rect 2222 1698 2226 1702
rect 2006 1688 2010 1692
rect 2446 1688 2450 1692
rect 2574 1688 2578 1692
rect 2702 1688 2706 1692
rect 454 1668 458 1672
rect 2326 1668 2330 1672
rect 926 1658 930 1662
rect 2462 1658 2466 1662
rect 2374 1648 2378 1652
rect 2382 1648 2386 1652
rect 2406 1648 2410 1652
rect 1998 1628 2002 1632
rect 1902 1618 1906 1622
rect 2662 1608 2666 1612
rect 578 1603 582 1607
rect 586 1603 589 1607
rect 589 1603 590 1607
rect 1602 1603 1606 1607
rect 1610 1603 1613 1607
rect 1613 1603 1614 1607
rect 2334 1588 2338 1592
rect 294 1568 298 1572
rect 38 1558 42 1562
rect 142 1558 146 1562
rect 502 1548 506 1552
rect 742 1548 746 1552
rect 1350 1538 1354 1542
rect 1798 1538 1802 1542
rect 2678 1538 2682 1542
rect 2414 1528 2418 1532
rect 2510 1528 2514 1532
rect 2542 1518 2546 1522
rect 1998 1508 2002 1512
rect 2382 1508 2386 1512
rect 1082 1503 1086 1507
rect 1090 1503 1093 1507
rect 1093 1503 1094 1507
rect 2106 1503 2110 1507
rect 2114 1503 2117 1507
rect 2117 1503 2118 1507
rect 294 1478 298 1482
rect 2158 1478 2162 1482
rect 1886 1468 1890 1472
rect 2134 1468 2138 1472
rect 2422 1468 2426 1472
rect 38 1458 42 1462
rect 1414 1458 1418 1462
rect 1422 1458 1426 1462
rect 2318 1458 2322 1462
rect 2510 1458 2514 1462
rect 2246 1448 2250 1452
rect 1902 1438 1906 1442
rect 2006 1418 2010 1422
rect 2582 1418 2586 1422
rect 578 1403 582 1407
rect 586 1403 589 1407
rect 589 1403 590 1407
rect 1602 1403 1606 1407
rect 1610 1403 1613 1407
rect 1613 1403 1614 1407
rect 390 1398 394 1402
rect 742 1398 746 1402
rect 1758 1398 1762 1402
rect 382 1388 386 1392
rect 502 1388 506 1392
rect 2006 1388 2010 1392
rect 2246 1388 2250 1392
rect 2582 1378 2586 1382
rect 1774 1368 1778 1372
rect 190 1358 194 1362
rect 270 1358 274 1362
rect 2414 1358 2418 1362
rect 126 1348 130 1352
rect 1174 1348 1178 1352
rect 2254 1348 2258 1352
rect 2422 1348 2426 1352
rect 2662 1348 2666 1352
rect 1766 1338 1770 1342
rect 1806 1338 1810 1342
rect 2086 1338 2090 1342
rect 2302 1338 2306 1342
rect 1174 1328 1178 1332
rect 2070 1328 2074 1332
rect 2254 1328 2258 1332
rect 2342 1328 2346 1332
rect 2622 1328 2626 1332
rect 2702 1328 2706 1332
rect 390 1318 394 1322
rect 2054 1318 2058 1322
rect 126 1308 130 1312
rect 886 1308 890 1312
rect 2302 1308 2306 1312
rect 2318 1308 2322 1312
rect 1082 1303 1086 1307
rect 1090 1303 1093 1307
rect 1093 1303 1094 1307
rect 2106 1303 2110 1307
rect 2114 1303 2117 1307
rect 2117 1303 2118 1307
rect 2430 1298 2434 1302
rect 1590 1288 1594 1292
rect 1134 1278 1138 1282
rect 1254 1278 1258 1282
rect 1262 1278 1266 1282
rect 1742 1278 1746 1282
rect 2174 1278 2178 1282
rect 190 1258 194 1262
rect 1462 1268 1466 1272
rect 2238 1268 2242 1272
rect 2494 1268 2498 1272
rect 2678 1268 2682 1272
rect 2054 1258 2058 1262
rect 2406 1258 2410 1262
rect 1134 1248 1138 1252
rect 270 1238 274 1242
rect 1214 1238 1218 1242
rect 1406 1238 1410 1242
rect 2214 1238 2218 1242
rect 2230 1238 2234 1242
rect 2350 1238 2354 1242
rect 974 1228 978 1232
rect 2174 1228 2178 1232
rect 2326 1218 2330 1222
rect 1214 1208 1218 1212
rect 578 1203 582 1207
rect 586 1203 589 1207
rect 589 1203 590 1207
rect 1602 1203 1606 1207
rect 1610 1203 1613 1207
rect 1613 1203 1614 1207
rect 950 1198 954 1202
rect 2302 1198 2306 1202
rect 2478 1198 2482 1202
rect 2430 1188 2434 1192
rect 1358 1178 1362 1182
rect 1862 1168 1866 1172
rect 1942 1168 1946 1172
rect 2390 1168 2394 1172
rect 2406 1168 2410 1172
rect 2422 1158 2426 1162
rect 750 1148 754 1152
rect 1334 1148 1338 1152
rect 1814 1148 1818 1152
rect 174 1138 178 1142
rect 310 1138 314 1142
rect 1366 1138 1370 1142
rect 1958 1138 1962 1142
rect 2006 1138 2010 1142
rect 2070 1138 2074 1142
rect 2302 1138 2306 1142
rect 2502 1138 2506 1142
rect 110 1128 114 1132
rect 270 1128 274 1132
rect 1334 1128 1338 1132
rect 2086 1128 2090 1132
rect 2574 1128 2578 1132
rect 1006 1118 1010 1122
rect 46 1108 50 1112
rect 630 1108 634 1112
rect 1894 1108 1898 1112
rect 2534 1108 2538 1112
rect 2614 1108 2618 1112
rect 1082 1103 1086 1107
rect 1090 1103 1093 1107
rect 1093 1103 1094 1107
rect 2106 1103 2110 1107
rect 2114 1103 2117 1107
rect 2117 1103 2118 1107
rect 1382 1098 1386 1102
rect 2006 1098 2010 1102
rect 2014 1098 2018 1102
rect 2438 1098 2442 1102
rect 2478 1098 2482 1102
rect 2006 1088 2010 1092
rect 2014 1078 2018 1082
rect 902 1068 906 1072
rect 1590 1068 1594 1072
rect 1742 1068 1746 1072
rect 1782 1068 1786 1072
rect 1822 1068 1826 1072
rect 2222 1068 2226 1072
rect 2302 1068 2306 1072
rect 46 1058 50 1062
rect 102 1058 106 1062
rect 1702 1058 1706 1062
rect 2198 1058 2202 1062
rect 2318 1058 2322 1062
rect 1006 1048 1010 1052
rect 1214 1048 1218 1052
rect 1414 1048 1418 1052
rect 142 1038 146 1042
rect 2238 1038 2242 1042
rect 2438 1018 2442 1022
rect 2478 1018 2482 1022
rect 578 1003 582 1007
rect 586 1003 589 1007
rect 589 1003 590 1007
rect 1602 1003 1606 1007
rect 1610 1003 1613 1007
rect 1613 1003 1614 1007
rect 1894 998 1898 1002
rect 2358 998 2362 1002
rect 982 988 986 992
rect 2494 988 2498 992
rect 1822 978 1826 982
rect 2662 978 2666 982
rect 6 968 10 972
rect 1038 968 1042 972
rect 2390 968 2394 972
rect 502 958 506 962
rect 1406 958 1410 962
rect 1622 958 1626 962
rect 1686 958 1690 962
rect 2350 958 2354 962
rect 6 948 10 952
rect 254 948 258 952
rect 494 948 498 952
rect 502 948 506 952
rect 750 948 754 952
rect 886 948 890 952
rect 950 948 954 952
rect 1254 948 1258 952
rect 2406 948 2410 952
rect 2534 948 2538 952
rect 222 938 226 942
rect 1382 938 1386 942
rect 2158 938 2162 942
rect 350 928 354 932
rect 558 928 562 932
rect 606 928 610 932
rect 1430 928 1434 932
rect 1798 928 1802 932
rect 2006 928 2010 932
rect 2542 928 2546 932
rect 1686 918 1690 922
rect 2382 918 2386 922
rect 2094 908 2098 912
rect 1082 903 1086 907
rect 1090 903 1093 907
rect 1093 903 1094 907
rect 2106 903 2110 907
rect 2114 903 2117 907
rect 2117 903 2118 907
rect 2590 898 2594 902
rect 302 888 306 892
rect 1590 888 1594 892
rect 270 878 274 882
rect 1886 888 1890 892
rect 1910 888 1914 892
rect 2518 888 2522 892
rect 2526 888 2530 892
rect 1958 878 1962 882
rect 2150 878 2154 882
rect 2678 878 2682 882
rect 902 868 906 872
rect 1702 868 1706 872
rect 2062 868 2066 872
rect 2254 868 2258 872
rect 2334 868 2338 872
rect 2550 868 2554 872
rect 2622 868 2626 872
rect 1958 858 1962 862
rect 2222 858 2226 862
rect 2238 858 2242 862
rect 110 848 114 852
rect 350 848 354 852
rect 2078 848 2082 852
rect 2198 848 2202 852
rect 2574 848 2578 852
rect 494 838 498 842
rect 1782 838 1786 842
rect 2054 838 2058 842
rect 2350 838 2354 842
rect 654 828 658 832
rect 1406 818 1410 822
rect 578 803 582 807
rect 586 803 589 807
rect 589 803 590 807
rect 1602 803 1606 807
rect 1610 803 1613 807
rect 1613 803 1614 807
rect 982 798 986 802
rect 558 788 562 792
rect 86 778 90 782
rect 182 778 186 782
rect 302 778 306 782
rect 126 768 130 772
rect 2294 768 2298 772
rect 2566 768 2570 772
rect 238 758 242 762
rect 1590 758 1594 762
rect 1942 758 1946 762
rect 2286 758 2290 762
rect 54 748 58 752
rect 94 748 98 752
rect 270 748 274 752
rect 286 748 290 752
rect 494 748 498 752
rect 1958 748 1962 752
rect 246 738 250 742
rect 702 738 706 742
rect 950 738 954 742
rect 1022 738 1026 742
rect 1886 738 1890 742
rect 2590 748 2594 752
rect 2070 738 2074 742
rect 2094 738 2098 742
rect 262 728 266 732
rect 598 728 602 732
rect 1038 728 1042 732
rect 1046 728 1050 732
rect 1798 728 1802 732
rect 2278 728 2282 732
rect 2638 728 2642 732
rect 134 718 138 722
rect 174 718 178 722
rect 230 718 234 722
rect 790 718 794 722
rect 886 718 890 722
rect 2214 718 2218 722
rect 2302 718 2306 722
rect 2438 718 2442 722
rect 2686 718 2690 722
rect 222 708 226 712
rect 310 708 314 712
rect 1622 708 1626 712
rect 2054 708 2058 712
rect 2270 708 2274 712
rect 1082 703 1086 707
rect 1090 703 1093 707
rect 1093 703 1094 707
rect 2106 703 2110 707
rect 2114 703 2117 707
rect 2117 703 2118 707
rect 254 688 258 692
rect 2046 688 2050 692
rect 182 678 186 682
rect 230 678 234 682
rect 1350 678 1354 682
rect 2006 678 2010 682
rect 86 668 90 672
rect 222 668 226 672
rect 2150 668 2154 672
rect 2382 668 2386 672
rect 206 658 210 662
rect 790 658 794 662
rect 974 658 978 662
rect 2382 658 2386 662
rect 2478 658 2482 662
rect 2662 658 2666 662
rect 318 648 322 652
rect 654 648 658 652
rect 2286 648 2290 652
rect 2294 648 2298 652
rect 86 638 90 642
rect 710 638 714 642
rect 1110 628 1114 632
rect 1422 618 1426 622
rect 578 603 582 607
rect 586 603 589 607
rect 589 603 590 607
rect 1602 603 1606 607
rect 1610 603 1613 607
rect 1613 603 1614 607
rect 1814 598 1818 602
rect 494 588 498 592
rect 1046 578 1050 582
rect 1326 568 1330 572
rect 206 558 210 562
rect 326 538 330 542
rect 366 538 370 542
rect 1302 548 1306 552
rect 2046 548 2050 552
rect 2334 548 2338 552
rect 2614 548 2618 552
rect 1326 538 1330 542
rect 822 528 826 532
rect 1246 528 1250 532
rect 1766 528 1770 532
rect 694 508 698 512
rect 2270 508 2274 512
rect 2550 508 2554 512
rect 1082 503 1086 507
rect 1090 503 1093 507
rect 1093 503 1094 507
rect 2106 503 2110 507
rect 2114 503 2117 507
rect 2117 503 2118 507
rect 718 498 722 502
rect 2278 498 2282 502
rect 638 488 642 492
rect 1214 488 1218 492
rect 2638 488 2642 492
rect 2534 478 2538 482
rect 142 468 146 472
rect 1478 468 1482 472
rect 318 448 322 452
rect 1294 448 1298 452
rect 1110 438 1114 442
rect 2526 438 2530 442
rect 1574 418 1578 422
rect 2598 418 2602 422
rect 822 408 826 412
rect 578 403 582 407
rect 586 403 589 407
rect 589 403 590 407
rect 1602 403 1606 407
rect 1610 403 1613 407
rect 1613 403 1614 407
rect 1062 388 1066 392
rect 2334 388 2338 392
rect 1110 378 1114 382
rect 1198 378 1202 382
rect 2590 378 2594 382
rect 1230 358 1234 362
rect 1294 358 1298 362
rect 1406 358 1410 362
rect 2542 358 2546 362
rect 158 348 162 352
rect 326 348 330 352
rect 1814 348 1818 352
rect 2246 348 2250 352
rect 2462 348 2466 352
rect 150 338 154 342
rect 990 338 994 342
rect 1238 338 1242 342
rect 2206 338 2210 342
rect 1422 328 1426 332
rect 1766 328 1770 332
rect 2422 328 2426 332
rect 2438 328 2442 332
rect 142 318 146 322
rect 1278 318 1282 322
rect 2246 318 2250 322
rect 2598 318 2602 322
rect 1854 308 1858 312
rect 2206 308 2210 312
rect 2374 308 2378 312
rect 1082 303 1086 307
rect 1090 303 1093 307
rect 1093 303 1094 307
rect 2106 303 2110 307
rect 2114 303 2117 307
rect 2117 303 2118 307
rect 206 298 210 302
rect 2518 298 2522 302
rect 1214 288 1218 292
rect 2382 288 2386 292
rect 222 278 226 282
rect 1190 278 1194 282
rect 2374 268 2378 272
rect 1278 258 1282 262
rect 2638 258 2642 262
rect 1102 248 1106 252
rect 1366 248 1370 252
rect 2422 238 2426 242
rect 2438 238 2442 242
rect 2574 218 2578 222
rect 990 208 994 212
rect 578 203 582 207
rect 586 203 589 207
rect 589 203 590 207
rect 1602 203 1606 207
rect 1610 203 1613 207
rect 1613 203 1614 207
rect 2382 188 2386 192
rect 678 168 682 172
rect 838 168 842 172
rect 1478 168 1482 172
rect 2070 168 2074 172
rect 1134 158 1138 162
rect 718 148 722 152
rect 918 148 922 152
rect 1222 148 1226 152
rect 1230 148 1234 152
rect 1574 148 1578 152
rect 2334 148 2338 152
rect 2462 148 2466 152
rect 670 138 674 142
rect 678 138 682 142
rect 894 138 898 142
rect 1478 138 1482 142
rect 2526 138 2530 142
rect 2590 138 2594 142
rect 950 128 954 132
rect 1006 128 1010 132
rect 1022 128 1026 132
rect 1198 128 1202 132
rect 2070 128 2074 132
rect 2566 128 2570 132
rect 1238 118 1242 122
rect 1246 118 1250 122
rect 1342 118 1346 122
rect 1054 108 1058 112
rect 2630 108 2634 112
rect 1082 103 1086 107
rect 1090 103 1093 107
rect 1093 103 1094 107
rect 2106 103 2110 107
rect 2114 103 2117 107
rect 2117 103 2118 107
rect 734 88 738 92
rect 1062 88 1066 92
rect 1174 78 1178 82
rect 1222 78 1226 82
rect 1310 78 1314 82
rect 2686 78 2690 82
rect 382 68 386 72
rect 702 68 706 72
rect 734 68 738 72
rect 806 68 810 72
rect 894 68 898 72
rect 990 68 994 72
rect 1038 68 1042 72
rect 1262 48 1266 52
rect 838 18 842 22
rect 578 3 582 7
rect 586 3 589 7
rect 589 3 590 7
rect 1602 3 1606 7
rect 1610 3 1613 7
rect 1613 3 1614 7
<< metal4 >>
rect 576 1803 578 1807
rect 582 1803 585 1807
rect 590 1803 592 1807
rect 1600 1803 1602 1807
rect 1606 1803 1609 1807
rect 1614 1803 1616 1807
rect 450 1798 457 1801
rect 142 1562 145 1718
rect 454 1672 457 1798
rect 576 1603 578 1607
rect 582 1603 585 1607
rect 590 1603 592 1607
rect 38 1462 41 1558
rect 294 1482 297 1568
rect 742 1552 745 1788
rect 2230 1748 2238 1751
rect 926 1662 929 1748
rect 1080 1703 1082 1707
rect 1086 1703 1089 1707
rect 1094 1703 1096 1707
rect 1998 1632 2001 1738
rect 2006 1692 2009 1728
rect 2104 1703 2106 1707
rect 2110 1703 2113 1707
rect 2118 1703 2120 1707
rect 2158 1702 2161 1718
rect 2190 1712 2193 1748
rect 2230 1742 2233 1748
rect 2146 1698 2150 1701
rect 2218 1698 2222 1701
rect 1600 1603 1602 1607
rect 1606 1603 1609 1607
rect 1614 1603 1616 1607
rect 126 1312 129 1348
rect 190 1262 193 1358
rect 270 1242 273 1358
rect 46 1062 49 1108
rect 94 1058 102 1061
rect 6 952 9 968
rect 86 772 89 778
rect 54 752 57 758
rect 94 752 97 1058
rect 110 852 113 1128
rect 134 1038 142 1041
rect 122 768 126 771
rect 134 722 137 1038
rect 174 722 177 1138
rect 262 1128 270 1131
rect 182 682 185 778
rect 222 712 225 938
rect 234 758 238 761
rect 246 742 249 748
rect 230 682 233 718
rect 254 692 257 948
rect 262 732 265 1128
rect 270 752 273 878
rect 302 782 305 888
rect 282 748 286 751
rect 310 712 313 1138
rect 350 852 353 928
rect 86 642 89 668
rect 206 562 209 658
rect 142 322 145 468
rect 150 348 158 351
rect 150 342 153 348
rect 206 302 209 558
rect 222 282 225 668
rect 318 452 321 648
rect 370 538 374 541
rect 326 352 329 538
rect 382 72 385 1388
rect 390 1322 393 1398
rect 502 1392 505 1548
rect 576 1403 578 1407
rect 582 1403 585 1407
rect 590 1403 592 1407
rect 742 1402 745 1548
rect 1080 1503 1082 1507
rect 1086 1503 1089 1507
rect 1094 1503 1096 1507
rect 1174 1332 1177 1348
rect 576 1203 578 1207
rect 582 1203 585 1207
rect 590 1203 592 1207
rect 634 1108 641 1111
rect 576 1003 578 1007
rect 582 1003 585 1007
rect 590 1003 592 1007
rect 502 952 505 958
rect 494 842 497 948
rect 598 928 606 931
rect 558 792 561 928
rect 576 803 578 807
rect 582 803 585 807
rect 590 803 592 807
rect 494 592 497 748
rect 598 732 601 928
rect 576 603 578 607
rect 582 603 585 607
rect 590 603 592 607
rect 638 492 641 1108
rect 750 952 753 1148
rect 886 952 889 1308
rect 1080 1303 1082 1307
rect 1086 1303 1089 1307
rect 1094 1303 1096 1307
rect 1134 1252 1137 1278
rect 654 652 657 828
rect 706 738 710 741
rect 886 722 889 948
rect 902 872 905 1068
rect 950 952 953 1198
rect 950 742 953 948
rect 790 662 793 718
rect 974 662 977 1228
rect 1214 1212 1217 1238
rect 1006 1052 1009 1118
rect 1080 1103 1082 1107
rect 1086 1103 1089 1107
rect 1094 1103 1096 1107
rect 1214 1052 1217 1208
rect 982 802 985 988
rect 1018 738 1022 741
rect 1038 732 1041 968
rect 1254 952 1257 1278
rect 1262 1272 1265 1278
rect 1334 1132 1337 1148
rect 1080 903 1082 907
rect 1086 903 1089 907
rect 1094 903 1096 907
rect 714 638 721 641
rect 576 403 578 407
rect 582 403 585 407
rect 590 403 592 407
rect 576 203 578 207
rect 582 203 585 207
rect 590 203 592 207
rect 670 142 673 148
rect 678 142 681 168
rect 694 71 697 508
rect 718 502 721 638
rect 1046 582 1049 728
rect 1080 703 1082 707
rect 1086 703 1089 707
rect 1094 703 1096 707
rect 1350 682 1353 1538
rect 1798 1532 1801 1538
rect 1890 1468 1894 1471
rect 1426 1458 1433 1461
rect 1358 1141 1361 1178
rect 1358 1138 1366 1141
rect 1382 942 1385 1098
rect 1406 962 1409 1238
rect 1414 1052 1417 1458
rect 1430 932 1433 1458
rect 1902 1442 1905 1618
rect 1998 1512 2001 1628
rect 2006 1422 2009 1688
rect 2104 1503 2106 1507
rect 2110 1503 2113 1507
rect 2118 1503 2120 1507
rect 2130 1468 2134 1471
rect 1600 1403 1602 1407
rect 1606 1403 1609 1407
rect 1614 1403 1616 1407
rect 1762 1398 1769 1401
rect 1766 1342 1769 1398
rect 1458 1268 1462 1271
rect 1590 1072 1593 1288
rect 1600 1203 1602 1207
rect 1606 1203 1609 1207
rect 1614 1203 1616 1207
rect 1742 1072 1745 1278
rect 1774 1071 1777 1368
rect 1806 1151 1809 1338
rect 1806 1148 1814 1151
rect 1774 1068 1782 1071
rect 1600 1003 1602 1007
rect 1606 1003 1609 1007
rect 1614 1003 1616 1007
rect 822 412 825 528
rect 1080 503 1082 507
rect 1086 503 1089 507
rect 1094 503 1096 507
rect 1110 442 1113 628
rect 990 212 993 338
rect 714 148 718 151
rect 734 72 737 88
rect 694 68 702 71
rect 810 68 814 71
rect 838 22 841 168
rect 922 148 926 151
rect 890 138 894 141
rect 1022 132 1025 138
rect 1010 128 1014 131
rect 950 122 953 128
rect 1046 108 1054 111
rect 1046 92 1049 108
rect 1062 92 1065 388
rect 1110 382 1113 438
rect 1190 378 1198 381
rect 1080 303 1082 307
rect 1086 303 1089 307
rect 1094 303 1096 307
rect 1190 282 1193 378
rect 1214 292 1217 488
rect 1106 248 1110 251
rect 1134 142 1137 158
rect 1230 152 1233 358
rect 1246 341 1249 528
rect 1302 451 1305 548
rect 1326 542 1329 568
rect 1350 542 1353 678
rect 1298 448 1305 451
rect 1294 362 1297 448
rect 1406 362 1409 818
rect 1590 762 1593 888
rect 1600 803 1602 807
rect 1606 803 1609 807
rect 1614 803 1616 807
rect 1622 712 1625 958
rect 1686 922 1689 958
rect 1702 872 1705 1058
rect 1782 842 1785 1068
rect 1822 982 1825 1068
rect 1798 732 1801 928
rect 1242 338 1249 341
rect 1422 332 1425 618
rect 1600 603 1602 607
rect 1606 603 1609 607
rect 1614 603 1616 607
rect 1278 262 1281 318
rect 1362 248 1366 251
rect 1478 172 1481 468
rect 1198 132 1201 138
rect 1080 103 1082 107
rect 1086 103 1089 107
rect 1094 103 1096 107
rect 1174 82 1177 128
rect 1222 82 1225 148
rect 1246 122 1249 148
rect 1478 142 1481 168
rect 1574 152 1577 418
rect 1600 403 1602 407
rect 1606 403 1609 407
rect 1614 403 1616 407
rect 1766 332 1769 528
rect 1814 352 1817 598
rect 1862 311 1865 1168
rect 1894 1002 1897 1108
rect 1882 888 1886 891
rect 1894 741 1897 998
rect 1902 891 1905 918
rect 1902 888 1910 891
rect 1942 762 1945 1168
rect 2006 1142 2009 1388
rect 2090 1338 2094 1341
rect 2054 1262 2057 1318
rect 2070 1142 2073 1328
rect 2104 1303 2106 1307
rect 2110 1303 2113 1307
rect 2118 1303 2120 1307
rect 1958 882 1961 1138
rect 2006 1102 2009 1138
rect 2006 932 2009 1088
rect 2014 1082 2017 1098
rect 1958 752 1961 858
rect 1890 738 1897 741
rect 2006 682 2009 928
rect 2066 868 2070 871
rect 2086 851 2089 1128
rect 2104 1103 2106 1107
rect 2110 1103 2113 1107
rect 2118 1103 2120 1107
rect 2158 942 2161 1478
rect 2246 1392 2249 1448
rect 2254 1332 2257 1348
rect 2302 1312 2305 1338
rect 2318 1312 2321 1458
rect 2174 1232 2177 1278
rect 2222 1238 2230 1241
rect 2082 848 2089 851
rect 2054 712 2057 838
rect 2094 742 2097 908
rect 2104 903 2106 907
rect 2110 903 2113 907
rect 2118 903 2120 907
rect 2074 738 2078 741
rect 2046 552 2049 688
rect 2054 672 2057 708
rect 2104 703 2106 707
rect 2110 703 2113 707
rect 2118 703 2120 707
rect 2150 672 2153 878
rect 2198 852 2201 1058
rect 2214 722 2217 1238
rect 2222 1072 2225 1238
rect 2238 1042 2241 1268
rect 2302 1202 2305 1308
rect 2306 1138 2310 1141
rect 2238 862 2241 888
rect 2254 862 2257 868
rect 2226 858 2230 861
rect 2270 512 2273 708
rect 2104 503 2106 507
rect 2110 503 2113 507
rect 2118 503 2120 507
rect 2278 502 2281 728
rect 2286 652 2289 758
rect 2294 652 2297 768
rect 2302 722 2305 1068
rect 2318 1062 2321 1308
rect 2326 1222 2329 1668
rect 2446 1662 2449 1688
rect 2466 1658 2470 1661
rect 2370 1648 2374 1651
rect 2402 1648 2406 1651
rect 2334 872 2337 1588
rect 2382 1512 2385 1648
rect 2414 1362 2417 1528
rect 2426 1468 2433 1471
rect 2342 1332 2345 1338
rect 2354 1238 2361 1241
rect 2358 1002 2361 1238
rect 2406 1172 2409 1258
rect 2390 972 2393 1168
rect 2334 552 2337 868
rect 2350 842 2353 958
rect 2406 952 2409 1168
rect 2422 1162 2425 1348
rect 2430 1302 2433 1468
rect 2510 1462 2513 1528
rect 2430 1192 2433 1298
rect 2478 1102 2481 1198
rect 2438 1022 2441 1098
rect 2378 918 2382 921
rect 2438 722 2441 738
rect 2382 662 2385 668
rect 2478 662 2481 1018
rect 2494 992 2497 1268
rect 2506 1138 2510 1141
rect 2534 1112 2537 1728
rect 2542 1522 2545 1528
rect 2334 392 2337 548
rect 1858 308 1865 311
rect 2206 312 2209 338
rect 2246 322 2249 348
rect 2104 303 2106 307
rect 2110 303 2113 307
rect 2118 303 2120 307
rect 1600 203 1602 207
rect 1606 203 1609 207
rect 1614 203 1616 207
rect 2070 132 2073 168
rect 2334 152 2337 388
rect 2374 272 2377 308
rect 2382 192 2385 288
rect 2422 242 2425 328
rect 2438 242 2441 328
rect 2462 152 2465 348
rect 2518 302 2521 888
rect 2526 872 2529 888
rect 2534 482 2537 948
rect 2542 932 2545 1518
rect 2574 1132 2577 1688
rect 2582 1382 2585 1418
rect 2662 1352 2665 1608
rect 2526 142 2529 438
rect 2542 362 2545 928
rect 2550 512 2553 868
rect 2566 132 2569 768
rect 2574 222 2577 848
rect 2590 752 2593 898
rect 2614 552 2617 1108
rect 2622 872 2625 1328
rect 2662 982 2665 1348
rect 2678 1272 2681 1538
rect 2702 1332 2705 1688
rect 2630 728 2638 731
rect 2590 142 2593 378
rect 2598 322 2601 418
rect 1338 118 1342 121
rect 1238 82 1241 118
rect 2630 112 2633 728
rect 2662 662 2665 978
rect 2678 882 2681 1268
rect 2638 262 2641 488
rect 2104 103 2106 107
rect 2110 103 2113 107
rect 2118 103 2120 107
rect 890 68 894 71
rect 994 68 998 71
rect 1034 68 1038 71
rect 1262 52 1265 88
rect 2686 82 2689 718
rect 1314 78 1318 81
rect 576 3 578 7
rect 582 3 585 7
rect 590 3 592 7
rect 1600 3 1602 7
rect 1606 3 1609 7
rect 1614 3 1616 7
<< m5contact >>
rect 578 1803 582 1807
rect 585 1803 586 1807
rect 586 1803 589 1807
rect 1602 1803 1606 1807
rect 1609 1803 1610 1807
rect 1610 1803 1613 1807
rect 578 1603 582 1607
rect 585 1603 586 1607
rect 586 1603 589 1607
rect 1082 1703 1086 1707
rect 1089 1703 1090 1707
rect 1090 1703 1093 1707
rect 2106 1703 2110 1707
rect 2113 1703 2114 1707
rect 2114 1703 2117 1707
rect 2142 1698 2146 1702
rect 2214 1698 2218 1702
rect 1602 1603 1606 1607
rect 1609 1603 1610 1607
rect 1610 1603 1613 1607
rect 86 768 90 772
rect 54 758 58 762
rect 118 768 122 772
rect 230 758 234 762
rect 246 748 250 752
rect 278 748 282 752
rect 374 538 378 542
rect 578 1403 582 1407
rect 585 1403 586 1407
rect 586 1403 589 1407
rect 1082 1503 1086 1507
rect 1089 1503 1090 1507
rect 1090 1503 1093 1507
rect 578 1203 582 1207
rect 585 1203 586 1207
rect 586 1203 589 1207
rect 578 1003 582 1007
rect 585 1003 586 1007
rect 586 1003 589 1007
rect 578 803 582 807
rect 585 803 586 807
rect 586 803 589 807
rect 578 603 582 607
rect 585 603 586 607
rect 586 603 589 607
rect 1082 1303 1086 1307
rect 1089 1303 1090 1307
rect 1090 1303 1093 1307
rect 710 738 714 742
rect 1082 1103 1086 1107
rect 1089 1103 1090 1107
rect 1090 1103 1093 1107
rect 1014 738 1018 742
rect 1262 1268 1266 1272
rect 1082 903 1086 907
rect 1089 903 1090 907
rect 1090 903 1093 907
rect 578 403 582 407
rect 585 403 586 407
rect 586 403 589 407
rect 578 203 582 207
rect 585 203 586 207
rect 586 203 589 207
rect 670 148 674 152
rect 1082 703 1086 707
rect 1089 703 1090 707
rect 1090 703 1093 707
rect 1798 1528 1802 1532
rect 1894 1468 1898 1472
rect 2106 1503 2110 1507
rect 2113 1503 2114 1507
rect 2114 1503 2117 1507
rect 2126 1468 2130 1472
rect 1602 1403 1606 1407
rect 1609 1403 1610 1407
rect 1610 1403 1613 1407
rect 1454 1268 1458 1272
rect 1602 1203 1606 1207
rect 1609 1203 1610 1207
rect 1610 1203 1613 1207
rect 1602 1003 1606 1007
rect 1609 1003 1610 1007
rect 1610 1003 1613 1007
rect 1082 503 1086 507
rect 1089 503 1090 507
rect 1090 503 1093 507
rect 710 148 714 152
rect 814 68 818 72
rect 926 148 930 152
rect 886 138 890 142
rect 1022 138 1026 142
rect 1014 128 1018 132
rect 950 118 954 122
rect 1082 303 1086 307
rect 1089 303 1090 307
rect 1090 303 1093 307
rect 1110 248 1114 252
rect 1350 538 1354 542
rect 1602 803 1606 807
rect 1609 803 1610 807
rect 1610 803 1613 807
rect 1602 603 1606 607
rect 1609 603 1610 607
rect 1610 603 1613 607
rect 1358 248 1362 252
rect 1246 148 1250 152
rect 1134 138 1138 142
rect 1198 138 1202 142
rect 1174 128 1178 132
rect 1082 103 1086 107
rect 1089 103 1090 107
rect 1090 103 1093 107
rect 1046 88 1050 92
rect 1602 403 1606 407
rect 1609 403 1610 407
rect 1610 403 1613 407
rect 1878 888 1882 892
rect 1902 918 1906 922
rect 2094 1338 2098 1342
rect 2106 1303 2110 1307
rect 2113 1303 2114 1307
rect 2114 1303 2117 1307
rect 2070 868 2074 872
rect 2106 1103 2110 1107
rect 2113 1103 2114 1107
rect 2114 1103 2117 1107
rect 2106 903 2110 907
rect 2113 903 2114 907
rect 2114 903 2117 907
rect 2078 738 2082 742
rect 2106 703 2110 707
rect 2113 703 2114 707
rect 2114 703 2117 707
rect 2310 1138 2314 1142
rect 2238 888 2242 892
rect 2230 858 2234 862
rect 2254 858 2258 862
rect 2054 668 2058 672
rect 2106 503 2110 507
rect 2113 503 2114 507
rect 2114 503 2117 507
rect 2446 1658 2450 1662
rect 2470 1658 2474 1662
rect 2366 1648 2370 1652
rect 2398 1648 2402 1652
rect 2342 1338 2346 1342
rect 2374 918 2378 922
rect 2438 738 2442 742
rect 2382 668 2386 672
rect 2510 1138 2514 1142
rect 2542 1528 2546 1532
rect 2106 303 2110 307
rect 2113 303 2114 307
rect 2114 303 2117 307
rect 1602 203 1606 207
rect 1609 203 1610 207
rect 1610 203 1613 207
rect 2526 868 2530 872
rect 1334 118 1338 122
rect 2106 103 2110 107
rect 2113 103 2114 107
rect 2114 103 2117 107
rect 1262 88 1266 92
rect 1238 78 1242 82
rect 886 68 890 72
rect 998 68 1002 72
rect 1030 68 1034 72
rect 1318 78 1322 82
rect 578 3 582 7
rect 585 3 586 7
rect 586 3 589 7
rect 1602 3 1606 7
rect 1609 3 1610 7
rect 1610 3 1613 7
<< metal5 >>
rect 582 1803 585 1807
rect 582 1802 586 1803
rect 1606 1803 1609 1807
rect 1606 1802 1610 1803
rect 1086 1703 1089 1707
rect 1086 1702 1090 1703
rect 2110 1703 2113 1707
rect 2110 1702 2114 1703
rect 2146 1698 2214 1701
rect 2450 1658 2470 1661
rect 2370 1648 2398 1651
rect 582 1603 585 1607
rect 582 1602 586 1603
rect 1606 1603 1609 1607
rect 1606 1602 1610 1603
rect 1802 1528 2542 1531
rect 1086 1503 1089 1507
rect 1086 1502 1090 1503
rect 2110 1503 2113 1507
rect 2110 1502 2114 1503
rect 1898 1468 2126 1471
rect 582 1403 585 1407
rect 582 1402 586 1403
rect 1606 1403 1609 1407
rect 1606 1402 1610 1403
rect 2098 1338 2342 1341
rect 1086 1303 1089 1307
rect 1086 1302 1090 1303
rect 2110 1303 2113 1307
rect 2110 1302 2114 1303
rect 1266 1268 1454 1271
rect 582 1203 585 1207
rect 582 1202 586 1203
rect 1606 1203 1609 1207
rect 1606 1202 1610 1203
rect 2314 1138 2510 1141
rect 1086 1103 1089 1107
rect 1086 1102 1090 1103
rect 2110 1103 2113 1107
rect 2110 1102 2114 1103
rect 582 1003 585 1007
rect 582 1002 586 1003
rect 1606 1003 1609 1007
rect 1606 1002 1610 1003
rect 1906 918 2374 921
rect 1086 903 1089 907
rect 1086 902 1090 903
rect 2110 903 2113 907
rect 2110 902 2114 903
rect 1882 888 2238 891
rect 2074 868 2526 871
rect 2234 858 2254 861
rect 582 803 585 807
rect 582 802 586 803
rect 1606 803 1609 807
rect 1606 802 1610 803
rect 90 768 118 771
rect 58 758 230 761
rect 250 748 278 751
rect 714 738 1014 741
rect 2082 738 2438 741
rect 1086 703 1089 707
rect 1086 702 1090 703
rect 2110 703 2113 707
rect 2110 702 2114 703
rect 2058 668 2382 671
rect 582 603 585 607
rect 582 602 586 603
rect 1606 603 1609 607
rect 1606 602 1610 603
rect 378 538 1350 541
rect 1086 503 1089 507
rect 1086 502 1090 503
rect 2110 503 2113 507
rect 2110 502 2114 503
rect 582 403 585 407
rect 582 402 586 403
rect 1606 403 1609 407
rect 1606 402 1610 403
rect 1086 303 1089 307
rect 1086 302 1090 303
rect 2110 303 2113 307
rect 2110 302 2114 303
rect 1114 248 1358 251
rect 582 203 585 207
rect 582 202 586 203
rect 1606 203 1609 207
rect 1606 202 1610 203
rect 674 148 710 151
rect 930 148 1246 151
rect 890 138 1022 141
rect 1138 138 1198 141
rect 1018 128 1174 131
rect 954 118 1334 121
rect 1086 103 1089 107
rect 1086 102 1090 103
rect 2110 103 2113 107
rect 2110 102 2114 103
rect 1050 88 1262 91
rect 1242 78 1318 81
rect 818 68 886 71
rect 1002 68 1030 71
rect 582 3 585 7
rect 582 2 586 3
rect 1606 3 1609 7
rect 1606 2 1610 3
<< m6contact >>
rect 576 1807 582 1808
rect 586 1807 592 1808
rect 576 1803 578 1807
rect 578 1803 582 1807
rect 586 1803 589 1807
rect 589 1803 592 1807
rect 576 1802 582 1803
rect 586 1802 592 1803
rect 1600 1807 1606 1808
rect 1610 1807 1616 1808
rect 1600 1803 1602 1807
rect 1602 1803 1606 1807
rect 1610 1803 1613 1807
rect 1613 1803 1616 1807
rect 1600 1802 1606 1803
rect 1610 1802 1616 1803
rect 1080 1707 1086 1708
rect 1090 1707 1096 1708
rect 1080 1703 1082 1707
rect 1082 1703 1086 1707
rect 1090 1703 1093 1707
rect 1093 1703 1096 1707
rect 1080 1702 1086 1703
rect 1090 1702 1096 1703
rect 2104 1707 2110 1708
rect 2114 1707 2120 1708
rect 2104 1703 2106 1707
rect 2106 1703 2110 1707
rect 2114 1703 2117 1707
rect 2117 1703 2120 1707
rect 2104 1702 2110 1703
rect 2114 1702 2120 1703
rect 576 1607 582 1608
rect 586 1607 592 1608
rect 576 1603 578 1607
rect 578 1603 582 1607
rect 586 1603 589 1607
rect 589 1603 592 1607
rect 576 1602 582 1603
rect 586 1602 592 1603
rect 1600 1607 1606 1608
rect 1610 1607 1616 1608
rect 1600 1603 1602 1607
rect 1602 1603 1606 1607
rect 1610 1603 1613 1607
rect 1613 1603 1616 1607
rect 1600 1602 1606 1603
rect 1610 1602 1616 1603
rect 1080 1507 1086 1508
rect 1090 1507 1096 1508
rect 1080 1503 1082 1507
rect 1082 1503 1086 1507
rect 1090 1503 1093 1507
rect 1093 1503 1096 1507
rect 1080 1502 1086 1503
rect 1090 1502 1096 1503
rect 2104 1507 2110 1508
rect 2114 1507 2120 1508
rect 2104 1503 2106 1507
rect 2106 1503 2110 1507
rect 2114 1503 2117 1507
rect 2117 1503 2120 1507
rect 2104 1502 2110 1503
rect 2114 1502 2120 1503
rect 576 1407 582 1408
rect 586 1407 592 1408
rect 576 1403 578 1407
rect 578 1403 582 1407
rect 586 1403 589 1407
rect 589 1403 592 1407
rect 576 1402 582 1403
rect 586 1402 592 1403
rect 1600 1407 1606 1408
rect 1610 1407 1616 1408
rect 1600 1403 1602 1407
rect 1602 1403 1606 1407
rect 1610 1403 1613 1407
rect 1613 1403 1616 1407
rect 1600 1402 1606 1403
rect 1610 1402 1616 1403
rect 1080 1307 1086 1308
rect 1090 1307 1096 1308
rect 1080 1303 1082 1307
rect 1082 1303 1086 1307
rect 1090 1303 1093 1307
rect 1093 1303 1096 1307
rect 1080 1302 1086 1303
rect 1090 1302 1096 1303
rect 2104 1307 2110 1308
rect 2114 1307 2120 1308
rect 2104 1303 2106 1307
rect 2106 1303 2110 1307
rect 2114 1303 2117 1307
rect 2117 1303 2120 1307
rect 2104 1302 2110 1303
rect 2114 1302 2120 1303
rect 576 1207 582 1208
rect 586 1207 592 1208
rect 576 1203 578 1207
rect 578 1203 582 1207
rect 586 1203 589 1207
rect 589 1203 592 1207
rect 576 1202 582 1203
rect 586 1202 592 1203
rect 1600 1207 1606 1208
rect 1610 1207 1616 1208
rect 1600 1203 1602 1207
rect 1602 1203 1606 1207
rect 1610 1203 1613 1207
rect 1613 1203 1616 1207
rect 1600 1202 1606 1203
rect 1610 1202 1616 1203
rect 1080 1107 1086 1108
rect 1090 1107 1096 1108
rect 1080 1103 1082 1107
rect 1082 1103 1086 1107
rect 1090 1103 1093 1107
rect 1093 1103 1096 1107
rect 1080 1102 1086 1103
rect 1090 1102 1096 1103
rect 2104 1107 2110 1108
rect 2114 1107 2120 1108
rect 2104 1103 2106 1107
rect 2106 1103 2110 1107
rect 2114 1103 2117 1107
rect 2117 1103 2120 1107
rect 2104 1102 2110 1103
rect 2114 1102 2120 1103
rect 576 1007 582 1008
rect 586 1007 592 1008
rect 576 1003 578 1007
rect 578 1003 582 1007
rect 586 1003 589 1007
rect 589 1003 592 1007
rect 576 1002 582 1003
rect 586 1002 592 1003
rect 1600 1007 1606 1008
rect 1610 1007 1616 1008
rect 1600 1003 1602 1007
rect 1602 1003 1606 1007
rect 1610 1003 1613 1007
rect 1613 1003 1616 1007
rect 1600 1002 1606 1003
rect 1610 1002 1616 1003
rect 1080 907 1086 908
rect 1090 907 1096 908
rect 1080 903 1082 907
rect 1082 903 1086 907
rect 1090 903 1093 907
rect 1093 903 1096 907
rect 1080 902 1086 903
rect 1090 902 1096 903
rect 2104 907 2110 908
rect 2114 907 2120 908
rect 2104 903 2106 907
rect 2106 903 2110 907
rect 2114 903 2117 907
rect 2117 903 2120 907
rect 2104 902 2110 903
rect 2114 902 2120 903
rect 576 807 582 808
rect 586 807 592 808
rect 576 803 578 807
rect 578 803 582 807
rect 586 803 589 807
rect 589 803 592 807
rect 576 802 582 803
rect 586 802 592 803
rect 1600 807 1606 808
rect 1610 807 1616 808
rect 1600 803 1602 807
rect 1602 803 1606 807
rect 1610 803 1613 807
rect 1613 803 1616 807
rect 1600 802 1606 803
rect 1610 802 1616 803
rect 1080 707 1086 708
rect 1090 707 1096 708
rect 1080 703 1082 707
rect 1082 703 1086 707
rect 1090 703 1093 707
rect 1093 703 1096 707
rect 1080 702 1086 703
rect 1090 702 1096 703
rect 2104 707 2110 708
rect 2114 707 2120 708
rect 2104 703 2106 707
rect 2106 703 2110 707
rect 2114 703 2117 707
rect 2117 703 2120 707
rect 2104 702 2110 703
rect 2114 702 2120 703
rect 576 607 582 608
rect 586 607 592 608
rect 576 603 578 607
rect 578 603 582 607
rect 586 603 589 607
rect 589 603 592 607
rect 576 602 582 603
rect 586 602 592 603
rect 1600 607 1606 608
rect 1610 607 1616 608
rect 1600 603 1602 607
rect 1602 603 1606 607
rect 1610 603 1613 607
rect 1613 603 1616 607
rect 1600 602 1606 603
rect 1610 602 1616 603
rect 1080 507 1086 508
rect 1090 507 1096 508
rect 1080 503 1082 507
rect 1082 503 1086 507
rect 1090 503 1093 507
rect 1093 503 1096 507
rect 1080 502 1086 503
rect 1090 502 1096 503
rect 2104 507 2110 508
rect 2114 507 2120 508
rect 2104 503 2106 507
rect 2106 503 2110 507
rect 2114 503 2117 507
rect 2117 503 2120 507
rect 2104 502 2110 503
rect 2114 502 2120 503
rect 576 407 582 408
rect 586 407 592 408
rect 576 403 578 407
rect 578 403 582 407
rect 586 403 589 407
rect 589 403 592 407
rect 576 402 582 403
rect 586 402 592 403
rect 1600 407 1606 408
rect 1610 407 1616 408
rect 1600 403 1602 407
rect 1602 403 1606 407
rect 1610 403 1613 407
rect 1613 403 1616 407
rect 1600 402 1606 403
rect 1610 402 1616 403
rect 1080 307 1086 308
rect 1090 307 1096 308
rect 1080 303 1082 307
rect 1082 303 1086 307
rect 1090 303 1093 307
rect 1093 303 1096 307
rect 1080 302 1086 303
rect 1090 302 1096 303
rect 2104 307 2110 308
rect 2114 307 2120 308
rect 2104 303 2106 307
rect 2106 303 2110 307
rect 2114 303 2117 307
rect 2117 303 2120 307
rect 2104 302 2110 303
rect 2114 302 2120 303
rect 576 207 582 208
rect 586 207 592 208
rect 576 203 578 207
rect 578 203 582 207
rect 586 203 589 207
rect 589 203 592 207
rect 576 202 582 203
rect 586 202 592 203
rect 1600 207 1606 208
rect 1610 207 1616 208
rect 1600 203 1602 207
rect 1602 203 1606 207
rect 1610 203 1613 207
rect 1613 203 1616 207
rect 1600 202 1606 203
rect 1610 202 1616 203
rect 1080 107 1086 108
rect 1090 107 1096 108
rect 1080 103 1082 107
rect 1082 103 1086 107
rect 1090 103 1093 107
rect 1093 103 1096 107
rect 1080 102 1086 103
rect 1090 102 1096 103
rect 2104 107 2110 108
rect 2114 107 2120 108
rect 2104 103 2106 107
rect 2106 103 2110 107
rect 2114 103 2117 107
rect 2117 103 2120 107
rect 2104 102 2110 103
rect 2114 102 2120 103
rect 576 7 582 8
rect 586 7 592 8
rect 576 3 578 7
rect 578 3 582 7
rect 586 3 589 7
rect 589 3 592 7
rect 576 2 582 3
rect 586 2 592 3
rect 1600 7 1606 8
rect 1610 7 1616 8
rect 1600 3 1602 7
rect 1602 3 1606 7
rect 1610 3 1613 7
rect 1613 3 1616 7
rect 1600 2 1606 3
rect 1610 2 1616 3
<< metal6 >>
rect 576 1808 592 1830
rect 582 1802 586 1808
rect 576 1608 592 1802
rect 582 1602 586 1608
rect 576 1408 592 1602
rect 582 1402 586 1408
rect 576 1208 592 1402
rect 582 1202 586 1208
rect 576 1008 592 1202
rect 582 1002 586 1008
rect 576 808 592 1002
rect 582 802 586 808
rect 576 608 592 802
rect 582 602 586 608
rect 576 408 592 602
rect 582 402 586 408
rect 576 208 592 402
rect 582 202 586 208
rect 576 8 592 202
rect 582 2 586 8
rect 576 -30 592 2
rect 1080 1708 1096 1830
rect 1086 1702 1090 1708
rect 1080 1508 1096 1702
rect 1086 1502 1090 1508
rect 1080 1308 1096 1502
rect 1086 1302 1090 1308
rect 1080 1108 1096 1302
rect 1086 1102 1090 1108
rect 1080 908 1096 1102
rect 1086 902 1090 908
rect 1080 708 1096 902
rect 1086 702 1090 708
rect 1080 508 1096 702
rect 1086 502 1090 508
rect 1080 308 1096 502
rect 1086 302 1090 308
rect 1080 108 1096 302
rect 1086 102 1090 108
rect 1080 -30 1096 102
rect 1600 1808 1616 1830
rect 1606 1802 1610 1808
rect 1600 1608 1616 1802
rect 1606 1602 1610 1608
rect 1600 1408 1616 1602
rect 1606 1402 1610 1408
rect 1600 1208 1616 1402
rect 1606 1202 1610 1208
rect 1600 1008 1616 1202
rect 1606 1002 1610 1008
rect 1600 808 1616 1002
rect 1606 802 1610 808
rect 1600 608 1616 802
rect 1606 602 1610 608
rect 1600 408 1616 602
rect 1606 402 1610 408
rect 1600 208 1616 402
rect 1606 202 1610 208
rect 1600 8 1616 202
rect 1606 2 1610 8
rect 1600 -30 1616 2
rect 2104 1708 2120 1830
rect 2110 1702 2114 1708
rect 2104 1508 2120 1702
rect 2110 1502 2114 1508
rect 2104 1308 2120 1502
rect 2110 1302 2114 1308
rect 2104 1108 2120 1302
rect 2110 1102 2114 1108
rect 2104 908 2120 1102
rect 2110 902 2114 908
rect 2104 708 2120 902
rect 2110 702 2114 708
rect 2104 508 2120 702
rect 2110 502 2114 508
rect 2104 308 2120 502
rect 2110 302 2114 308
rect 2104 108 2120 302
rect 2110 102 2114 108
rect 2104 -30 2120 102
use INVX1  INVX1_78
timestamp 1626400951
transform 1 0 4 0 1 1705
box -2 -3 18 103
use OAI22X1  OAI22X1_4
timestamp 1626400951
transform 1 0 20 0 1 1705
box -2 -3 42 103
use NAND2X1  NAND2X1_35
timestamp 1626400951
transform -1 0 84 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_36
timestamp 1626400951
transform -1 0 108 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_79
timestamp 1626400951
transform -1 0 124 0 1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_32
timestamp 1626400951
transform 1 0 124 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_74
timestamp 1626400951
transform -1 0 164 0 1 1705
box -2 -3 18 103
use INVX1  INVX1_45
timestamp 1626400951
transform 1 0 164 0 1 1705
box -2 -3 18 103
use AOI22X1  AOI22X1_6
timestamp 1626400951
transform -1 0 220 0 1 1705
box -2 -3 42 103
use INVX1  INVX1_44
timestamp 1626400951
transform -1 0 236 0 1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_46
timestamp 1626400951
transform -1 0 260 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_46
timestamp 1626400951
transform 1 0 260 0 1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_12
timestamp 1626400951
transform -1 0 300 0 1 1705
box -2 -3 26 103
use OR2X2  OR2X2_4
timestamp 1626400951
transform 1 0 300 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_69
timestamp 1626400951
transform 1 0 332 0 1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_30
timestamp 1626400951
transform -1 0 372 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_70
timestamp 1626400951
transform 1 0 372 0 1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_31
timestamp 1626400951
transform -1 0 412 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_41
timestamp 1626400951
transform 1 0 412 0 1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_10
timestamp 1626400951
transform -1 0 452 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_11
timestamp 1626400951
transform 1 0 452 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_42
timestamp 1626400951
transform -1 0 492 0 1 1705
box -2 -3 18 103
use BUFX2  BUFX2_9
timestamp 1626400951
transform 1 0 492 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_18
timestamp 1626400951
transform -1 0 612 0 1 1705
box -2 -3 98 103
use FILL  FILL_17_0_0
timestamp 1626400951
transform 1 0 612 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_0_1
timestamp 1626400951
transform 1 0 620 0 1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_16
timestamp 1626400951
transform 1 0 628 0 1 1705
box -2 -3 98 103
use BUFX2  BUFX2_7
timestamp 1626400951
transform 1 0 724 0 1 1705
box -2 -3 26 103
use BUFX2  BUFX2_4
timestamp 1626400951
transform 1 0 748 0 1 1705
box -2 -3 26 103
use BUFX2  BUFX2_6
timestamp 1626400951
transform 1 0 772 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_33
timestamp 1626400951
transform 1 0 796 0 1 1705
box -2 -3 98 103
use INVX1  INVX1_15
timestamp 1626400951
transform 1 0 892 0 1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_15
timestamp 1626400951
transform 1 0 908 0 1 1705
box -2 -3 26 103
use BUFX2  BUFX2_24
timestamp 1626400951
transform 1 0 932 0 1 1705
box -2 -3 26 103
use BUFX2  BUFX2_13
timestamp 1626400951
transform 1 0 956 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_14
timestamp 1626400951
transform 1 0 980 0 1 1705
box -2 -3 98 103
use BUFX2  BUFX2_10
timestamp 1626400951
transform 1 0 1076 0 1 1705
box -2 -3 26 103
use FILL  FILL_17_1_0
timestamp 1626400951
transform 1 0 1100 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_1_1
timestamp 1626400951
transform 1 0 1108 0 1 1705
box -2 -3 10 103
use BUFX2  BUFX2_5
timestamp 1626400951
transform 1 0 1116 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_31
timestamp 1626400951
transform -1 0 1236 0 1 1705
box -2 -3 98 103
use BUFX2  BUFX2_21
timestamp 1626400951
transform -1 0 1260 0 1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_13
timestamp 1626400951
transform -1 0 1284 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_13
timestamp 1626400951
transform -1 0 1300 0 1 1705
box -2 -3 18 103
use BUFX2  BUFX2_22
timestamp 1626400951
transform 1 0 1300 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_17
timestamp 1626400951
transform 1 0 1324 0 1 1705
box -2 -3 98 103
use BUFX2  BUFX2_26
timestamp 1626400951
transform 1 0 1420 0 1 1705
box -2 -3 26 103
use BUFX2  BUFX2_25
timestamp 1626400951
transform 1 0 1444 0 1 1705
box -2 -3 26 103
use BUFX2  BUFX2_8
timestamp 1626400951
transform 1 0 1468 0 1 1705
box -2 -3 26 103
use BUFX2  BUFX2_18
timestamp 1626400951
transform 1 0 1492 0 1 1705
box -2 -3 26 103
use BUFX2  BUFX2_2
timestamp 1626400951
transform -1 0 1540 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_37
timestamp 1626400951
transform -1 0 1636 0 1 1705
box -2 -3 98 103
use FILL  FILL_17_2_0
timestamp 1626400951
transform 1 0 1636 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_2_1
timestamp 1626400951
transform 1 0 1644 0 1 1705
box -2 -3 10 103
use INVX1  INVX1_3
timestamp 1626400951
transform 1 0 1652 0 1 1705
box -2 -3 18 103
use BUFX2  BUFX2_28
timestamp 1626400951
transform 1 0 1668 0 1 1705
box -2 -3 26 103
use BUFX2  BUFX2_20
timestamp 1626400951
transform -1 0 1716 0 1 1705
box -2 -3 26 103
use BUFX2  BUFX2_31
timestamp 1626400951
transform 1 0 1716 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_25
timestamp 1626400951
transform 1 0 1740 0 1 1705
box -2 -3 98 103
use NOR2X1  NOR2X1_22
timestamp 1626400951
transform -1 0 1860 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_24
timestamp 1626400951
transform -1 0 1876 0 1 1705
box -2 -3 18 103
use BUFX2  BUFX2_16
timestamp 1626400951
transform 1 0 1876 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_130
timestamp 1626400951
transform 1 0 1900 0 1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_137
timestamp 1626400951
transform 1 0 1996 0 1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_90
timestamp 1626400951
transform 1 0 2028 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_134
timestamp 1626400951
transform 1 0 2060 0 1 1705
box -2 -3 98 103
use FILL  FILL_17_3_0
timestamp 1626400951
transform -1 0 2164 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_3_1
timestamp 1626400951
transform -1 0 2172 0 1 1705
box -2 -3 10 103
use NOR2X1  NOR2X1_177
timestamp 1626400951
transform -1 0 2196 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_138
timestamp 1626400951
transform 1 0 2196 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_126
timestamp 1626400951
transform -1 0 2252 0 1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_91
timestamp 1626400951
transform 1 0 2252 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_133
timestamp 1626400951
transform 1 0 2284 0 1 1705
box -2 -3 98 103
use NAND2X1  NAND2X1_108
timestamp 1626400951
transform 1 0 2380 0 1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_163
timestamp 1626400951
transform 1 0 2404 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_182
timestamp 1626400951
transform 1 0 2428 0 1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_164
timestamp 1626400951
transform -1 0 2468 0 1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_165
timestamp 1626400951
transform -1 0 2492 0 1 1705
box -2 -3 26 103
use AND2X2  AND2X2_20
timestamp 1626400951
transform 1 0 2492 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_21
timestamp 1626400951
transform -1 0 2548 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_163
timestamp 1626400951
transform 1 0 2548 0 1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_24
timestamp 1626400951
transform 1 0 2564 0 1 1705
box -2 -3 98 103
use INVX1  INVX1_23
timestamp 1626400951
transform -1 0 2676 0 1 1705
box -2 -3 18 103
use BUFX2  BUFX2_15
timestamp 1626400951
transform 1 0 2676 0 1 1705
box -2 -3 26 103
use FILL  FILL_18_1
timestamp 1626400951
transform 1 0 2700 0 1 1705
box -2 -3 10 103
use BUFX2  BUFX2_39
timestamp 1626400951
transform 1 0 4 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_49
timestamp 1626400951
transform -1 0 60 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_76
timestamp 1626400951
transform 1 0 60 0 -1 1705
box -2 -3 18 103
use NAND3X1  NAND3X1_26
timestamp 1626400951
transform 1 0 76 0 -1 1705
box -2 -3 34 103
use AOI22X1  AOI22X1_13
timestamp 1626400951
transform 1 0 108 0 -1 1705
box -2 -3 42 103
use INVX1  INVX1_77
timestamp 1626400951
transform -1 0 164 0 -1 1705
box -2 -3 18 103
use INVX1  INVX1_75
timestamp 1626400951
transform -1 0 180 0 -1 1705
box -2 -3 18 103
use INVX1  INVX1_73
timestamp 1626400951
transform 1 0 180 0 -1 1705
box -2 -3 18 103
use AOI22X1  AOI22X1_12
timestamp 1626400951
transform -1 0 236 0 -1 1705
box -2 -3 42 103
use NOR2X1  NOR2X1_63
timestamp 1626400951
transform 1 0 236 0 -1 1705
box -2 -3 26 103
use INVX1  INVX1_72
timestamp 1626400951
transform -1 0 276 0 -1 1705
box -2 -3 18 103
use NAND3X1  NAND3X1_20
timestamp 1626400951
transform 1 0 276 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_47
timestamp 1626400951
transform 1 0 308 0 -1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_13
timestamp 1626400951
transform -1 0 348 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_39
timestamp 1626400951
transform 1 0 348 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_71
timestamp 1626400951
transform 1 0 380 0 -1 1705
box -2 -3 18 103
use INVX2  INVX2_4
timestamp 1626400951
transform 1 0 396 0 -1 1705
box -2 -3 18 103
use NAND3X1  NAND3X1_19
timestamp 1626400951
transform -1 0 444 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_43
timestamp 1626400951
transform 1 0 444 0 -1 1705
box -2 -3 18 103
use AOI22X1  AOI22X1_5
timestamp 1626400951
transform -1 0 500 0 -1 1705
box -2 -3 42 103
use INVX2  INVX2_2
timestamp 1626400951
transform 1 0 500 0 -1 1705
box -2 -3 18 103
use AOI21X1  AOI21X1_37
timestamp 1626400951
transform -1 0 548 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_47
timestamp 1626400951
transform -1 0 572 0 -1 1705
box -2 -3 26 103
use FILL  FILL_16_0_0
timestamp 1626400951
transform 1 0 572 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_0_1
timestamp 1626400951
transform 1 0 580 0 -1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_38
timestamp 1626400951
transform 1 0 588 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_33
timestamp 1626400951
transform 1 0 620 0 -1 1705
box -2 -3 18 103
use AOI21X1  AOI21X1_24
timestamp 1626400951
transform 1 0 636 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_22
timestamp 1626400951
transform -1 0 700 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_31
timestamp 1626400951
transform -1 0 716 0 -1 1705
box -2 -3 18 103
use AOI21X1  AOI21X1_21
timestamp 1626400951
transform -1 0 748 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_30
timestamp 1626400951
transform -1 0 764 0 -1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_15
timestamp 1626400951
transform -1 0 860 0 -1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_22
timestamp 1626400951
transform 1 0 860 0 -1 1705
box -2 -3 98 103
use INVX1  INVX1_21
timestamp 1626400951
transform 1 0 956 0 -1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_19
timestamp 1626400951
transform 1 0 972 0 -1 1705
box -2 -3 26 103
use AOI22X1  AOI22X1_3
timestamp 1626400951
transform -1 0 1036 0 -1 1705
box -2 -3 42 103
use INVX1  INVX1_17
timestamp 1626400951
transform -1 0 1052 0 -1 1705
box -2 -3 18 103
use FILL  FILL_16_1_0
timestamp 1626400951
transform 1 0 1052 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_1_1
timestamp 1626400951
transform 1 0 1060 0 -1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_19
timestamp 1626400951
transform 1 0 1068 0 -1 1705
box -2 -3 98 103
use INVX1  INVX1_29
timestamp 1626400951
transform 1 0 1164 0 -1 1705
box -2 -3 18 103
use AOI21X1  AOI21X1_20
timestamp 1626400951
transform 1 0 1180 0 -1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_30
timestamp 1626400951
transform -1 0 1308 0 -1 1705
box -2 -3 98 103
use INVX1  INVX1_12
timestamp 1626400951
transform 1 0 1308 0 -1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_12
timestamp 1626400951
transform 1 0 1324 0 -1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_23
timestamp 1626400951
transform -1 0 1380 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_32
timestamp 1626400951
transform -1 0 1396 0 -1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_16
timestamp 1626400951
transform -1 0 1420 0 -1 1705
box -2 -3 26 103
use INVX1  INVX1_16
timestamp 1626400951
transform -1 0 1436 0 -1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_34
timestamp 1626400951
transform -1 0 1532 0 -1 1705
box -2 -3 98 103
use INVX1  INVX1_26
timestamp 1626400951
transform 1 0 1532 0 -1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_11
timestamp 1626400951
transform -1 0 1644 0 -1 1705
box -2 -3 98 103
use FILL  FILL_16_2_0
timestamp 1626400951
transform 1 0 1644 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_2_1
timestamp 1626400951
transform 1 0 1652 0 -1 1705
box -2 -3 10 103
use NOR2X1  NOR2X1_4
timestamp 1626400951
transform 1 0 1660 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_11
timestamp 1626400951
transform -1 0 1708 0 -1 1705
box -2 -3 26 103
use INVX1  INVX1_11
timestamp 1626400951
transform -1 0 1724 0 -1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_29
timestamp 1626400951
transform 1 0 1724 0 -1 1705
box -2 -3 98 103
use NOR2X1  NOR2X1_7
timestamp 1626400951
transform -1 0 1844 0 -1 1705
box -2 -3 26 103
use INVX1  INVX1_6
timestamp 1626400951
transform -1 0 1860 0 -1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_40
timestamp 1626400951
transform -1 0 1956 0 -1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_131
timestamp 1626400951
transform 1 0 1956 0 -1 1705
box -2 -3 98 103
use AOI21X1  AOI21X1_94
timestamp 1626400951
transform -1 0 2084 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_180
timestamp 1626400951
transform 1 0 2084 0 -1 1705
box -2 -3 26 103
use FILL  FILL_16_3_0
timestamp 1626400951
transform -1 0 2116 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_3_1
timestamp 1626400951
transform -1 0 2124 0 -1 1705
box -2 -3 10 103
use NAND2X1  NAND2X1_130
timestamp 1626400951
transform -1 0 2148 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_141
timestamp 1626400951
transform -1 0 2180 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_176
timestamp 1626400951
transform 1 0 2180 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_125
timestamp 1626400951
transform -1 0 2228 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_107
timestamp 1626400951
transform 1 0 2228 0 -1 1705
box -2 -3 26 103
use INVX1  INVX1_181
timestamp 1626400951
transform 1 0 2252 0 -1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_160
timestamp 1626400951
transform 1 0 2268 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_119
timestamp 1626400951
transform 1 0 2292 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_120
timestamp 1626400951
transform 1 0 2324 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_121
timestamp 1626400951
transform 1 0 2356 0 -1 1705
box -2 -3 34 103
use OAI22X1  OAI22X1_8
timestamp 1626400951
transform -1 0 2428 0 -1 1705
box -2 -3 42 103
use AND2X2  AND2X2_19
timestamp 1626400951
transform -1 0 2460 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_122
timestamp 1626400951
transform 1 0 2460 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_31
timestamp 1626400951
transform -1 0 2524 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_123
timestamp 1626400951
transform 1 0 2524 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_77
timestamp 1626400951
transform -1 0 2588 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_76
timestamp 1626400951
transform -1 0 2620 0 -1 1705
box -2 -3 34 103
use XOR2X1  XOR2X1_10
timestamp 1626400951
transform -1 0 2676 0 -1 1705
box -2 -3 58 103
use BUFX4  BUFX4_33
timestamp 1626400951
transform 1 0 2676 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_49
timestamp 1626400951
transform 1 0 4 0 1 1505
box -2 -3 18 103
use AOI22X1  AOI22X1_7
timestamp 1626400951
transform -1 0 60 0 1 1505
box -2 -3 42 103
use INVX1  INVX1_48
timestamp 1626400951
transform -1 0 76 0 1 1505
box -2 -3 18 103
use INVX1  INVX1_51
timestamp 1626400951
transform 1 0 76 0 1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_16
timestamp 1626400951
transform -1 0 116 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_33
timestamp 1626400951
transform 1 0 116 0 1 1505
box -2 -3 26 103
use NAND3X1  NAND3X1_24
timestamp 1626400951
transform 1 0 140 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_51
timestamp 1626400951
transform -1 0 196 0 1 1505
box -2 -3 26 103
use OR2X2  OR2X2_7
timestamp 1626400951
transform 1 0 196 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_52
timestamp 1626400951
transform 1 0 228 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_34
timestamp 1626400951
transform 1 0 260 0 1 1505
box -2 -3 26 103
use NAND3X1  NAND3X1_23
timestamp 1626400951
transform -1 0 316 0 1 1505
box -2 -3 34 103
use AOI22X1  AOI22X1_11
timestamp 1626400951
transform 1 0 316 0 1 1505
box -2 -3 42 103
use AOI21X1  AOI21X1_46
timestamp 1626400951
transform 1 0 356 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_64
timestamp 1626400951
transform -1 0 412 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_51
timestamp 1626400951
transform 1 0 412 0 1 1505
box -2 -3 34 103
use BUFX2  BUFX2_11
timestamp 1626400951
transform -1 0 468 0 1 1505
box -2 -3 26 103
use INVX1  INVX1_19
timestamp 1626400951
transform 1 0 468 0 1 1505
box -2 -3 18 103
use NOR2X1  NOR2X1_17
timestamp 1626400951
transform 1 0 484 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_20
timestamp 1626400951
transform -1 0 604 0 1 1505
box -2 -3 98 103
use FILL  FILL_15_0_0
timestamp 1626400951
transform 1 0 604 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_0_1
timestamp 1626400951
transform 1 0 612 0 1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_13
timestamp 1626400951
transform 1 0 620 0 1 1505
box -2 -3 98 103
use BUFX4  BUFX4_44
timestamp 1626400951
transform -1 0 748 0 1 1505
box -2 -3 34 103
use BUFX2  BUFX2_27
timestamp 1626400951
transform 1 0 748 0 1 1505
box -2 -3 26 103
use INVX1  INVX1_2
timestamp 1626400951
transform 1 0 772 0 1 1505
box -2 -3 18 103
use NOR2X1  NOR2X1_3
timestamp 1626400951
transform 1 0 788 0 1 1505
box -2 -3 26 103
use BUFX4  BUFX4_40
timestamp 1626400951
transform -1 0 844 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_17
timestamp 1626400951
transform -1 0 876 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_2
timestamp 1626400951
transform -1 0 900 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_20
timestamp 1626400951
transform 1 0 900 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_6
timestamp 1626400951
transform 1 0 932 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_27
timestamp 1626400951
transform -1 0 980 0 1 1505
box -2 -3 26 103
use INVX1  INVX1_34
timestamp 1626400951
transform 1 0 980 0 1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_5
timestamp 1626400951
transform 1 0 996 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_24
timestamp 1626400951
transform -1 0 1044 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_21
timestamp 1626400951
transform -1 0 1076 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_3
timestamp 1626400951
transform -1 0 1100 0 1 1505
box -2 -3 26 103
use FILL  FILL_15_1_0
timestamp 1626400951
transform -1 0 1108 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_1_1
timestamp 1626400951
transform -1 0 1116 0 1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_3
timestamp 1626400951
transform -1 0 1212 0 1 1505
box -2 -3 98 103
use BUFX2  BUFX2_1
timestamp 1626400951
transform -1 0 1236 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_35
timestamp 1626400951
transform 1 0 1236 0 1 1505
box -2 -3 98 103
use OR2X2  OR2X2_1
timestamp 1626400951
transform 1 0 1332 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_18
timestamp 1626400951
transform -1 0 1396 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_27
timestamp 1626400951
transform -1 0 1412 0 1 1505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_12
timestamp 1626400951
transform 1 0 1412 0 1 1505
box -2 -3 98 103
use AOI22X1  AOI22X1_4
timestamp 1626400951
transform -1 0 1548 0 1 1505
box -2 -3 42 103
use BUFX2  BUFX2_3
timestamp 1626400951
transform 1 0 1548 0 1 1505
box -2 -3 26 103
use FILL  FILL_15_2_0
timestamp 1626400951
transform -1 0 1580 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_2_1
timestamp 1626400951
transform -1 0 1588 0 1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_136
timestamp 1626400951
transform -1 0 1684 0 1 1505
box -2 -3 98 103
use AOI21X1  AOI21X1_103
timestamp 1626400951
transform -1 0 1716 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_150
timestamp 1626400951
transform -1 0 1748 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_192
timestamp 1626400951
transform -1 0 1772 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_140
timestamp 1626400951
transform -1 0 1796 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_109
timestamp 1626400951
transform 1 0 1796 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_169
timestamp 1626400951
transform 1 0 1820 0 1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_93
timestamp 1626400951
transform -1 0 1876 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_140
timestamp 1626400951
transform -1 0 1908 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_178
timestamp 1626400951
transform -1 0 1932 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_139
timestamp 1626400951
transform 1 0 1932 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_92
timestamp 1626400951
transform 1 0 1964 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_128
timestamp 1626400951
transform -1 0 2020 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_132
timestamp 1626400951
transform 1 0 2020 0 1 1505
box -2 -3 98 103
use FILL  FILL_15_3_0
timestamp 1626400951
transform -1 0 2124 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_3_1
timestamp 1626400951
transform -1 0 2132 0 1 1505
box -2 -3 10 103
use AND2X2  AND2X2_21
timestamp 1626400951
transform -1 0 2164 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_167
timestamp 1626400951
transform 1 0 2164 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_125
timestamp 1626400951
transform 1 0 2188 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_126
timestamp 1626400951
transform 1 0 2220 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_171
timestamp 1626400951
transform -1 0 2268 0 1 1505
box -2 -3 18 103
use NOR2X1  NOR2X1_166
timestamp 1626400951
transform -1 0 2292 0 1 1505
box -2 -3 26 103
use BUFX4  BUFX4_30
timestamp 1626400951
transform 1 0 2292 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_152
timestamp 1626400951
transform 1 0 2324 0 1 1505
box -2 -3 26 103
use XNOR2X1  XNOR2X1_24
timestamp 1626400951
transform -1 0 2404 0 1 1505
box -2 -3 58 103
use NOR2X1  NOR2X1_162
timestamp 1626400951
transform -1 0 2428 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_150
timestamp 1626400951
transform -1 0 2452 0 1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_75
timestamp 1626400951
transform 1 0 2452 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_114
timestamp 1626400951
transform 1 0 2484 0 1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_71
timestamp 1626400951
transform -1 0 2540 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_124
timestamp 1626400951
transform 1 0 2540 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_143
timestamp 1626400951
transform -1 0 2596 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_144
timestamp 1626400951
transform 1 0 2596 0 1 1505
box -2 -3 26 103
use INVX1  INVX1_168
timestamp 1626400951
transform -1 0 2636 0 1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_100
timestamp 1626400951
transform -1 0 2660 0 1 1505
box -2 -3 26 103
use OR2X2  OR2X2_18
timestamp 1626400951
transform -1 0 2692 0 1 1505
box -2 -3 34 103
use FILL  FILL_16_1
timestamp 1626400951
transform 1 0 2692 0 1 1505
box -2 -3 10 103
use FILL  FILL_16_2
timestamp 1626400951
transform 1 0 2700 0 1 1505
box -2 -3 10 103
use NOR2X1  NOR2X1_52
timestamp 1626400951
transform 1 0 4 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_50
timestamp 1626400951
transform 1 0 28 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_36
timestamp 1626400951
transform 1 0 60 0 -1 1505
box -2 -3 34 103
use OAI22X1  OAI22X1_2
timestamp 1626400951
transform -1 0 132 0 -1 1505
box -2 -3 42 103
use INVX1  INVX1_50
timestamp 1626400951
transform 1 0 132 0 -1 1505
box -2 -3 18 103
use NAND3X1  NAND3X1_22
timestamp 1626400951
transform -1 0 180 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_15
timestamp 1626400951
transform -1 0 204 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_37
timestamp 1626400951
transform 1 0 204 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_47
timestamp 1626400951
transform 1 0 236 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_38
timestamp 1626400951
transform 1 0 268 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_64
timestamp 1626400951
transform 1 0 300 0 -1 1505
box -2 -3 98 103
use INVX1  INVX1_217
timestamp 1626400951
transform 1 0 396 0 -1 1505
box -2 -3 18 103
use OAI22X1  OAI22X1_11
timestamp 1626400951
transform 1 0 412 0 -1 1505
box -2 -3 42 103
use INVX1  INVX1_218
timestamp 1626400951
transform -1 0 468 0 -1 1505
box -2 -3 18 103
use NOR3X1  NOR3X1_7
timestamp 1626400951
transform -1 0 532 0 -1 1505
box -2 -3 66 103
use OAI21X1  OAI21X1_164
timestamp 1626400951
transform -1 0 564 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_219
timestamp 1626400951
transform -1 0 580 0 -1 1505
box -2 -3 18 103
use FILL  FILL_14_0_0
timestamp 1626400951
transform -1 0 588 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_0_1
timestamp 1626400951
transform -1 0 596 0 -1 1505
box -2 -3 10 103
use INVX1  INVX1_28
timestamp 1626400951
transform -1 0 612 0 -1 1505
box -2 -3 18 103
use AOI21X1  AOI21X1_19
timestamp 1626400951
transform 1 0 612 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_147
timestamp 1626400951
transform 1 0 644 0 -1 1505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_36
timestamp 1626400951
transform -1 0 836 0 -1 1505
box -2 -3 98 103
use NAND2X1  NAND2X1_2
timestamp 1626400951
transform -1 0 860 0 -1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_5
timestamp 1626400951
transform 1 0 860 0 -1 1505
box -2 -3 98 103
use NOR2X1  NOR2X1_28
timestamp 1626400951
transform 1 0 956 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_22
timestamp 1626400951
transform -1 0 1012 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_35
timestamp 1626400951
transform -1 0 1028 0 -1 1505
box -2 -3 18 103
use NAND3X1  NAND3X1_17
timestamp 1626400951
transform 1 0 1028 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_4
timestamp 1626400951
transform -1 0 1084 0 -1 1505
box -2 -3 26 103
use FILL  FILL_14_1_0
timestamp 1626400951
transform 1 0 1084 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_1_1
timestamp 1626400951
transform 1 0 1092 0 -1 1505
box -2 -3 10 103
use NOR2X1  NOR2X1_26
timestamp 1626400951
transform 1 0 1100 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_1
timestamp 1626400951
transform 1 0 1124 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_1
timestamp 1626400951
transform 1 0 1148 0 -1 1505
box -2 -3 26 103
use NAND3X1  NAND3X1_48
timestamp 1626400951
transform 1 0 1172 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_220
timestamp 1626400951
transform -1 0 1220 0 -1 1505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_4
timestamp 1626400951
transform -1 0 1316 0 -1 1505
box -2 -3 98 103
use INVX2  INVX2_1
timestamp 1626400951
transform 1 0 1316 0 -1 1505
box -2 -3 18 103
use AOI21X1  AOI21X1_17
timestamp 1626400951
transform 1 0 1332 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_1
timestamp 1626400951
transform 1 0 1364 0 -1 1505
box -2 -3 18 103
use AOI22X1  AOI22X1_1
timestamp 1626400951
transform 1 0 1380 0 -1 1505
box -2 -3 42 103
use AOI22X1  AOI22X1_2
timestamp 1626400951
transform -1 0 1460 0 -1 1505
box -2 -3 42 103
use INVX1  INVX1_9
timestamp 1626400951
transform -1 0 1476 0 -1 1505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_27
timestamp 1626400951
transform -1 0 1572 0 -1 1505
box -2 -3 98 103
use BUFX4  BUFX4_39
timestamp 1626400951
transform -1 0 1604 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_2_0
timestamp 1626400951
transform 1 0 1604 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_2_1
timestamp 1626400951
transform 1 0 1612 0 -1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_137
timestamp 1626400951
transform 1 0 1620 0 -1 1505
box -2 -3 98 103
use INVX1  INVX1_195
timestamp 1626400951
transform 1 0 1716 0 -1 1505
box -2 -3 18 103
use NOR2X1  NOR2X1_174
timestamp 1626400951
transform 1 0 1732 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_135
timestamp 1626400951
transform -1 0 1788 0 -1 1505
box -2 -3 34 103
use AND2X2  AND2X2_22
timestamp 1626400951
transform -1 0 1820 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_183
timestamp 1626400951
transform 1 0 1820 0 -1 1505
box -2 -3 18 103
use NOR2X1  NOR2X1_170
timestamp 1626400951
transform -1 0 1860 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_171
timestamp 1626400951
transform 1 0 1860 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_127
timestamp 1626400951
transform 1 0 1884 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_175
timestamp 1626400951
transform 1 0 1916 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_136
timestamp 1626400951
transform 1 0 1940 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_135
timestamp 1626400951
transform -1 0 2068 0 -1 1505
box -2 -3 98 103
use AOI21X1  AOI21X1_89
timestamp 1626400951
transform -1 0 2100 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_123
timestamp 1626400951
transform -1 0 2124 0 -1 1505
box -2 -3 26 103
use FILL  FILL_14_3_0
timestamp 1626400951
transform 1 0 2124 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_3_1
timestamp 1626400951
transform 1 0 2132 0 -1 1505
box -2 -3 10 103
use AOI21X1  AOI21X1_78
timestamp 1626400951
transform 1 0 2140 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_79
timestamp 1626400951
transform 1 0 2172 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_128
timestamp 1626400951
transform -1 0 2236 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_168
timestamp 1626400951
transform -1 0 2260 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_149
timestamp 1626400951
transform 1 0 2260 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_145
timestamp 1626400951
transform -1 0 2308 0 -1 1505
box -2 -3 26 103
use BUFX4  BUFX4_48
timestamp 1626400951
transform 1 0 2308 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_47
timestamp 1626400951
transform 1 0 2340 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_151
timestamp 1626400951
transform -1 0 2396 0 -1 1505
box -2 -3 26 103
use INVX1  INVX1_169
timestamp 1626400951
transform 1 0 2396 0 -1 1505
box -2 -3 18 103
use NOR2X1  NOR2X1_142
timestamp 1626400951
transform -1 0 2436 0 -1 1505
box -2 -3 26 103
use NAND3X1  NAND3X1_36
timestamp 1626400951
transform 1 0 2436 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_161
timestamp 1626400951
transform -1 0 2492 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_105
timestamp 1626400951
transform -1 0 2524 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_106
timestamp 1626400951
transform -1 0 2556 0 -1 1505
box -2 -3 34 103
use AND2X2  AND2X2_18
timestamp 1626400951
transform -1 0 2588 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_146
timestamp 1626400951
transform 1 0 2588 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_103
timestamp 1626400951
transform -1 0 2644 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_141
timestamp 1626400951
transform -1 0 2668 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_98
timestamp 1626400951
transform 1 0 2668 0 -1 1505
box -2 -3 26 103
use INVX1  INVX1_167
timestamp 1626400951
transform -1 0 2708 0 -1 1505
box -2 -3 18 103
use NAND3X1  NAND3X1_25
timestamp 1626400951
transform -1 0 36 0 1 1305
box -2 -3 34 103
use OR2X2  OR2X2_6
timestamp 1626400951
transform -1 0 68 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_34
timestamp 1626400951
transform -1 0 92 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_62
timestamp 1626400951
transform -1 0 116 0 1 1305
box -2 -3 26 103
use INVX2  INVX2_5
timestamp 1626400951
transform -1 0 132 0 1 1305
box -2 -3 18 103
use INVX2  INVX2_3
timestamp 1626400951
transform 1 0 132 0 1 1305
box -2 -3 18 103
use NAND2X1  NAND2X1_14
timestamp 1626400951
transform 1 0 148 0 1 1305
box -2 -3 26 103
use OR2X2  OR2X2_3
timestamp 1626400951
transform 1 0 172 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_21
timestamp 1626400951
transform 1 0 204 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_35
timestamp 1626400951
transform -1 0 260 0 1 1305
box -2 -3 26 103
use AND2X2  AND2X2_7
timestamp 1626400951
transform -1 0 292 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_44
timestamp 1626400951
transform 1 0 292 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_56
timestamp 1626400951
transform 1 0 316 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_57
timestamp 1626400951
transform -1 0 380 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_94
timestamp 1626400951
transform -1 0 396 0 1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_66
timestamp 1626400951
transform 1 0 396 0 1 1305
box -2 -3 98 103
use NOR2X1  NOR2X1_206
timestamp 1626400951
transform 1 0 492 0 1 1305
box -2 -3 26 103
use AND2X2  AND2X2_37
timestamp 1626400951
transform 1 0 516 0 1 1305
box -2 -3 34 103
use OAI22X1  OAI22X1_10
timestamp 1626400951
transform -1 0 588 0 1 1305
box -2 -3 42 103
use FILL  FILL_13_0_0
timestamp 1626400951
transform 1 0 588 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_0_1
timestamp 1626400951
transform 1 0 596 0 1 1305
box -2 -3 10 103
use INVX1  INVX1_216
timestamp 1626400951
transform 1 0 604 0 1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_65
timestamp 1626400951
transform -1 0 716 0 1 1305
box -2 -3 98 103
use BUFX4  BUFX4_43
timestamp 1626400951
transform -1 0 748 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_62
timestamp 1626400951
transform -1 0 844 0 1 1305
box -2 -3 98 103
use BUFX4  BUFX4_38
timestamp 1626400951
transform -1 0 876 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_18
timestamp 1626400951
transform 1 0 876 0 1 1305
box -2 -3 18 103
use BUFX2  BUFX2_35
timestamp 1626400951
transform 1 0 892 0 1 1305
box -2 -3 26 103
use CLKBUF1  CLKBUF1_11
timestamp 1626400951
transform -1 0 988 0 1 1305
box -2 -3 74 103
use INVX1  INVX1_221
timestamp 1626400951
transform 1 0 988 0 1 1305
box -2 -3 18 103
use NAND2X1  NAND2X1_152
timestamp 1626400951
transform 1 0 1004 0 1 1305
box -2 -3 26 103
use NOR3X1  NOR3X1_8
timestamp 1626400951
transform -1 0 1092 0 1 1305
box -2 -3 66 103
use FILL  FILL_13_1_0
timestamp 1626400951
transform -1 0 1100 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_1_1
timestamp 1626400951
transform -1 0 1108 0 1 1305
box -2 -3 10 103
use NOR2X1  NOR2X1_29
timestamp 1626400951
transform -1 0 1132 0 1 1305
box -2 -3 26 103
use AND2X2  AND2X2_2
timestamp 1626400951
transform 1 0 1132 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_32
timestamp 1626400951
transform -1 0 1188 0 1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_6
timestamp 1626400951
transform -1 0 1284 0 1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_60
timestamp 1626400951
transform -1 0 1380 0 1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_43
timestamp 1626400951
transform -1 0 1476 0 1 1305
box -2 -3 98 103
use BUFX2  BUFX2_41
timestamp 1626400951
transform 1 0 1476 0 1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_8
timestamp 1626400951
transform -1 0 1596 0 1 1305
box -2 -3 98 103
use FILL  FILL_13_2_0
timestamp 1626400951
transform 1 0 1596 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_2_1
timestamp 1626400951
transform 1 0 1604 0 1 1305
box -2 -3 10 103
use CLKBUF1  CLKBUF1_10
timestamp 1626400951
transform 1 0 1612 0 1 1305
box -2 -3 74 103
use CLKBUF1  CLKBUF1_12
timestamp 1626400951
transform 1 0 1684 0 1 1305
box -2 -3 74 103
use NAND3X1  NAND3X1_41
timestamp 1626400951
transform 1 0 1756 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_37
timestamp 1626400951
transform 1 0 1788 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_21
timestamp 1626400951
transform 1 0 1820 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_19
timestamp 1626400951
transform 1 0 1852 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_20
timestamp 1626400951
transform 1 0 1884 0 1 1305
box -2 -3 34 103
use INVX4  INVX4_2
timestamp 1626400951
transform -1 0 1940 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_179
timestamp 1626400951
transform 1 0 1940 0 1 1305
box -2 -3 26 103
use NAND3X1  NAND3X1_42
timestamp 1626400951
transform 1 0 1964 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_196
timestamp 1626400951
transform -1 0 2012 0 1 1305
box -2 -3 18 103
use NAND2X1  NAND2X1_129
timestamp 1626400951
transform -1 0 2036 0 1 1305
box -2 -3 26 103
use INVX1  INVX1_149
timestamp 1626400951
transform 1 0 2036 0 1 1305
box -2 -3 18 103
use NOR2X1  NOR2X1_116
timestamp 1626400951
transform -1 0 2076 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_131
timestamp 1626400951
transform -1 0 2108 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_3_0
timestamp 1626400951
transform -1 0 2116 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_3_1
timestamp 1626400951
transform -1 0 2124 0 1 1305
box -2 -3 10 103
use AOI21X1  AOI21X1_80
timestamp 1626400951
transform -1 0 2156 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_78
timestamp 1626400951
transform 1 0 2156 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_99
timestamp 1626400951
transform 1 0 2180 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_101
timestamp 1626400951
transform 1 0 2204 0 1 1305
box -2 -3 26 103
use INVX1  INVX1_184
timestamp 1626400951
transform -1 0 2244 0 1 1305
box -2 -3 18 103
use NAND2X1  NAND2X1_80
timestamp 1626400951
transform 1 0 2244 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_81
timestamp 1626400951
transform 1 0 2268 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_82
timestamp 1626400951
transform 1 0 2292 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_96
timestamp 1626400951
transform 1 0 2316 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_97
timestamp 1626400951
transform 1 0 2340 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_115
timestamp 1626400951
transform 1 0 2364 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_136
timestamp 1626400951
transform 1 0 2388 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_140
timestamp 1626400951
transform -1 0 2436 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_102
timestamp 1626400951
transform -1 0 2468 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_101
timestamp 1626400951
transform 1 0 2468 0 1 1305
box -2 -3 34 103
use OAI22X1  OAI22X1_7
timestamp 1626400951
transform 1 0 2500 0 1 1305
box -2 -3 42 103
use OAI21X1  OAI21X1_104
timestamp 1626400951
transform 1 0 2540 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_100
timestamp 1626400951
transform -1 0 2604 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_138
timestamp 1626400951
transform -1 0 2628 0 1 1305
box -2 -3 26 103
use AND2X2  AND2X2_17
timestamp 1626400951
transform -1 0 2660 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_32
timestamp 1626400951
transform 1 0 2660 0 1 1305
box -2 -3 34 103
use FILL  FILL_14_1
timestamp 1626400951
transform 1 0 2692 0 1 1305
box -2 -3 10 103
use FILL  FILL_14_2
timestamp 1626400951
transform 1 0 2700 0 1 1305
box -2 -3 10 103
use XNOR2X1  XNOR2X1_7
timestamp 1626400951
transform 1 0 4 0 -1 1305
box -2 -3 58 103
use AOI21X1  AOI21X1_45
timestamp 1626400951
transform 1 0 60 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_61
timestamp 1626400951
transform 1 0 92 0 -1 1305
box -2 -3 26 103
use INVX1  INVX1_91
timestamp 1626400951
transform -1 0 132 0 -1 1305
box -2 -3 18 103
use XNOR2X1  XNOR2X1_1
timestamp 1626400951
transform 1 0 132 0 -1 1305
box -2 -3 58 103
use NOR2X1  NOR2X1_45
timestamp 1626400951
transform -1 0 212 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_36
timestamp 1626400951
transform 1 0 212 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_63
timestamp 1626400951
transform 1 0 244 0 -1 1305
box -2 -3 18 103
use NOR2X1  NOR2X1_44
timestamp 1626400951
transform -1 0 284 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_54
timestamp 1626400951
transform 1 0 284 0 -1 1305
box -2 -3 34 103
use AOI22X1  AOI22X1_16
timestamp 1626400951
transform -1 0 356 0 -1 1305
box -2 -3 42 103
use INVX1  INVX1_92
timestamp 1626400951
transform 1 0 356 0 -1 1305
box -2 -3 18 103
use NAND2X1  NAND2X1_43
timestamp 1626400951
transform -1 0 396 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_44
timestamp 1626400951
transform -1 0 428 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_66
timestamp 1626400951
transform -1 0 444 0 -1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_63
timestamp 1626400951
transform 1 0 444 0 -1 1305
box -2 -3 98 103
use AND2X2  AND2X2_9
timestamp 1626400951
transform 1 0 540 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_0_0
timestamp 1626400951
transform -1 0 580 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_0_1
timestamp 1626400951
transform -1 0 588 0 -1 1305
box -2 -3 10 103
use OR2X2  OR2X2_8
timestamp 1626400951
transform -1 0 620 0 -1 1305
box -2 -3 34 103
use OR2X2  OR2X2_5
timestamp 1626400951
transform 1 0 620 0 -1 1305
box -2 -3 34 103
use AND2X2  AND2X2_6
timestamp 1626400951
transform 1 0 652 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_56
timestamp 1626400951
transform -1 0 780 0 -1 1305
box -2 -3 98 103
use AOI21X1  AOI21X1_13
timestamp 1626400951
transform -1 0 812 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_13
timestamp 1626400951
transform -1 0 844 0 -1 1305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_8
timestamp 1626400951
transform 1 0 844 0 -1 1305
box -2 -3 74 103
use NOR2X1  NOR2X1_25
timestamp 1626400951
transform 1 0 916 0 -1 1305
box -2 -3 26 103
use BUFX4  BUFX4_22
timestamp 1626400951
transform -1 0 972 0 -1 1305
box -2 -3 34 103
use AND2X2  AND2X2_3
timestamp 1626400951
transform 1 0 972 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_7
timestamp 1626400951
transform 1 0 1004 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_23
timestamp 1626400951
transform 1 0 1028 0 -1 1305
box -2 -3 34 103
use OR2X2  OR2X2_2
timestamp 1626400951
transform 1 0 1060 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_1_0
timestamp 1626400951
transform -1 0 1100 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_1_1
timestamp 1626400951
transform -1 0 1108 0 -1 1305
box -2 -3 10 103
use NAND2X1  NAND2X1_151
timestamp 1626400951
transform -1 0 1132 0 -1 1305
box -2 -3 26 103
use NAND3X1  NAND3X1_1
timestamp 1626400951
transform 1 0 1132 0 -1 1305
box -2 -3 34 103
use AND2X2  AND2X2_1
timestamp 1626400951
transform -1 0 1196 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_222
timestamp 1626400951
transform -1 0 1212 0 -1 1305
box -2 -3 18 103
use NOR2X1  NOR2X1_209
timestamp 1626400951
transform -1 0 1236 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_28
timestamp 1626400951
transform 1 0 1236 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_33
timestamp 1626400951
transform 1 0 1268 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_7
timestamp 1626400951
transform 1 0 1292 0 -1 1305
box -2 -3 98 103
use AOI21X1  AOI21X1_25
timestamp 1626400951
transform 1 0 1388 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_24
timestamp 1626400951
transform -1 0 1452 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_207
timestamp 1626400951
transform -1 0 1476 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_26
timestamp 1626400951
transform 1 0 1476 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_8
timestamp 1626400951
transform 1 0 1508 0 -1 1305
box -2 -3 26 103
use INVX1  INVX1_36
timestamp 1626400951
transform -1 0 1548 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_25
timestamp 1626400951
transform 1 0 1548 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_30
timestamp 1626400951
transform -1 0 1604 0 -1 1305
box -2 -3 26 103
use FILL  FILL_12_2_0
timestamp 1626400951
transform 1 0 1604 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_2_1
timestamp 1626400951
transform 1 0 1612 0 -1 1305
box -2 -3 10 103
use BUFX4  BUFX4_42
timestamp 1626400951
transform 1 0 1620 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_110
timestamp 1626400951
transform 1 0 1652 0 -1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_127
timestamp 1626400951
transform -1 0 1772 0 -1 1305
box -2 -3 26 103
use BUFX4  BUFX4_18
timestamp 1626400951
transform -1 0 1804 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_121
timestamp 1626400951
transform -1 0 1828 0 -1 1305
box -2 -3 26 103
use BUFX4  BUFX4_17
timestamp 1626400951
transform -1 0 1860 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_124
timestamp 1626400951
transform -1 0 1884 0 -1 1305
box -2 -3 26 103
use INVX2  INVX2_14
timestamp 1626400951
transform 1 0 1884 0 -1 1305
box -2 -3 18 103
use NAND2X1  NAND2X1_122
timestamp 1626400951
transform -1 0 1924 0 -1 1305
box -2 -3 26 103
use NAND3X1  NAND3X1_45
timestamp 1626400951
transform -1 0 1956 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_105
timestamp 1626400951
transform -1 0 2052 0 -1 1305
box -2 -3 98 103
use NOR2X1  NOR2X1_112
timestamp 1626400951
transform 1 0 2052 0 -1 1305
box -2 -3 26 103
use INVX2  INVX2_10
timestamp 1626400951
transform 1 0 2076 0 -1 1305
box -2 -3 18 103
use INVX2  INVX2_11
timestamp 1626400951
transform 1 0 2092 0 -1 1305
box -2 -3 18 103
use FILL  FILL_12_3_0
timestamp 1626400951
transform 1 0 2108 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_3_1
timestamp 1626400951
transform 1 0 2116 0 -1 1305
box -2 -3 10 103
use NOR2X1  NOR2X1_113
timestamp 1626400951
transform 1 0 2124 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_129
timestamp 1626400951
transform 1 0 2148 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_72
timestamp 1626400951
transform -1 0 2204 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_148
timestamp 1626400951
transform 1 0 2204 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_119
timestamp 1626400951
transform 1 0 2228 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_79
timestamp 1626400951
transform 1 0 2252 0 -1 1305
box -2 -3 26 103
use INVX2  INVX2_12
timestamp 1626400951
transform 1 0 2276 0 -1 1305
box -2 -3 18 103
use INVX8  INVX8_2
timestamp 1626400951
transform -1 0 2332 0 -1 1305
box -2 -3 42 103
use NOR2X1  NOR2X1_118
timestamp 1626400951
transform -1 0 2356 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_117
timestamp 1626400951
transform 1 0 2356 0 -1 1305
box -2 -3 26 103
use INVX1  INVX1_165
timestamp 1626400951
transform 1 0 2380 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_98
timestamp 1626400951
transform 1 0 2396 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_151
timestamp 1626400951
transform 1 0 2428 0 -1 1305
box -2 -3 18 103
use NOR2X1  NOR2X1_139
timestamp 1626400951
transform -1 0 2468 0 -1 1305
box -2 -3 26 103
use INVX1  INVX1_166
timestamp 1626400951
transform -1 0 2484 0 -1 1305
box -2 -3 18 103
use NOR2X1  NOR2X1_137
timestamp 1626400951
transform -1 0 2508 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_99
timestamp 1626400951
transform 1 0 2508 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_164
timestamp 1626400951
transform -1 0 2556 0 -1 1305
box -2 -3 18 103
use AOI21X1  AOI21X1_70
timestamp 1626400951
transform -1 0 2588 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_152
timestamp 1626400951
transform 1 0 2588 0 -1 1305
box -2 -3 18 103
use AOI21X1  AOI21X1_69
timestamp 1626400951
transform 1 0 2604 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_68
timestamp 1626400951
transform -1 0 2668 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_95
timestamp 1626400951
transform -1 0 2692 0 -1 1305
box -2 -3 26 103
use FILL  FILL_13_1
timestamp 1626400951
transform -1 0 2700 0 -1 1305
box -2 -3 10 103
use FILL  FILL_13_2
timestamp 1626400951
transform -1 0 2708 0 -1 1305
box -2 -3 10 103
use INVX1  INVX1_90
timestamp 1626400951
transform 1 0 4 0 1 1105
box -2 -3 18 103
use NOR2X1  NOR2X1_60
timestamp 1626400951
transform -1 0 44 0 1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_44
timestamp 1626400951
transform 1 0 44 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_59
timestamp 1626400951
transform 1 0 76 0 1 1105
box -2 -3 26 103
use INVX1  INVX1_89
timestamp 1626400951
transform -1 0 116 0 1 1105
box -2 -3 18 103
use XNOR2X1  XNOR2X1_8
timestamp 1626400951
transform -1 0 172 0 1 1105
box -2 -3 58 103
use OAI21X1  OAI21X1_48
timestamp 1626400951
transform 1 0 172 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_24
timestamp 1626400951
transform 1 0 204 0 1 1105
box -2 -3 26 103
use AND2X2  AND2X2_4
timestamp 1626400951
transform 1 0 228 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_43
timestamp 1626400951
transform 1 0 260 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_41
timestamp 1626400951
transform 1 0 292 0 1 1105
box -2 -3 34 103
use AOI22X1  AOI22X1_10
timestamp 1626400951
transform -1 0 364 0 1 1105
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_61
timestamp 1626400951
transform 1 0 364 0 1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_23
timestamp 1626400951
transform 1 0 460 0 1 1105
box -2 -3 26 103
use INVX1  INVX1_64
timestamp 1626400951
transform -1 0 500 0 1 1105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_80
timestamp 1626400951
transform 1 0 500 0 1 1105
box -2 -3 98 103
use FILL  FILL_11_0_0
timestamp 1626400951
transform -1 0 604 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_0_1
timestamp 1626400951
transform -1 0 612 0 1 1105
box -2 -3 10 103
use OR2X2  OR2X2_14
timestamp 1626400951
transform -1 0 644 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_96
timestamp 1626400951
transform 1 0 644 0 1 1105
box -2 -3 98 103
use NAND3X1  NAND3X1_13
timestamp 1626400951
transform 1 0 740 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_58
timestamp 1626400951
transform -1 0 868 0 1 1105
box -2 -3 98 103
use NOR2X1  NOR2X1_93
timestamp 1626400951
transform -1 0 892 0 1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_82
timestamp 1626400951
transform 1 0 892 0 1 1105
box -2 -3 98 103
use INVX1  INVX1_118
timestamp 1626400951
transform -1 0 1004 0 1 1105
box -2 -3 18 103
use INVX1  INVX1_125
timestamp 1626400951
transform 1 0 1004 0 1 1105
box -2 -3 18 103
use AOI22X1  AOI22X1_18
timestamp 1626400951
transform -1 0 1060 0 1 1105
box -2 -3 42 103
use NOR2X1  NOR2X1_107
timestamp 1626400951
transform -1 0 1084 0 1 1105
box -2 -3 26 103
use FILL  FILL_11_1_0
timestamp 1626400951
transform -1 0 1092 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_1_1
timestamp 1626400951
transform -1 0 1100 0 1 1105
box -2 -3 10 103
use INVX1  INVX1_124
timestamp 1626400951
transform -1 0 1116 0 1 1105
box -2 -3 18 103
use INVX1  INVX1_123
timestamp 1626400951
transform -1 0 1132 0 1 1105
box -2 -3 18 103
use NAND2X1  NAND2X1_60
timestamp 1626400951
transform 1 0 1132 0 1 1105
box -2 -3 26 103
use INVX1  INVX1_126
timestamp 1626400951
transform -1 0 1172 0 1 1105
box -2 -3 18 103
use NAND2X1  NAND2X1_59
timestamp 1626400951
transform 1 0 1172 0 1 1105
box -2 -3 26 103
use INVX1  INVX1_122
timestamp 1626400951
transform -1 0 1212 0 1 1105
box -2 -3 18 103
use BUFX2  BUFX2_36
timestamp 1626400951
transform -1 0 1236 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_208
timestamp 1626400951
transform 1 0 1236 0 1 1105
box -2 -3 26 103
use INVX1  INVX1_37
timestamp 1626400951
transform 1 0 1260 0 1 1105
box -2 -3 18 103
use NAND3X1  NAND3X1_18
timestamp 1626400951
transform 1 0 1276 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_38
timestamp 1626400951
transform -1 0 1324 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_27
timestamp 1626400951
transform -1 0 1356 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_28
timestamp 1626400951
transform 1 0 1356 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_29
timestamp 1626400951
transform -1 0 1420 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_29
timestamp 1626400951
transform -1 0 1452 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_39
timestamp 1626400951
transform -1 0 1468 0 1 1105
box -2 -3 18 103
use AOI21X1  AOI21X1_27
timestamp 1626400951
transform -1 0 1500 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_9
timestamp 1626400951
transform 1 0 1500 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_26
timestamp 1626400951
transform 1 0 1524 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_45
timestamp 1626400951
transform -1 0 1588 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_2_0
timestamp 1626400951
transform 1 0 1588 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_2_1
timestamp 1626400951
transform 1 0 1596 0 1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_109
timestamp 1626400951
transform 1 0 1604 0 1 1105
box -2 -3 98 103
use INVX2  INVX2_13
timestamp 1626400951
transform 1 0 1700 0 1 1105
box -2 -3 18 103
use NOR3X1  NOR3X1_4
timestamp 1626400951
transform 1 0 1716 0 1 1105
box -2 -3 66 103
use AND2X2  AND2X2_25
timestamp 1626400951
transform -1 0 1812 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_128
timestamp 1626400951
transform 1 0 1812 0 1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_127
timestamp 1626400951
transform 1 0 1908 0 1 1105
box -2 -3 98 103
use INVX8  INVX8_3
timestamp 1626400951
transform 1 0 2004 0 1 1105
box -2 -3 42 103
use NOR2X1  NOR2X1_183
timestamp 1626400951
transform -1 0 2068 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_134
timestamp 1626400951
transform -1 0 2092 0 1 1105
box -2 -3 26 103
use INVX1  INVX1_180
timestamp 1626400951
transform 1 0 2092 0 1 1105
box -2 -3 18 103
use FILL  FILL_11_3_0
timestamp 1626400951
transform 1 0 2108 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_3_1
timestamp 1626400951
transform 1 0 2116 0 1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_118
timestamp 1626400951
transform 1 0 2124 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_150
timestamp 1626400951
transform 1 0 2156 0 1 1105
box -2 -3 18 103
use NOR2X1  NOR2X1_120
timestamp 1626400951
transform -1 0 2196 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_124
timestamp 1626400951
transform 1 0 2196 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_130
timestamp 1626400951
transform -1 0 2252 0 1 1105
box -2 -3 34 103
use AND2X2  AND2X2_15
timestamp 1626400951
transform 1 0 2252 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_84
timestamp 1626400951
transform 1 0 2284 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_154
timestamp 1626400951
transform -1 0 2332 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_159
timestamp 1626400951
transform 1 0 2332 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_85
timestamp 1626400951
transform 1 0 2356 0 1 1105
box -2 -3 26 103
use AND2X2  AND2X2_16
timestamp 1626400951
transform 1 0 2380 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_93
timestamp 1626400951
transform 1 0 2412 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_88
timestamp 1626400951
transform -1 0 2460 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_83
timestamp 1626400951
transform 1 0 2460 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_86
timestamp 1626400951
transform -1 0 2508 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_122
timestamp 1626400951
transform -1 0 2532 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_121
timestamp 1626400951
transform -1 0 2556 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_135
timestamp 1626400951
transform -1 0 2580 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_134
timestamp 1626400951
transform -1 0 2604 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_96
timestamp 1626400951
transform 1 0 2604 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_97
timestamp 1626400951
transform 1 0 2636 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_94
timestamp 1626400951
transform -1 0 2692 0 1 1105
box -2 -3 26 103
use FILL  FILL_12_1
timestamp 1626400951
transform 1 0 2692 0 1 1105
box -2 -3 10 103
use FILL  FILL_12_2
timestamp 1626400951
transform 1 0 2700 0 1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_47
timestamp 1626400951
transform 1 0 4 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_42
timestamp 1626400951
transform 1 0 36 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_65
timestamp 1626400951
transform -1 0 84 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_49
timestamp 1626400951
transform 1 0 84 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_47
timestamp 1626400951
transform 1 0 116 0 -1 1105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_9
timestamp 1626400951
transform -1 0 196 0 -1 1105
box -2 -3 58 103
use INVX1  INVX1_62
timestamp 1626400951
transform 1 0 196 0 -1 1105
box -2 -3 18 103
use NOR2X1  NOR2X1_43
timestamp 1626400951
transform 1 0 212 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_79
timestamp 1626400951
transform -1 0 332 0 -1 1105
box -2 -3 98 103
use INVX1  INVX1_116
timestamp 1626400951
transform 1 0 332 0 -1 1105
box -2 -3 18 103
use NOR2X1  NOR2X1_91
timestamp 1626400951
transform 1 0 348 0 -1 1105
box -2 -3 26 103
use NOR3X1  NOR3X1_3
timestamp 1626400951
transform -1 0 436 0 -1 1105
box -2 -3 66 103
use INVX1  INVX1_107
timestamp 1626400951
transform -1 0 452 0 -1 1105
box -2 -3 18 103
use NOR2X1  NOR2X1_80
timestamp 1626400951
transform 1 0 452 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_68
timestamp 1626400951
transform 1 0 476 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_82
timestamp 1626400951
transform -1 0 532 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_69
timestamp 1626400951
transform -1 0 564 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_0_0
timestamp 1626400951
transform -1 0 572 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_0_1
timestamp 1626400951
transform -1 0 580 0 -1 1105
box -2 -3 10 103
use AOI21X1  AOI21X1_53
timestamp 1626400951
transform -1 0 612 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_54
timestamp 1626400951
transform 1 0 612 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_30
timestamp 1626400951
transform -1 0 676 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_57
timestamp 1626400951
transform -1 0 772 0 -1 1105
box -2 -3 98 103
use AOI21X1  AOI21X1_14
timestamp 1626400951
transform -1 0 804 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_14
timestamp 1626400951
transform -1 0 836 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_15
timestamp 1626400951
transform -1 0 868 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_15
timestamp 1626400951
transform -1 0 900 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_61
timestamp 1626400951
transform 1 0 900 0 -1 1105
box -2 -3 26 103
use INVX1  INVX1_127
timestamp 1626400951
transform -1 0 940 0 -1 1105
box -2 -3 18 103
use NAND3X1  NAND3X1_32
timestamp 1626400951
transform -1 0 972 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_95
timestamp 1626400951
transform -1 0 996 0 -1 1105
box -2 -3 26 103
use OR2X2  OR2X2_16
timestamp 1626400951
transform 1 0 996 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_79
timestamp 1626400951
transform 1 0 1028 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_31
timestamp 1626400951
transform -1 0 1092 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_1_0
timestamp 1626400951
transform -1 0 1100 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_1_1
timestamp 1626400951
transform -1 0 1108 0 -1 1105
box -2 -3 10 103
use AOI22X1  AOI22X1_17
timestamp 1626400951
transform -1 0 1148 0 -1 1105
box -2 -3 42 103
use AOI21X1  AOI21X1_62
timestamp 1626400951
transform 1 0 1148 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_108
timestamp 1626400951
transform -1 0 1204 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_78
timestamp 1626400951
transform -1 0 1236 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_10
timestamp 1626400951
transform -1 0 1332 0 -1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_9
timestamp 1626400951
transform -1 0 1428 0 -1 1105
box -2 -3 98 103
use NOR2X1  NOR2X1_31
timestamp 1626400951
transform -1 0 1452 0 -1 1105
box -2 -3 26 103
use NOR3X1  NOR3X1_5
timestamp 1626400951
transform -1 0 1516 0 -1 1105
box -2 -3 66 103
use AND2X2  AND2X2_26
timestamp 1626400951
transform -1 0 1548 0 -1 1105
box -2 -3 34 103
use OR2X2  OR2X2_20
timestamp 1626400951
transform 1 0 1548 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_84
timestamp 1626400951
transform 1 0 1580 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_2_0
timestamp 1626400951
transform -1 0 1620 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_2_1
timestamp 1626400951
transform -1 0 1628 0 -1 1105
box -2 -3 10 103
use INVX1  INVX1_186
timestamp 1626400951
transform -1 0 1644 0 -1 1105
box -2 -3 18 103
use NAND3X1  NAND3X1_39
timestamp 1626400951
transform -1 0 1676 0 -1 1105
box -2 -3 34 103
use AND2X2  AND2X2_24
timestamp 1626400951
transform 1 0 1676 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_38
timestamp 1626400951
transform 1 0 1708 0 -1 1105
box -2 -3 34 103
use INVX2  INVX2_15
timestamp 1626400951
transform 1 0 1740 0 -1 1105
box -2 -3 18 103
use NAND3X1  NAND3X1_44
timestamp 1626400951
transform -1 0 1788 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_96
timestamp 1626400951
transform -1 0 1820 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_143
timestamp 1626400951
transform 1 0 1820 0 -1 1105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_23
timestamp 1626400951
transform -1 0 1908 0 -1 1105
box -2 -3 58 103
use AOI21X1  AOI21X1_97
timestamp 1626400951
transform -1 0 1940 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_144
timestamp 1626400951
transform 1 0 1940 0 -1 1105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_22
timestamp 1626400951
transform -1 0 2028 0 -1 1105
box -2 -3 58 103
use NAND2X1  NAND2X1_106
timestamp 1626400951
transform 1 0 2028 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_117
timestamp 1626400951
transform 1 0 2052 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_74
timestamp 1626400951
transform -1 0 2116 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_3_0
timestamp 1626400951
transform -1 0 2124 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_3_1
timestamp 1626400951
transform -1 0 2132 0 -1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_116
timestamp 1626400951
transform -1 0 2164 0 -1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_2
timestamp 1626400951
transform 1 0 2164 0 -1 1105
box -2 -3 50 103
use INVX1  INVX1_172
timestamp 1626400951
transform -1 0 2228 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_129
timestamp 1626400951
transform -1 0 2260 0 -1 1105
box -2 -3 34 103
use AND2X2  AND2X2_23
timestamp 1626400951
transform 1 0 2260 0 -1 1105
box -2 -3 34 103
use BUFX4  BUFX4_49
timestamp 1626400951
transform -1 0 2324 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_153
timestamp 1626400951
transform 1 0 2324 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_155
timestamp 1626400951
transform 1 0 2348 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_123
timestamp 1626400951
transform -1 0 2396 0 -1 1105
box -2 -3 26 103
use INVX1  INVX1_153
timestamp 1626400951
transform 1 0 2396 0 -1 1105
box -2 -3 18 103
use XOR2X1  XOR2X1_13
timestamp 1626400951
transform 1 0 2412 0 -1 1105
box -2 -3 58 103
use NOR2X1  NOR2X1_133
timestamp 1626400951
transform -1 0 2492 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_67
timestamp 1626400951
transform -1 0 2524 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_93
timestamp 1626400951
transform 1 0 2524 0 -1 1105
box -2 -3 34 103
use XOR2X1  XOR2X1_14
timestamp 1626400951
transform 1 0 2556 0 -1 1105
box -2 -3 58 103
use OAI21X1  OAI21X1_94
timestamp 1626400951
transform -1 0 2644 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_95
timestamp 1626400951
transform -1 0 2676 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_162
timestamp 1626400951
transform -1 0 2692 0 -1 1105
box -2 -3 18 103
use FILL  FILL_11_1
timestamp 1626400951
transform -1 0 2700 0 -1 1105
box -2 -3 10 103
use FILL  FILL_11_2
timestamp 1626400951
transform -1 0 2708 0 -1 1105
box -2 -3 10 103
use INVX1  INVX1_82
timestamp 1626400951
transform 1 0 4 0 1 905
box -2 -3 18 103
use OAI22X1  OAI22X1_3
timestamp 1626400951
transform 1 0 20 0 1 905
box -2 -3 42 103
use INVX1  INVX1_83
timestamp 1626400951
transform 1 0 60 0 1 905
box -2 -3 18 103
use AOI22X1  AOI22X1_15
timestamp 1626400951
transform -1 0 116 0 1 905
box -2 -3 42 103
use NAND2X1  NAND2X1_45
timestamp 1626400951
transform -1 0 140 0 1 905
box -2 -3 26 103
use AND2X2  AND2X2_8
timestamp 1626400951
transform 1 0 140 0 1 905
box -2 -3 34 103
use XOR2X1  XOR2X1_5
timestamp 1626400951
transform -1 0 228 0 1 905
box -2 -3 58 103
use OAI21X1  OAI21X1_35
timestamp 1626400951
transform 1 0 228 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_22
timestamp 1626400951
transform -1 0 284 0 1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_35
timestamp 1626400951
transform 1 0 284 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_42
timestamp 1626400951
transform 1 0 316 0 1 905
box -2 -3 26 103
use INVX1  INVX1_61
timestamp 1626400951
transform -1 0 356 0 1 905
box -2 -3 18 103
use INVX1  INVX1_143
timestamp 1626400951
transform 1 0 356 0 1 905
box -2 -3 18 103
use XNOR2X1  XNOR2X1_13
timestamp 1626400951
transform -1 0 428 0 1 905
box -2 -3 58 103
use NOR2X1  NOR2X1_105
timestamp 1626400951
transform -1 0 452 0 1 905
box -2 -3 26 103
use INVX1  INVX1_106
timestamp 1626400951
transform -1 0 468 0 1 905
box -2 -3 18 103
use AOI21X1  AOI21X1_61
timestamp 1626400951
transform -1 0 500 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_81
timestamp 1626400951
transform 1 0 500 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_67
timestamp 1626400951
transform -1 0 556 0 1 905
box -2 -3 34 103
use INVX1  INVX1_105
timestamp 1626400951
transform 1 0 556 0 1 905
box -2 -3 18 103
use FILL  FILL_9_0_0
timestamp 1626400951
transform -1 0 580 0 1 905
box -2 -3 10 103
use FILL  FILL_9_0_1
timestamp 1626400951
transform -1 0 588 0 1 905
box -2 -3 10 103
use AOI21X1  AOI21X1_12
timestamp 1626400951
transform -1 0 620 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_95
timestamp 1626400951
transform 1 0 620 0 1 905
box -2 -3 98 103
use NAND3X1  NAND3X1_12
timestamp 1626400951
transform 1 0 716 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_83
timestamp 1626400951
transform 1 0 748 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_56
timestamp 1626400951
transform -1 0 796 0 1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_14
timestamp 1626400951
transform -1 0 828 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_15
timestamp 1626400951
transform -1 0 860 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_14
timestamp 1626400951
transform -1 0 892 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_6
timestamp 1626400951
transform -1 0 924 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_29
timestamp 1626400951
transform -1 0 956 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_70
timestamp 1626400951
transform -1 0 988 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_55
timestamp 1626400951
transform -1 0 1020 0 1 905
box -2 -3 34 103
use INVX1  INVX1_108
timestamp 1626400951
transform -1 0 1036 0 1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_99
timestamp 1626400951
transform 1 0 1036 0 1 905
box -2 -3 98 103
use FILL  FILL_9_1_0
timestamp 1626400951
transform 1 0 1132 0 1 905
box -2 -3 10 103
use FILL  FILL_9_1_1
timestamp 1626400951
transform 1 0 1140 0 1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_59
timestamp 1626400951
transform 1 0 1148 0 1 905
box -2 -3 98 103
use INVX2  INVX2_8
timestamp 1626400951
transform -1 0 1260 0 1 905
box -2 -3 18 103
use INVX1  INVX1_119
timestamp 1626400951
transform 1 0 1260 0 1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_81
timestamp 1626400951
transform -1 0 1372 0 1 905
box -2 -3 98 103
use AOI21X1  AOI21X1_30
timestamp 1626400951
transform 1 0 1372 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_30
timestamp 1626400951
transform -1 0 1436 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_18
timestamp 1626400951
transform 1 0 1436 0 1 905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_7
timestamp 1626400951
transform 1 0 1468 0 1 905
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_108
timestamp 1626400951
transform 1 0 1540 0 1 905
box -2 -3 98 103
use FILL  FILL_9_2_0
timestamp 1626400951
transform -1 0 1644 0 1 905
box -2 -3 10 103
use FILL  FILL_9_2_1
timestamp 1626400951
transform -1 0 1652 0 1 905
box -2 -3 10 103
use AOI21X1  AOI21X1_83
timestamp 1626400951
transform -1 0 1684 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_113
timestamp 1626400951
transform -1 0 1708 0 1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_81
timestamp 1626400951
transform 1 0 1708 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_124
timestamp 1626400951
transform 1 0 1740 0 1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_137
timestamp 1626400951
transform 1 0 1836 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_147
timestamp 1626400951
transform 1 0 1860 0 1 905
box -2 -3 34 103
use INVX1  INVX1_200
timestamp 1626400951
transform -1 0 1908 0 1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_129
timestamp 1626400951
transform 1 0 1908 0 1 905
box -2 -3 98 103
use AOI21X1  AOI21X1_95
timestamp 1626400951
transform -1 0 2036 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_142
timestamp 1626400951
transform -1 0 2068 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_102
timestamp 1626400951
transform 1 0 2068 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_181
timestamp 1626400951
transform -1 0 2116 0 1 905
box -2 -3 26 103
use FILL  FILL_9_3_0
timestamp 1626400951
transform -1 0 2124 0 1 905
box -2 -3 10 103
use FILL  FILL_9_3_1
timestamp 1626400951
transform -1 0 2132 0 1 905
box -2 -3 10 103
use NAND2X1  NAND2X1_132
timestamp 1626400951
transform -1 0 2156 0 1 905
box -2 -3 26 103
use XOR2X1  XOR2X1_11
timestamp 1626400951
transform 1 0 2156 0 1 905
box -2 -3 58 103
use NOR2X1  NOR2X1_147
timestamp 1626400951
transform -1 0 2236 0 1 905
box -2 -3 26 103
use BUFX4  BUFX4_36
timestamp 1626400951
transform 1 0 2236 0 1 905
box -2 -3 34 103
use INVX1  INVX1_176
timestamp 1626400951
transform -1 0 2284 0 1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_103
timestamp 1626400951
transform -1 0 2308 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_89
timestamp 1626400951
transform -1 0 2332 0 1 905
box -2 -3 26 103
use BUFX4  BUFX4_50
timestamp 1626400951
transform 1 0 2332 0 1 905
box -2 -3 34 103
use OR2X2  OR2X2_19
timestamp 1626400951
transform -1 0 2396 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_91
timestamp 1626400951
transform -1 0 2420 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_156
timestamp 1626400951
transform 1 0 2420 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_130
timestamp 1626400951
transform -1 0 2468 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_125
timestamp 1626400951
transform 1 0 2468 0 1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_1
timestamp 1626400951
transform 1 0 2492 0 1 905
box -2 -3 50 103
use NOR2X1  NOR2X1_188
timestamp 1626400951
transform 1 0 2540 0 1 905
box -2 -3 26 103
use XOR2X1  XOR2X1_16
timestamp 1626400951
transform 1 0 2564 0 1 905
box -2 -3 58 103
use XNOR2X1  XNOR2X1_20
timestamp 1626400951
transform -1 0 2676 0 1 905
box -2 -3 58 103
use NOR2X1  NOR2X1_131
timestamp 1626400951
transform -1 0 2700 0 1 905
box -2 -3 26 103
use FILL  FILL_10_1
timestamp 1626400951
transform 1 0 2700 0 1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_46
timestamp 1626400951
transform -1 0 36 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_80
timestamp 1626400951
transform -1 0 52 0 -1 905
box -2 -3 18 103
use AOI22X1  AOI22X1_14
timestamp 1626400951
transform 1 0 52 0 -1 905
box -2 -3 42 103
use INVX1  INVX1_81
timestamp 1626400951
transform -1 0 108 0 -1 905
box -2 -3 18 103
use XOR2X1  XOR2X1_4
timestamp 1626400951
transform 1 0 108 0 -1 905
box -2 -3 58 103
use NAND2X1  NAND2X1_37
timestamp 1626400951
transform -1 0 188 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_53
timestamp 1626400951
transform 1 0 188 0 -1 905
box -2 -3 26 103
use XNOR2X1  XNOR2X1_3
timestamp 1626400951
transform 1 0 212 0 -1 905
box -2 -3 58 103
use XNOR2X1  XNOR2X1_2
timestamp 1626400951
transform -1 0 324 0 -1 905
box -2 -3 58 103
use XOR2X1  XOR2X1_2
timestamp 1626400951
transform 1 0 324 0 -1 905
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_55
timestamp 1626400951
transform -1 0 476 0 -1 905
box -2 -3 98 103
use NOR2X1  NOR2X1_106
timestamp 1626400951
transform -1 0 500 0 -1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_33
timestamp 1626400951
transform -1 0 532 0 -1 905
box -2 -3 34 103
use OR2X2  OR2X2_15
timestamp 1626400951
transform -1 0 564 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_62
timestamp 1626400951
transform -1 0 588 0 -1 905
box -2 -3 26 103
use FILL  FILL_8_0_0
timestamp 1626400951
transform -1 0 596 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_0_1
timestamp 1626400951
transform -1 0 604 0 -1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_12
timestamp 1626400951
transform -1 0 636 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_11
timestamp 1626400951
transform -1 0 668 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_94
timestamp 1626400951
transform -1 0 764 0 -1 905
box -2 -3 98 103
use NOR2X1  NOR2X1_79
timestamp 1626400951
transform 1 0 764 0 -1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_98
timestamp 1626400951
transform 1 0 788 0 -1 905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_97
timestamp 1626400951
transform -1 0 980 0 -1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_16
timestamp 1626400951
transform 1 0 980 0 -1 905
box -2 -3 34 103
use BUFX4  BUFX4_1
timestamp 1626400951
transform -1 0 1044 0 -1 905
box -2 -3 34 103
use INVX8  INVX8_1
timestamp 1626400951
transform -1 0 1084 0 -1 905
box -2 -3 42 103
use FILL  FILL_8_1_0
timestamp 1626400951
transform -1 0 1092 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_1_1
timestamp 1626400951
transform -1 0 1100 0 -1 905
box -2 -3 10 103
use AOI21X1  AOI21X1_16
timestamp 1626400951
transform -1 0 1132 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_16
timestamp 1626400951
transform 1 0 1132 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_121
timestamp 1626400951
transform 1 0 1164 0 -1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_58
timestamp 1626400951
transform -1 0 1204 0 -1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_83
timestamp 1626400951
transform -1 0 1300 0 -1 905
box -2 -3 98 103
use NOR2X1  NOR2X1_94
timestamp 1626400951
transform 1 0 1300 0 -1 905
box -2 -3 26 103
use INVX1  INVX1_117
timestamp 1626400951
transform 1 0 1324 0 -1 905
box -2 -3 18 103
use NOR2X1  NOR2X1_92
timestamp 1626400951
transform 1 0 1340 0 -1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_2
timestamp 1626400951
transform 1 0 1364 0 -1 905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_113
timestamp 1626400951
transform -1 0 1556 0 -1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_110
timestamp 1626400951
transform 1 0 1556 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_132
timestamp 1626400951
transform -1 0 1612 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_2_0
timestamp 1626400951
transform -1 0 1620 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_2_1
timestamp 1626400951
transform -1 0 1628 0 -1 905
box -2 -3 10 103
use AOI21X1  AOI21X1_85
timestamp 1626400951
transform -1 0 1660 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_185
timestamp 1626400951
transform 1 0 1660 0 -1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_112
timestamp 1626400951
transform 1 0 1676 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_111
timestamp 1626400951
transform -1 0 1724 0 -1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_106
timestamp 1626400951
transform 1 0 1724 0 -1 905
box -2 -3 98 103
use INVX1  INVX1_187
timestamp 1626400951
transform -1 0 1836 0 -1 905
box -2 -3 18 103
use NOR2X1  NOR2X1_182
timestamp 1626400951
transform 1 0 1836 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_133
timestamp 1626400951
transform -1 0 1884 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_100
timestamp 1626400951
transform -1 0 1916 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_187
timestamp 1626400951
transform -1 0 1940 0 -1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_43
timestamp 1626400951
transform -1 0 1972 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_157
timestamp 1626400951
transform 1 0 1972 0 -1 905
box -2 -3 18 103
use NOR2X1  NOR2X1_186
timestamp 1626400951
transform -1 0 2012 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_148
timestamp 1626400951
transform 1 0 2012 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_136
timestamp 1626400951
transform -1 0 2068 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_157
timestamp 1626400951
transform 1 0 2068 0 -1 905
box -2 -3 26 103
use INVX1  INVX1_174
timestamp 1626400951
transform 1 0 2092 0 -1 905
box -2 -3 18 103
use FILL  FILL_8_3_0
timestamp 1626400951
transform 1 0 2108 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_3_1
timestamp 1626400951
transform 1 0 2116 0 -1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_108
timestamp 1626400951
transform 1 0 2124 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_111
timestamp 1626400951
transform -1 0 2188 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_73
timestamp 1626400951
transform -1 0 2220 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_109
timestamp 1626400951
transform 1 0 2220 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_110
timestamp 1626400951
transform 1 0 2252 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_177
timestamp 1626400951
transform -1 0 2300 0 -1 905
box -2 -3 18 103
use INVX1  INVX1_173
timestamp 1626400951
transform -1 0 2316 0 -1 905
box -2 -3 18 103
use XOR2X1  XOR2X1_12
timestamp 1626400951
transform 1 0 2316 0 -1 905
box -2 -3 58 103
use INVX1  INVX1_155
timestamp 1626400951
transform 1 0 2372 0 -1 905
box -2 -3 18 103
use INVX4  INVX4_1
timestamp 1626400951
transform -1 0 2412 0 -1 905
box -2 -3 26 103
use INVX1  INVX1_158
timestamp 1626400951
transform 1 0 2412 0 -1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_89
timestamp 1626400951
transform 1 0 2428 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_90
timestamp 1626400951
transform 1 0 2460 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_132
timestamp 1626400951
transform -1 0 2516 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_92
timestamp 1626400951
transform 1 0 2516 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_91
timestamp 1626400951
transform 1 0 2548 0 -1 905
box -2 -3 34 103
use XOR2X1  XOR2X1_15
timestamp 1626400951
transform 1 0 2580 0 -1 905
box -2 -3 58 103
use XNOR2X1  XNOR2X1_21
timestamp 1626400951
transform -1 0 2692 0 -1 905
box -2 -3 58 103
use FILL  FILL_9_1
timestamp 1626400951
transform -1 0 2700 0 -1 905
box -2 -3 10 103
use FILL  FILL_9_2
timestamp 1626400951
transform -1 0 2708 0 -1 905
box -2 -3 10 103
use INVX1  INVX1_55
timestamp 1626400951
transform 1 0 4 0 1 705
box -2 -3 18 103
use AOI22X1  AOI22X1_9
timestamp 1626400951
transform -1 0 60 0 1 705
box -2 -3 42 103
use OAI22X1  OAI22X1_1
timestamp 1626400951
transform -1 0 100 0 1 705
box -2 -3 42 103
use INVX1  INVX1_54
timestamp 1626400951
transform -1 0 116 0 1 705
box -2 -3 18 103
use INVX1  INVX1_53
timestamp 1626400951
transform 1 0 116 0 1 705
box -2 -3 18 103
use AOI22X1  AOI22X1_8
timestamp 1626400951
transform -1 0 172 0 1 705
box -2 -3 42 103
use OAI21X1  OAI21X1_33
timestamp 1626400951
transform -1 0 204 0 1 705
box -2 -3 34 103
use INVX1  INVX1_52
timestamp 1626400951
transform -1 0 220 0 1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_25
timestamp 1626400951
transform 1 0 220 0 1 705
box -2 -3 26 103
use AND2X2  AND2X2_5
timestamp 1626400951
transform 1 0 244 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_34
timestamp 1626400951
transform 1 0 276 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_17
timestamp 1626400951
transform -1 0 332 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_36
timestamp 1626400951
transform 1 0 332 0 1 705
box -2 -3 26 103
use XOR2X1  XOR2X1_1
timestamp 1626400951
transform -1 0 412 0 1 705
box -2 -3 58 103
use INVX1  INVX1_128
timestamp 1626400951
transform 1 0 412 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_76
timestamp 1626400951
transform -1 0 460 0 1 705
box -2 -3 34 103
use AOI22X1  AOI22X1_19
timestamp 1626400951
transform 1 0 460 0 1 705
box -2 -3 42 103
use INVX1  INVX1_129
timestamp 1626400951
transform -1 0 516 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_77
timestamp 1626400951
transform 1 0 516 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_29
timestamp 1626400951
transform 1 0 548 0 1 705
box -2 -3 34 103
use FILL  FILL_7_0_0
timestamp 1626400951
transform -1 0 588 0 1 705
box -2 -3 10 103
use FILL  FILL_7_0_1
timestamp 1626400951
transform -1 0 596 0 1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_54
timestamp 1626400951
transform -1 0 692 0 1 705
box -2 -3 98 103
use AOI21X1  AOI21X1_11
timestamp 1626400951
transform -1 0 724 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_11
timestamp 1626400951
transform -1 0 756 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_66
timestamp 1626400951
transform -1 0 788 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_52
timestamp 1626400951
transform -1 0 884 0 1 705
box -2 -3 98 103
use INVX1  INVX1_104
timestamp 1626400951
transform -1 0 900 0 1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_55
timestamp 1626400951
transform -1 0 924 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_65
timestamp 1626400951
transform 1 0 924 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_78
timestamp 1626400951
transform -1 0 980 0 1 705
box -2 -3 26 103
use BUFX4  BUFX4_26
timestamp 1626400951
transform -1 0 1012 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_63
timestamp 1626400951
transform 1 0 1012 0 1 705
box -2 -3 34 103
use FILL  FILL_7_1_0
timestamp 1626400951
transform 1 0 1044 0 1 705
box -2 -3 10 103
use FILL  FILL_7_1_1
timestamp 1626400951
transform 1 0 1052 0 1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_93
timestamp 1626400951
transform 1 0 1060 0 1 705
box -2 -3 98 103
use BUFX4  BUFX4_13
timestamp 1626400951
transform 1 0 1156 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_53
timestamp 1626400951
transform 1 0 1188 0 1 705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_44
timestamp 1626400951
transform -1 0 1380 0 1 705
box -2 -3 98 103
use BUFX4  BUFX4_4
timestamp 1626400951
transform 1 0 1380 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_19
timestamp 1626400951
transform 1 0 1412 0 1 705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_5
timestamp 1626400951
transform -1 0 1516 0 1 705
box -2 -3 74 103
use CLKBUF1  CLKBUF1_9
timestamp 1626400951
transform -1 0 1588 0 1 705
box -2 -3 74 103
use FILL  FILL_7_2_0
timestamp 1626400951
transform 1 0 1588 0 1 705
box -2 -3 10 103
use FILL  FILL_7_2_1
timestamp 1626400951
transform 1 0 1596 0 1 705
box -2 -3 10 103
use AND2X2  AND2X2_30
timestamp 1626400951
transform 1 0 1604 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_119
timestamp 1626400951
transform 1 0 1636 0 1 705
box -2 -3 26 103
use INVX1  INVX1_193
timestamp 1626400951
transform -1 0 1676 0 1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_114
timestamp 1626400951
transform 1 0 1676 0 1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_115
timestamp 1626400951
transform -1 0 1796 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_82
timestamp 1626400951
transform -1 0 1828 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_40
timestamp 1626400951
transform -1 0 1860 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_172
timestamp 1626400951
transform -1 0 1884 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_114
timestamp 1626400951
transform -1 0 1908 0 1 705
box -2 -3 26 103
use OR2X2  OR2X2_23
timestamp 1626400951
transform 1 0 1908 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_133
timestamp 1626400951
transform -1 0 1972 0 1 705
box -2 -3 34 103
use OR2X2  OR2X2_22
timestamp 1626400951
transform -1 0 2004 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_189
timestamp 1626400951
transform -1 0 2028 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_138
timestamp 1626400951
transform -1 0 2052 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_101
timestamp 1626400951
transform -1 0 2084 0 1 705
box -2 -3 34 103
use FILL  FILL_7_3_0
timestamp 1626400951
transform 1 0 2084 0 1 705
box -2 -3 10 103
use FILL  FILL_7_3_1
timestamp 1626400951
transform 1 0 2092 0 1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_123
timestamp 1626400951
transform 1 0 2100 0 1 705
box -2 -3 98 103
use INVX1  INVX1_201
timestamp 1626400951
transform -1 0 2212 0 1 705
box -2 -3 18 103
use INVX1  INVX1_175
timestamp 1626400951
transform 1 0 2212 0 1 705
box -2 -3 18 103
use INVX1  INVX1_170
timestamp 1626400951
transform -1 0 2244 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_113
timestamp 1626400951
transform 1 0 2244 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_37
timestamp 1626400951
transform 1 0 2276 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_115
timestamp 1626400951
transform 1 0 2308 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_114
timestamp 1626400951
transform -1 0 2372 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_158
timestamp 1626400951
transform 1 0 2372 0 1 705
box -2 -3 26 103
use INVX1  INVX1_179
timestamp 1626400951
transform -1 0 2412 0 1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_105
timestamp 1626400951
transform 1 0 2412 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_190
timestamp 1626400951
transform 1 0 2436 0 1 705
box -2 -3 26 103
use XOR2X1  XOR2X1_17
timestamp 1626400951
transform 1 0 2460 0 1 705
box -2 -3 58 103
use NAND3X1  NAND3X1_35
timestamp 1626400951
transform -1 0 2548 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_92
timestamp 1626400951
transform -1 0 2572 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_87
timestamp 1626400951
transform -1 0 2604 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_86
timestamp 1626400951
transform -1 0 2636 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_128
timestamp 1626400951
transform 1 0 2636 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_87
timestamp 1626400951
transform 1 0 2660 0 1 705
box -2 -3 26 103
use INVX1  INVX1_156
timestamp 1626400951
transform -1 0 2700 0 1 705
box -2 -3 18 103
use FILL  FILL_8_1
timestamp 1626400951
transform 1 0 2700 0 1 705
box -2 -3 10 103
use INVX1  INVX1_87
timestamp 1626400951
transform 1 0 4 0 -1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_41
timestamp 1626400951
transform 1 0 20 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_57
timestamp 1626400951
transform -1 0 68 0 -1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_42
timestamp 1626400951
transform -1 0 100 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_55
timestamp 1626400951
transform -1 0 132 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_66
timestamp 1626400951
transform -1 0 156 0 -1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_43
timestamp 1626400951
transform 1 0 156 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_46
timestamp 1626400951
transform -1 0 212 0 -1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_34
timestamp 1626400951
transform 1 0 212 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_48
timestamp 1626400951
transform 1 0 244 0 -1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_40
timestamp 1626400951
transform -1 0 300 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_27
timestamp 1626400951
transform 1 0 300 0 -1 705
box -2 -3 26 103
use INVX1  INVX1_131
timestamp 1626400951
transform -1 0 340 0 -1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_64
timestamp 1626400951
transform -1 0 364 0 -1 705
box -2 -3 26 103
use OAI22X1  OAI22X1_6
timestamp 1626400951
transform -1 0 404 0 -1 705
box -2 -3 42 103
use NAND3X1  NAND3X1_34
timestamp 1626400951
transform -1 0 436 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_63
timestamp 1626400951
transform -1 0 460 0 -1 705
box -2 -3 26 103
use INVX1  INVX1_130
timestamp 1626400951
transform -1 0 476 0 -1 705
box -2 -3 18 103
use NOR2X1  NOR2X1_96
timestamp 1626400951
transform 1 0 476 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_91
timestamp 1626400951
transform 1 0 500 0 -1 705
box -2 -3 98 103
use FILL  FILL_6_0_0
timestamp 1626400951
transform 1 0 596 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_0_1
timestamp 1626400951
transform 1 0 604 0 -1 705
box -2 -3 10 103
use NOR2X1  NOR2X1_76
timestamp 1626400951
transform 1 0 612 0 -1 705
box -2 -3 26 103
use NAND3X1  NAND3X1_8
timestamp 1626400951
transform 1 0 636 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_64
timestamp 1626400951
transform 1 0 668 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_77
timestamp 1626400951
transform -1 0 724 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_92
timestamp 1626400951
transform 1 0 724 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_9
timestamp 1626400951
transform -1 0 852 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_9
timestamp 1626400951
transform -1 0 884 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_9
timestamp 1626400951
transform 1 0 884 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_16
timestamp 1626400951
transform -1 0 948 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_25
timestamp 1626400951
transform -1 0 980 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_8
timestamp 1626400951
transform -1 0 1012 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_3
timestamp 1626400951
transform -1 0 1044 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_15
timestamp 1626400951
transform -1 0 1076 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_1_0
timestamp 1626400951
transform 1 0 1076 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_1_1
timestamp 1626400951
transform 1 0 1084 0 -1 705
box -2 -3 10 103
use BUFX4  BUFX4_2
timestamp 1626400951
transform 1 0 1092 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_7
timestamp 1626400951
transform 1 0 1124 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_10
timestamp 1626400951
transform 1 0 1156 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_10
timestamp 1626400951
transform -1 0 1220 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_4
timestamp 1626400951
transform -1 0 1252 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_10
timestamp 1626400951
transform -1 0 1284 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_27
timestamp 1626400951
transform 1 0 1284 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_23
timestamp 1626400951
transform 1 0 1316 0 -1 705
box -2 -3 34 103
use INVX8  INVX8_4
timestamp 1626400951
transform 1 0 1348 0 -1 705
box -2 -3 42 103
use OAI21X1  OAI21X1_1
timestamp 1626400951
transform -1 0 1420 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_1
timestamp 1626400951
transform 1 0 1420 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_2
timestamp 1626400951
transform 1 0 1452 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_2
timestamp 1626400951
transform 1 0 1484 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_45
timestamp 1626400951
transform -1 0 1612 0 -1 705
box -2 -3 98 103
use FILL  FILL_6_2_0
timestamp 1626400951
transform 1 0 1612 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_2_1
timestamp 1626400951
transform 1 0 1620 0 -1 705
box -2 -3 10 103
use NAND2X1  NAND2X1_120
timestamp 1626400951
transform 1 0 1628 0 -1 705
box -2 -3 26 103
use INVX1  INVX1_194
timestamp 1626400951
transform -1 0 1668 0 -1 705
box -2 -3 18 103
use BUFX4  BUFX4_46
timestamp 1626400951
transform -1 0 1700 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_41
timestamp 1626400951
transform 1 0 1700 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_190
timestamp 1626400951
transform -1 0 1748 0 -1 705
box -2 -3 18 103
use INVX1  INVX1_188
timestamp 1626400951
transform 1 0 1748 0 -1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_116
timestamp 1626400951
transform -1 0 1788 0 -1 705
box -2 -3 26 103
use MUX2X1  MUX2X1_4
timestamp 1626400951
transform 1 0 1788 0 -1 705
box -2 -3 50 103
use NOR2X1  NOR2X1_173
timestamp 1626400951
transform 1 0 1836 0 -1 705
box -2 -3 26 103
use OR2X2  OR2X2_21
timestamp 1626400951
transform 1 0 1860 0 -1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_3
timestamp 1626400951
transform -1 0 1940 0 -1 705
box -2 -3 50 103
use XNOR2X1  XNOR2X1_25
timestamp 1626400951
transform -1 0 1996 0 -1 705
box -2 -3 58 103
use BUFX2  BUFX2_38
timestamp 1626400951
transform -1 0 2020 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_131
timestamp 1626400951
transform 1 0 2020 0 -1 705
box -2 -3 26 103
use INVX1  INVX1_197
timestamp 1626400951
transform -1 0 2060 0 -1 705
box -2 -3 18 103
use INVX4  INVX4_3
timestamp 1626400951
transform -1 0 2084 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_185
timestamp 1626400951
transform 1 0 2084 0 -1 705
box -2 -3 26 103
use FILL  FILL_6_3_0
timestamp 1626400951
transform -1 0 2116 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_3_1
timestamp 1626400951
transform -1 0 2124 0 -1 705
box -2 -3 10 103
use NOR2X1  NOR2X1_184
timestamp 1626400951
transform -1 0 2148 0 -1 705
box -2 -3 26 103
use NAND3X1  NAND3X1_47
timestamp 1626400951
transform -1 0 2180 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_135
timestamp 1626400951
transform 1 0 2180 0 -1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_99
timestamp 1626400951
transform -1 0 2236 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_146
timestamp 1626400951
transform 1 0 2236 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_104
timestamp 1626400951
transform 1 0 2268 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_107
timestamp 1626400951
transform -1 0 2324 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_178
timestamp 1626400951
transform 1 0 2324 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_112
timestamp 1626400951
transform -1 0 2372 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_145
timestamp 1626400951
transform 1 0 2372 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_98
timestamp 1626400951
transform 1 0 2404 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_199
timestamp 1626400951
transform 1 0 2436 0 -1 705
box -2 -3 18 103
use INVX1  INVX1_198
timestamp 1626400951
transform 1 0 2452 0 -1 705
box -2 -3 18 103
use NAND3X1  NAND3X1_46
timestamp 1626400951
transform 1 0 2468 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_127
timestamp 1626400951
transform -1 0 2524 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_88
timestamp 1626400951
transform 1 0 2524 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_159
timestamp 1626400951
transform -1 0 2572 0 -1 705
box -2 -3 18 103
use XNOR2X1  XNOR2X1_19
timestamp 1626400951
transform 1 0 2572 0 -1 705
box -2 -3 58 103
use BUFX4  BUFX4_35
timestamp 1626400951
transform -1 0 2660 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_34
timestamp 1626400951
transform 1 0 2660 0 -1 705
box -2 -3 34 103
use FILL  FILL_7_1
timestamp 1626400951
transform -1 0 2700 0 -1 705
box -2 -3 10 103
use FILL  FILL_7_2
timestamp 1626400951
transform -1 0 2708 0 -1 705
box -2 -3 10 103
use XNOR2X1  XNOR2X1_10
timestamp 1626400951
transform 1 0 4 0 1 505
box -2 -3 58 103
use INVX1  INVX1_88
timestamp 1626400951
transform 1 0 60 0 1 505
box -2 -3 18 103
use NOR2X1  NOR2X1_58
timestamp 1626400951
transform -1 0 100 0 1 505
box -2 -3 26 103
use INVX1  INVX1_93
timestamp 1626400951
transform 1 0 100 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_53
timestamp 1626400951
transform -1 0 148 0 1 505
box -2 -3 34 103
use INVX1  INVX1_95
timestamp 1626400951
transform 1 0 148 0 1 505
box -2 -3 18 103
use NOR2X1  NOR2X1_67
timestamp 1626400951
transform 1 0 164 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_48
timestamp 1626400951
transform -1 0 220 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_48
timestamp 1626400951
transform -1 0 244 0 1 505
box -2 -3 26 103
use XNOR2X1  XNOR2X1_12
timestamp 1626400951
transform 1 0 244 0 1 505
box -2 -3 58 103
use OAI21X1  OAI21X1_42
timestamp 1626400951
transform -1 0 332 0 1 505
box -2 -3 34 103
use INVX1  INVX1_68
timestamp 1626400951
transform 1 0 332 0 1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_29
timestamp 1626400951
transform -1 0 372 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_39
timestamp 1626400951
transform 1 0 372 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_50
timestamp 1626400951
transform -1 0 428 0 1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_76
timestamp 1626400951
transform -1 0 524 0 1 505
box -2 -3 98 103
use OR2X2  OR2X2_12
timestamp 1626400951
transform -1 0 556 0 1 505
box -2 -3 34 103
use FILL  FILL_5_0_0
timestamp 1626400951
transform -1 0 564 0 1 505
box -2 -3 10 103
use FILL  FILL_5_0_1
timestamp 1626400951
transform -1 0 572 0 1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_51
timestamp 1626400951
transform -1 0 668 0 1 505
box -2 -3 98 103
use AOI21X1  AOI21X1_8
timestamp 1626400951
transform -1 0 700 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_63
timestamp 1626400951
transform -1 0 732 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_8
timestamp 1626400951
transform -1 0 764 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_7
timestamp 1626400951
transform 1 0 764 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_7
timestamp 1626400951
transform -1 0 828 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_49
timestamp 1626400951
transform -1 0 924 0 1 505
box -2 -3 98 103
use BUFX4  BUFX4_28
timestamp 1626400951
transform -1 0 956 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_24
timestamp 1626400951
transform -1 0 988 0 1 505
box -2 -3 34 103
use AND2X2  AND2X2_11
timestamp 1626400951
transform 1 0 988 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_72
timestamp 1626400951
transform 1 0 1020 0 1 505
box -2 -3 26 103
use BUFX4  BUFX4_5
timestamp 1626400951
transform -1 0 1076 0 1 505
box -2 -3 34 103
use FILL  FILL_5_1_0
timestamp 1626400951
transform -1 0 1084 0 1 505
box -2 -3 10 103
use FILL  FILL_5_1_1
timestamp 1626400951
transform -1 0 1092 0 1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_47
timestamp 1626400951
transform -1 0 1188 0 1 505
box -2 -3 98 103
use AOI21X1  AOI21X1_4
timestamp 1626400951
transform -1 0 1220 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_4
timestamp 1626400951
transform 1 0 1220 0 1 505
box -2 -3 34 103
use INVX2  INVX2_6
timestamp 1626400951
transform 1 0 1252 0 1 505
box -2 -3 18 103
use INVX1  INVX1_98
timestamp 1626400951
transform 1 0 1268 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_58
timestamp 1626400951
transform 1 0 1284 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_50
timestamp 1626400951
transform 1 0 1316 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_85
timestamp 1626400951
transform 1 0 1348 0 1 505
box -2 -3 98 103
use NAND3X1  NAND3X1_49
timestamp 1626400951
transform -1 0 1476 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_2
timestamp 1626400951
transform 1 0 1476 0 1 505
box -2 -3 34 103
use BUFX2  BUFX2_40
timestamp 1626400951
transform -1 0 1532 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_31
timestamp 1626400951
transform 1 0 1532 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_31
timestamp 1626400951
transform 1 0 1564 0 1 505
box -2 -3 34 103
use FILL  FILL_5_2_0
timestamp 1626400951
transform 1 0 1596 0 1 505
box -2 -3 10 103
use FILL  FILL_5_2_1
timestamp 1626400951
transform 1 0 1604 0 1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_119
timestamp 1626400951
transform 1 0 1612 0 1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_118
timestamp 1626400951
transform 1 0 1708 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_87
timestamp 1626400951
transform -1 0 1764 0 1 505
box -2 -3 34 103
use INVX1  INVX1_192
timestamp 1626400951
transform 1 0 1764 0 1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_117
timestamp 1626400951
transform 1 0 1780 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_86
timestamp 1626400951
transform -1 0 1836 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_107
timestamp 1626400951
transform 1 0 1836 0 1 505
box -2 -3 98 103
use INVX1  INVX1_191
timestamp 1626400951
transform -1 0 1948 0 1 505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_104
timestamp 1626400951
transform -1 0 2044 0 1 505
box -2 -3 98 103
use AOI21X1  AOI21X1_88
timestamp 1626400951
transform -1 0 2076 0 1 505
box -2 -3 34 103
use FILL  FILL_5_3_0
timestamp 1626400951
transform 1 0 2076 0 1 505
box -2 -3 10 103
use FILL  FILL_5_3_1
timestamp 1626400951
transform 1 0 2084 0 1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_116
timestamp 1626400951
transform 1 0 2092 0 1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_125
timestamp 1626400951
transform 1 0 2188 0 1 505
box -2 -3 98 103
use NOR2X1  NOR2X1_126
timestamp 1626400951
transform -1 0 2308 0 1 505
box -2 -3 26 103
use AND2X2  AND2X2_14
timestamp 1626400951
transform 1 0 2308 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_126
timestamp 1626400951
transform -1 0 2436 0 1 505
box -2 -3 98 103
use INVX1  INVX1_202
timestamp 1626400951
transform 1 0 2436 0 1 505
box -2 -3 18 103
use AND2X2  AND2X2_31
timestamp 1626400951
transform 1 0 2452 0 1 505
box -2 -3 34 103
use NOR3X1  NOR3X1_6
timestamp 1626400951
transform 1 0 2484 0 1 505
box -2 -3 66 103
use NOR2X1  NOR2X1_203
timestamp 1626400951
transform -1 0 2572 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_102
timestamp 1626400951
transform -1 0 2604 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_149
timestamp 1626400951
transform 1 0 2604 0 1 505
box -2 -3 34 103
use INVX1  INVX1_203
timestamp 1626400951
transform 1 0 2636 0 1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_139
timestamp 1626400951
transform 1 0 2652 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_191
timestamp 1626400951
transform 1 0 2676 0 1 505
box -2 -3 26 103
use FILL  FILL_6_1
timestamp 1626400951
transform 1 0 2700 0 1 505
box -2 -3 10 103
use XOR2X1  XOR2X1_6
timestamp 1626400951
transform -1 0 60 0 -1 505
box -2 -3 58 103
use NAND2X1  NAND2X1_38
timestamp 1626400951
transform 1 0 60 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_41
timestamp 1626400951
transform -1 0 116 0 -1 505
box -2 -3 34 103
use INVX1  INVX1_84
timestamp 1626400951
transform -1 0 132 0 -1 505
box -2 -3 18 103
use NOR2X1  NOR2X1_54
timestamp 1626400951
transform -1 0 156 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_40
timestamp 1626400951
transform -1 0 180 0 -1 505
box -2 -3 26 103
use XNOR2X1  XNOR2X1_11
timestamp 1626400951
transform 1 0 180 0 -1 505
box -2 -3 58 103
use INVX1  INVX1_96
timestamp 1626400951
transform 1 0 236 0 -1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_49
timestamp 1626400951
transform -1 0 276 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_56
timestamp 1626400951
transform 1 0 276 0 -1 505
box -2 -3 26 103
use INVX1  INVX1_86
timestamp 1626400951
transform -1 0 316 0 -1 505
box -2 -3 18 103
use XNOR2X1  XNOR2X1_6
timestamp 1626400951
transform 1 0 316 0 -1 505
box -2 -3 58 103
use INVX1  INVX1_58
timestamp 1626400951
transform -1 0 388 0 -1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_28
timestamp 1626400951
transform 1 0 388 0 -1 505
box -2 -3 26 103
use INVX1  INVX1_67
timestamp 1626400951
transform 1 0 412 0 -1 505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_77
timestamp 1626400951
transform -1 0 524 0 -1 505
box -2 -3 98 103
use OR2X2  OR2X2_13
timestamp 1626400951
transform -1 0 556 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_9
timestamp 1626400951
transform 1 0 556 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_0_0
timestamp 1626400951
transform 1 0 588 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_0_1
timestamp 1626400951
transform 1 0 596 0 -1 505
box -2 -3 10 103
use INVX1  INVX1_103
timestamp 1626400951
transform 1 0 604 0 -1 505
box -2 -3 18 103
use NOR3X1  NOR3X1_2
timestamp 1626400951
transform -1 0 684 0 -1 505
box -2 -3 66 103
use NOR2X1  NOR2X1_75
timestamp 1626400951
transform 1 0 684 0 -1 505
box -2 -3 26 103
use INVX1  INVX1_102
timestamp 1626400951
transform -1 0 724 0 -1 505
box -2 -3 18 103
use INVX1  INVX1_101
timestamp 1626400951
transform 1 0 724 0 -1 505
box -2 -3 18 103
use NOR2X1  NOR2X1_74
timestamp 1626400951
transform 1 0 740 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_7
timestamp 1626400951
transform -1 0 796 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_90
timestamp 1626400951
transform 1 0 796 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_6
timestamp 1626400951
transform -1 0 924 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_6
timestamp 1626400951
transform 1 0 924 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_5
timestamp 1626400951
transform 1 0 956 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_5
timestamp 1626400951
transform -1 0 1020 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_3
timestamp 1626400951
transform 1 0 1020 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_3
timestamp 1626400951
transform 1 0 1052 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_1_0
timestamp 1626400951
transform -1 0 1092 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_1_1
timestamp 1626400951
transform -1 0 1100 0 -1 505
box -2 -3 10 103
use NAND3X1  NAND3X1_3
timestamp 1626400951
transform -1 0 1132 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_86
timestamp 1626400951
transform -1 0 1228 0 -1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_52
timestamp 1626400951
transform 1 0 1228 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_71
timestamp 1626400951
transform -1 0 1276 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_51
timestamp 1626400951
transform -1 0 1308 0 -1 505
box -2 -3 34 103
use AND2X2  AND2X2_10
timestamp 1626400951
transform 1 0 1308 0 -1 505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_1
timestamp 1626400951
transform -1 0 1412 0 -1 505
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_84
timestamp 1626400951
transform 1 0 1412 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_1
timestamp 1626400951
transform 1 0 1508 0 -1 505
box -2 -3 98 103
use FILL  FILL_4_2_0
timestamp 1626400951
transform 1 0 1604 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_2_1
timestamp 1626400951
transform 1 0 1612 0 -1 505
box -2 -3 10 103
use NOR2X1  NOR2X1_69
timestamp 1626400951
transform 1 0 1620 0 -1 505
box -2 -3 26 103
use INVX1  INVX1_97
timestamp 1626400951
transform -1 0 1660 0 -1 505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_111
timestamp 1626400951
transform -1 0 1756 0 -1 505
box -2 -3 98 103
use INVX1  INVX1_189
timestamp 1626400951
transform 1 0 1756 0 -1 505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_112
timestamp 1626400951
transform -1 0 1868 0 -1 505
box -2 -3 98 103
use AND2X2  AND2X2_29
timestamp 1626400951
transform 1 0 1868 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_115
timestamp 1626400951
transform 1 0 1900 0 -1 505
box -2 -3 98 103
use AND2X2  AND2X2_28
timestamp 1626400951
transform -1 0 2028 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_134
timestamp 1626400951
transform 1 0 2028 0 -1 505
box -2 -3 34 103
use BUFX2  BUFX2_34
timestamp 1626400951
transform 1 0 2060 0 -1 505
box -2 -3 26 103
use FILL  FILL_4_3_0
timestamp 1626400951
transform 1 0 2084 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_3_1
timestamp 1626400951
transform 1 0 2092 0 -1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_117
timestamp 1626400951
transform 1 0 2100 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_139
timestamp 1626400951
transform 1 0 2196 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_140
timestamp 1626400951
transform -1 0 2388 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_122
timestamp 1626400951
transform -1 0 2484 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_153
timestamp 1626400951
transform 1 0 2484 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_155
timestamp 1626400951
transform -1 0 2548 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_104
timestamp 1626400951
transform 1 0 2548 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_141
timestamp 1626400951
transform -1 0 2676 0 -1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_90
timestamp 1626400951
transform -1 0 2700 0 -1 505
box -2 -3 26 103
use FILL  FILL_5_1
timestamp 1626400951
transform -1 0 2708 0 -1 505
box -2 -3 10 103
use XNOR2X1  XNOR2X1_4
timestamp 1626400951
transform 1 0 4 0 1 305
box -2 -3 58 103
use XOR2X1  XOR2X1_3
timestamp 1626400951
transform 1 0 60 0 1 305
box -2 -3 58 103
use INVX1  INVX1_85
timestamp 1626400951
transform 1 0 116 0 1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_39
timestamp 1626400951
transform 1 0 132 0 1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_55
timestamp 1626400951
transform -1 0 180 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_45
timestamp 1626400951
transform -1 0 212 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_37
timestamp 1626400951
transform 1 0 212 0 1 305
box -2 -3 26 103
use INVX1  INVX1_65
timestamp 1626400951
transform 1 0 236 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_40
timestamp 1626400951
transform 1 0 252 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_39
timestamp 1626400951
transform 1 0 284 0 1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_49
timestamp 1626400951
transform -1 0 332 0 1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_26
timestamp 1626400951
transform -1 0 356 0 1 305
box -2 -3 26 103
use XNOR2X1  XNOR2X1_5
timestamp 1626400951
transform -1 0 412 0 1 305
box -2 -3 58 103
use INVX1  INVX1_115
timestamp 1626400951
transform 1 0 412 0 1 305
box -2 -3 18 103
use NOR2X1  NOR2X1_90
timestamp 1626400951
transform 1 0 428 0 1 305
box -2 -3 26 103
use INVX2  INVX2_9
timestamp 1626400951
transform 1 0 452 0 1 305
box -2 -3 18 103
use BUFX4  BUFX4_12
timestamp 1626400951
transform -1 0 500 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_50
timestamp 1626400951
transform -1 0 596 0 1 305
box -2 -3 98 103
use FILL  FILL_3_0_0
timestamp 1626400951
transform -1 0 604 0 1 305
box -2 -3 10 103
use FILL  FILL_3_0_1
timestamp 1626400951
transform -1 0 612 0 1 305
box -2 -3 10 103
use NAND3X1  NAND3X1_28
timestamp 1626400951
transform -1 0 644 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_54
timestamp 1626400951
transform 1 0 644 0 1 305
box -2 -3 26 103
use INVX1  INVX1_100
timestamp 1626400951
transform 1 0 668 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_62
timestamp 1626400951
transform 1 0 684 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_48
timestamp 1626400951
transform -1 0 812 0 1 305
box -2 -3 98 103
use NAND3X1  NAND3X1_6
timestamp 1626400951
transform 1 0 812 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_5
timestamp 1626400951
transform 1 0 844 0 1 305
box -2 -3 34 103
use NOR3X1  NOR3X1_1
timestamp 1626400951
transform -1 0 940 0 1 305
box -2 -3 66 103
use INVX1  INVX1_99
timestamp 1626400951
transform -1 0 956 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_60
timestamp 1626400951
transform -1 0 988 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_75
timestamp 1626400951
transform 1 0 988 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_83
timestamp 1626400951
transform 1 0 1020 0 1 305
box -2 -3 34 103
use FILL  FILL_3_1_0
timestamp 1626400951
transform 1 0 1052 0 1 305
box -2 -3 10 103
use FILL  FILL_3_1_1
timestamp 1626400951
transform 1 0 1060 0 1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_46
timestamp 1626400951
transform 1 0 1068 0 1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_81
timestamp 1626400951
transform 1 0 1164 0 1 305
box -2 -3 34 103
use AOI22X1  AOI22X1_22
timestamp 1626400951
transform -1 0 1236 0 1 305
box -2 -3 42 103
use NAND3X1  NAND3X1_27
timestamp 1626400951
transform 1 0 1236 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_100
timestamp 1626400951
transform 1 0 1268 0 1 305
box -2 -3 98 103
use AND2X2  AND2X2_13
timestamp 1626400951
transform 1 0 1364 0 1 305
box -2 -3 34 103
use OR2X2  OR2X2_17
timestamp 1626400951
transform -1 0 1428 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_101
timestamp 1626400951
transform 1 0 1428 0 1 305
box -2 -3 98 103
use NAND2X1  NAND2X1_50
timestamp 1626400951
transform 1 0 1524 0 1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_51
timestamp 1626400951
transform 1 0 1548 0 1 305
box -2 -3 26 103
use INVX1  INVX1_120
timestamp 1626400951
transform -1 0 1588 0 1 305
box -2 -3 18 103
use FILL  FILL_3_2_0
timestamp 1626400951
transform -1 0 1596 0 1 305
box -2 -3 10 103
use FILL  FILL_3_2_1
timestamp 1626400951
transform -1 0 1604 0 1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_68
timestamp 1626400951
transform -1 0 1700 0 1 305
box -2 -3 98 103
use INVX1  INVX1_109
timestamp 1626400951
transform 1 0 1700 0 1 305
box -2 -3 18 103
use NOR2X1  NOR2X1_84
timestamp 1626400951
transform 1 0 1716 0 1 305
box -2 -3 26 103
use INVX1  INVX1_40
timestamp 1626400951
transform -1 0 1756 0 1 305
box -2 -3 18 103
use BUFX4  BUFX4_11
timestamp 1626400951
transform 1 0 1756 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_121
timestamp 1626400951
transform 1 0 1788 0 1 305
box -2 -3 98 103
use AOI21X1  AOI21X1_66
timestamp 1626400951
transform 1 0 1884 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_85
timestamp 1626400951
transform 1 0 1916 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_120
timestamp 1626400951
transform 1 0 1948 0 1 305
box -2 -3 98 103
use AND2X2  AND2X2_27
timestamp 1626400951
transform 1 0 2044 0 1 305
box -2 -3 34 103
use FILL  FILL_3_3_0
timestamp 1626400951
transform 1 0 2076 0 1 305
box -2 -3 10 103
use FILL  FILL_3_3_1
timestamp 1626400951
transform 1 0 2084 0 1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_118
timestamp 1626400951
transform 1 0 2092 0 1 305
box -2 -3 98 103
use AND2X2  AND2X2_36
timestamp 1626400951
transform 1 0 2188 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_143
timestamp 1626400951
transform 1 0 2220 0 1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_161
timestamp 1626400951
transform -1 0 2348 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_112
timestamp 1626400951
transform 1 0 2348 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_162
timestamp 1626400951
transform -1 0 2412 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_199
timestamp 1626400951
transform 1 0 2412 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_110
timestamp 1626400951
transform -1 0 2468 0 1 305
box -2 -3 34 103
use INVX4  INVX4_4
timestamp 1626400951
transform -1 0 2492 0 1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_202
timestamp 1626400951
transform 1 0 2492 0 1 305
box -2 -3 26 103
use INVX1  INVX1_211
timestamp 1626400951
transform 1 0 2516 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_158
timestamp 1626400951
transform 1 0 2532 0 1 305
box -2 -3 34 103
use AND2X2  AND2X2_34
timestamp 1626400951
transform -1 0 2596 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_154
timestamp 1626400951
transform 1 0 2596 0 1 305
box -2 -3 34 103
use INVX1  INVX1_212
timestamp 1626400951
transform -1 0 2644 0 1 305
box -2 -3 18 103
use AOI21X1  AOI21X1_108
timestamp 1626400951
transform -1 0 2676 0 1 305
box -2 -3 34 103
use INVX1  INVX1_215
timestamp 1626400951
transform 1 0 2676 0 1 305
box -2 -3 18 103
use FILL  FILL_4_1
timestamp 1626400951
transform 1 0 2692 0 1 305
box -2 -3 10 103
use FILL  FILL_4_2
timestamp 1626400951
transform 1 0 2700 0 1 305
box -2 -3 10 103
use INVX1  INVX1_60
timestamp 1626400951
transform 1 0 4 0 -1 305
box -2 -3 18 103
use NOR2X1  NOR2X1_41
timestamp 1626400951
transform -1 0 44 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_21
timestamp 1626400951
transform 1 0 44 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_33
timestamp 1626400951
transform 1 0 68 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_40
timestamp 1626400951
transform -1 0 124 0 -1 305
box -2 -3 26 103
use INVX1  INVX1_59
timestamp 1626400951
transform -1 0 140 0 -1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_18
timestamp 1626400951
transform 1 0 140 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_32
timestamp 1626400951
transform -1 0 196 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_56
timestamp 1626400951
transform -1 0 212 0 -1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_20
timestamp 1626400951
transform -1 0 236 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_32
timestamp 1626400951
transform -1 0 268 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_38
timestamp 1626400951
transform -1 0 292 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_19
timestamp 1626400951
transform 1 0 292 0 -1 305
box -2 -3 26 103
use INVX1  INVX1_57
timestamp 1626400951
transform -1 0 332 0 -1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_78
timestamp 1626400951
transform 1 0 332 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_73
timestamp 1626400951
transform 1 0 428 0 -1 305
box -2 -3 98 103
use NOR2X1  NOR2X1_89
timestamp 1626400951
transform -1 0 548 0 -1 305
box -2 -3 26 103
use INVX1  INVX1_114
timestamp 1626400951
transform -1 0 564 0 -1 305
box -2 -3 18 103
use FILL  FILL_2_0_0
timestamp 1626400951
transform 1 0 564 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_0_1
timestamp 1626400951
transform 1 0 572 0 -1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_74
timestamp 1626400951
transform 1 0 580 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_61
timestamp 1626400951
transform 1 0 676 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_73
timestamp 1626400951
transform -1 0 732 0 -1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_89
timestamp 1626400951
transform 1 0 732 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_88
timestamp 1626400951
transform -1 0 924 0 -1 305
box -2 -3 98 103
use NOR2X1  NOR2X1_72
timestamp 1626400951
transform 1 0 924 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_53
timestamp 1626400951
transform -1 0 972 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_65
timestamp 1626400951
transform 1 0 972 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_75
timestamp 1626400951
transform 1 0 1004 0 -1 305
box -2 -3 26 103
use INVX2  INVX2_7
timestamp 1626400951
transform -1 0 1044 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_59
timestamp 1626400951
transform 1 0 1044 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_1_0
timestamp 1626400951
transform 1 0 1076 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_1_1
timestamp 1626400951
transform 1 0 1084 0 -1 305
box -2 -3 10 103
use AOI21X1  AOI21X1_52
timestamp 1626400951
transform 1 0 1092 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_87
timestamp 1626400951
transform 1 0 1124 0 -1 305
box -2 -3 98 103
use INVX1  INVX1_144
timestamp 1626400951
transform 1 0 1220 0 -1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_71
timestamp 1626400951
transform -1 0 1260 0 -1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_70
timestamp 1626400951
transform 1 0 1260 0 -1 305
box -2 -3 26 103
use OR2X2  OR2X2_9
timestamp 1626400951
transform -1 0 1316 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_68
timestamp 1626400951
transform 1 0 1316 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_57
timestamp 1626400951
transform -1 0 1364 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_84
timestamp 1626400951
transform -1 0 1396 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_146
timestamp 1626400951
transform -1 0 1412 0 -1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_102
timestamp 1626400951
transform -1 0 1508 0 -1 305
box -2 -3 98 103
use AOI21X1  AOI21X1_56
timestamp 1626400951
transform 1 0 1508 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_67
timestamp 1626400951
transform 1 0 1540 0 -1 305
box -2 -3 98 103
use FILL  FILL_2_2_0
timestamp 1626400951
transform 1 0 1636 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_2_1
timestamp 1626400951
transform 1 0 1644 0 -1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_71
timestamp 1626400951
transform 1 0 1652 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_103
timestamp 1626400951
transform 1 0 1684 0 -1 305
box -2 -3 98 103
use NOR2X1  NOR2X1_193
timestamp 1626400951
transform 1 0 1780 0 -1 305
box -2 -3 26 103
use INVX1  INVX1_205
timestamp 1626400951
transform -1 0 1820 0 -1 305
box -2 -3 18 103
use CLKBUF1  CLKBUF1_2
timestamp 1626400951
transform 1 0 1820 0 -1 305
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_145
timestamp 1626400951
transform 1 0 1892 0 -1 305
box -2 -3 98 103
use INVX2  INVX2_18
timestamp 1626400951
transform 1 0 1988 0 -1 305
box -2 -3 18 103
use MUX2X1  MUX2X1_6
timestamp 1626400951
transform -1 0 2052 0 -1 305
box -2 -3 50 103
use AND2X2  AND2X2_32
timestamp 1626400951
transform -1 0 2084 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_152
timestamp 1626400951
transform 1 0 2084 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_3_0
timestamp 1626400951
transform -1 0 2124 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_3_1
timestamp 1626400951
transform -1 0 2132 0 -1 305
box -2 -3 10 103
use INVX1  INVX1_208
timestamp 1626400951
transform -1 0 2148 0 -1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_149
timestamp 1626400951
transform -1 0 2172 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_146
timestamp 1626400951
transform 1 0 2172 0 -1 305
box -2 -3 26 103
use INVX2  INVX2_21
timestamp 1626400951
transform -1 0 2212 0 -1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_150
timestamp 1626400951
transform 1 0 2212 0 -1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_204
timestamp 1626400951
transform 1 0 2236 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_156
timestamp 1626400951
transform 1 0 2260 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_109
timestamp 1626400951
transform 1 0 2292 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_141
timestamp 1626400951
transform -1 0 2348 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_157
timestamp 1626400951
transform -1 0 2380 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_111
timestamp 1626400951
transform 1 0 2380 0 -1 305
box -2 -3 34 103
use INVX4  INVX4_5
timestamp 1626400951
transform -1 0 2436 0 -1 305
box -2 -3 26 103
use XNOR2X1  XNOR2X1_26
timestamp 1626400951
transform 1 0 2436 0 -1 305
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_138
timestamp 1626400951
transform 1 0 2492 0 -1 305
box -2 -3 98 103
use INVX1  INVX1_161
timestamp 1626400951
transform 1 0 2588 0 -1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_142
timestamp 1626400951
transform 1 0 2604 0 -1 305
box -2 -3 98 103
use FILL  FILL_3_1
timestamp 1626400951
transform -1 0 2708 0 -1 305
box -2 -3 10 103
use INVX1  INVX1_14
timestamp 1626400951
transform -1 0 20 0 1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_14
timestamp 1626400951
transform 1 0 20 0 1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_32
timestamp 1626400951
transform -1 0 140 0 1 105
box -2 -3 98 103
use NOR2X1  NOR2X1_9
timestamp 1626400951
transform -1 0 164 0 1 105
box -2 -3 26 103
use INVX1  INVX1_8
timestamp 1626400951
transform -1 0 180 0 1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_42
timestamp 1626400951
transform -1 0 276 0 1 105
box -2 -3 98 103
use BUFX2  BUFX2_37
timestamp 1626400951
transform 1 0 276 0 1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_75
timestamp 1626400951
transform 1 0 300 0 1 105
box -2 -3 98 103
use OR2X2  OR2X2_11
timestamp 1626400951
transform -1 0 428 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_88
timestamp 1626400951
transform -1 0 452 0 1 105
box -2 -3 26 103
use INVX1  INVX1_113
timestamp 1626400951
transform -1 0 468 0 1 105
box -2 -3 18 103
use INVX1  INVX1_141
timestamp 1626400951
transform 1 0 468 0 1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_103
timestamp 1626400951
transform -1 0 508 0 1 105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_15
timestamp 1626400951
transform -1 0 564 0 1 105
box -2 -3 58 103
use FILL  FILL_1_0_0
timestamp 1626400951
transform -1 0 572 0 1 105
box -2 -3 10 103
use FILL  FILL_1_0_1
timestamp 1626400951
transform -1 0 580 0 1 105
box -2 -3 10 103
use AOI21X1  AOI21X1_60
timestamp 1626400951
transform -1 0 612 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_70
timestamp 1626400951
transform 1 0 612 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_74
timestamp 1626400951
transform -1 0 668 0 1 105
box -2 -3 34 103
use INVX1  INVX1_132
timestamp 1626400951
transform 1 0 668 0 1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_73
timestamp 1626400951
transform 1 0 684 0 1 105
box -2 -3 34 103
use AOI22X1  AOI22X1_20
timestamp 1626400951
transform 1 0 716 0 1 105
box -2 -3 42 103
use INVX1  INVX1_133
timestamp 1626400951
transform -1 0 772 0 1 105
box -2 -3 18 103
use CLKBUF1  CLKBUF1_6
timestamp 1626400951
transform -1 0 844 0 1 105
box -2 -3 74 103
use NOR2X1  NOR2X1_109
timestamp 1626400951
transform -1 0 868 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_59
timestamp 1626400951
transform 1 0 868 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_82
timestamp 1626400951
transform -1 0 932 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_110
timestamp 1626400951
transform -1 0 956 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_80
timestamp 1626400951
transform -1 0 988 0 1 105
box -2 -3 34 103
use INVX1  INVX1_145
timestamp 1626400951
transform -1 0 1004 0 1 105
box -2 -3 18 103
use INVX1  INVX1_136
timestamp 1626400951
transform 1 0 1004 0 1 105
box -2 -3 18 103
use AOI21X1  AOI21X1_57
timestamp 1626400951
transform 1 0 1020 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_68
timestamp 1626400951
transform -1 0 1076 0 1 105
box -2 -3 26 103
use FILL  FILL_1_1_0
timestamp 1626400951
transform -1 0 1084 0 1 105
box -2 -3 10 103
use FILL  FILL_1_1_1
timestamp 1626400951
transform -1 0 1092 0 1 105
box -2 -3 10 103
use OAI21X1  OAI21X1_72
timestamp 1626400951
transform -1 0 1124 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_100
timestamp 1626400951
transform 1 0 1124 0 1 105
box -2 -3 26 103
use INVX1  INVX1_138
timestamp 1626400951
transform -1 0 1164 0 1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_99
timestamp 1626400951
transform 1 0 1164 0 1 105
box -2 -3 26 103
use INVX1  INVX1_148
timestamp 1626400951
transform 1 0 1188 0 1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_77
timestamp 1626400951
transform -1 0 1228 0 1 105
box -2 -3 26 103
use INVX1  INVX1_137
timestamp 1626400951
transform -1 0 1244 0 1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_70
timestamp 1626400951
transform -1 0 1340 0 1 105
box -2 -3 98 103
use INVX1  INVX1_111
timestamp 1626400951
transform 1 0 1340 0 1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_86
timestamp 1626400951
transform 1 0 1356 0 1 105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_18
timestamp 1626400951
transform -1 0 1436 0 1 105
box -2 -3 58 103
use INVX1  INVX1_112
timestamp 1626400951
transform 1 0 1436 0 1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_87
timestamp 1626400951
transform 1 0 1452 0 1 105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_3
timestamp 1626400951
transform 1 0 1476 0 1 105
box -2 -3 74 103
use BUFX4  BUFX4_10
timestamp 1626400951
transform -1 0 1580 0 1 105
box -2 -3 34 103
use INVX1  INVX1_110
timestamp 1626400951
transform 1 0 1580 0 1 105
box -2 -3 18 103
use FILL  FILL_1_2_0
timestamp 1626400951
transform 1 0 1596 0 1 105
box -2 -3 10 103
use FILL  FILL_1_2_1
timestamp 1626400951
transform 1 0 1604 0 1 105
box -2 -3 10 103
use NOR2X1  NOR2X1_85
timestamp 1626400951
transform 1 0 1612 0 1 105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_4
timestamp 1626400951
transform 1 0 1636 0 1 105
box -2 -3 74 103
use BUFX2  BUFX2_14
timestamp 1626400951
transform -1 0 1732 0 1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_23
timestamp 1626400951
transform -1 0 1828 0 1 105
box -2 -3 98 103
use INVX1  INVX1_22
timestamp 1626400951
transform 1 0 1828 0 1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_20
timestamp 1626400951
transform 1 0 1844 0 1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_205
timestamp 1626400951
transform -1 0 1892 0 1 105
box -2 -3 26 103
use AND2X2  AND2X2_35
timestamp 1626400951
transform 1 0 1892 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_159
timestamp 1626400951
transform 1 0 1924 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_144
timestamp 1626400951
transform 1 0 1956 0 1 105
box -2 -3 98 103
use MUX2X1  MUX2X1_7
timestamp 1626400951
transform -1 0 2100 0 1 105
box -2 -3 50 103
use INVX2  INVX2_20
timestamp 1626400951
transform 1 0 2100 0 1 105
box -2 -3 18 103
use FILL  FILL_1_3_0
timestamp 1626400951
transform -1 0 2124 0 1 105
box -2 -3 10 103
use FILL  FILL_1_3_1
timestamp 1626400951
transform -1 0 2132 0 1 105
box -2 -3 10 103
use OAI21X1  OAI21X1_160
timestamp 1626400951
transform -1 0 2164 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_147
timestamp 1626400951
transform 1 0 2164 0 1 105
box -2 -3 26 103
use AND2X2  AND2X2_33
timestamp 1626400951
transform 1 0 2188 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_198
timestamp 1626400951
transform -1 0 2244 0 1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_142
timestamp 1626400951
transform -1 0 2268 0 1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_197
timestamp 1626400951
transform 1 0 2268 0 1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_144
timestamp 1626400951
transform 1 0 2292 0 1 105
box -2 -3 26 103
use INVX1  INVX1_210
timestamp 1626400951
transform 1 0 2316 0 1 105
box -2 -3 18 103
use AOI22X1  AOI22X1_23
timestamp 1626400951
transform -1 0 2372 0 1 105
box -2 -3 42 103
use OAI21X1  OAI21X1_151
timestamp 1626400951
transform -1 0 2404 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_194
timestamp 1626400951
transform -1 0 2428 0 1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_148
timestamp 1626400951
transform -1 0 2452 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_163
timestamp 1626400951
transform 1 0 2452 0 1 105
box -2 -3 34 103
use INVX2  INVX2_19
timestamp 1626400951
transform -1 0 2500 0 1 105
box -2 -3 18 103
use INVX2  INVX2_17
timestamp 1626400951
transform 1 0 2500 0 1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_23
timestamp 1626400951
transform -1 0 2540 0 1 105
box -2 -3 26 103
use INVX1  INVX1_25
timestamp 1626400951
transform -1 0 2556 0 1 105
box -2 -3 18 103
use INVX1  INVX1_160
timestamp 1626400951
transform -1 0 2572 0 1 105
box -2 -3 18 103
use AOI21X1  AOI21X1_107
timestamp 1626400951
transform -1 0 2604 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_26
timestamp 1626400951
transform 1 0 2604 0 1 105
box -2 -3 98 103
use FILL  FILL_2_1
timestamp 1626400951
transform 1 0 2700 0 1 105
box -2 -3 10 103
use BUFX2  BUFX2_23
timestamp 1626400951
transform -1 0 28 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_30
timestamp 1626400951
transform -1 0 52 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_5
timestamp 1626400951
transform 1 0 52 0 -1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_6
timestamp 1626400951
transform 1 0 68 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_39
timestamp 1626400951
transform -1 0 188 0 -1 105
box -2 -3 98 103
use BUFX2  BUFX2_33
timestamp 1626400951
transform -1 0 212 0 -1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_8
timestamp 1626400951
transform -1 0 236 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_7
timestamp 1626400951
transform -1 0 252 0 -1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_41
timestamp 1626400951
transform 1 0 252 0 -1 105
box -2 -3 98 103
use BUFX2  BUFX2_32
timestamp 1626400951
transform 1 0 348 0 -1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_18
timestamp 1626400951
transform -1 0 396 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_20
timestamp 1626400951
transform -1 0 412 0 -1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_21
timestamp 1626400951
transform 1 0 412 0 -1 105
box -2 -3 98 103
use BUFX2  BUFX2_12
timestamp 1626400951
transform 1 0 508 0 -1 105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_14
timestamp 1626400951
transform 1 0 532 0 -1 105
box -2 -3 58 103
use FILL  FILL_0_0_0
timestamp 1626400951
transform 1 0 588 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_0_1
timestamp 1626400951
transform 1 0 596 0 -1 105
box -2 -3 10 103
use NOR2X1  NOR2X1_104
timestamp 1626400951
transform 1 0 604 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_142
timestamp 1626400951
transform -1 0 644 0 -1 105
box -2 -3 18 103
use XOR2X1  XOR2X1_7
timestamp 1626400951
transform -1 0 700 0 -1 105
box -2 -3 58 103
use XOR2X1  XOR2X1_8
timestamp 1626400951
transform 1 0 700 0 -1 105
box -2 -3 58 103
use NOR2X1  NOR2X1_97
timestamp 1626400951
transform -1 0 780 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_134
timestamp 1626400951
transform 1 0 780 0 -1 105
box -2 -3 18 103
use OAI22X1  OAI22X1_5
timestamp 1626400951
transform 1 0 796 0 -1 105
box -2 -3 42 103
use AOI22X1  AOI22X1_21
timestamp 1626400951
transform 1 0 836 0 -1 105
box -2 -3 42 103
use INVX1  INVX1_135
timestamp 1626400951
transform -1 0 892 0 -1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_73
timestamp 1626400951
transform -1 0 916 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_65
timestamp 1626400951
transform 1 0 916 0 -1 105
box -2 -3 26 103
use AND2X2  AND2X2_12
timestamp 1626400951
transform 1 0 940 0 -1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_58
timestamp 1626400951
transform -1 0 1004 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_101
timestamp 1626400951
transform -1 0 1028 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_69
timestamp 1626400951
transform -1 0 1052 0 -1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_102
timestamp 1626400951
transform 1 0 1052 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_140
timestamp 1626400951
transform -1 0 1092 0 -1 105
box -2 -3 18 103
use FILL  FILL_0_1_0
timestamp 1626400951
transform -1 0 1100 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_1_1
timestamp 1626400951
transform -1 0 1108 0 -1 105
box -2 -3 10 103
use XNOR2X1  XNOR2X1_16
timestamp 1626400951
transform -1 0 1164 0 -1 105
box -2 -3 58 103
use NAND2X1  NAND2X1_66
timestamp 1626400951
transform -1 0 1188 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_139
timestamp 1626400951
transform -1 0 1204 0 -1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_98
timestamp 1626400951
transform 1 0 1204 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_67
timestamp 1626400951
transform -1 0 1252 0 -1 105
box -2 -3 26 103
use XOR2X1  XOR2X1_9
timestamp 1626400951
transform -1 0 1308 0 -1 105
box -2 -3 58 103
use AOI21X1  AOI21X1_64
timestamp 1626400951
transform 1 0 1308 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_111
timestamp 1626400951
transform 1 0 1340 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_76
timestamp 1626400951
transform 1 0 1364 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_147
timestamp 1626400951
transform -1 0 1404 0 -1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_74
timestamp 1626400951
transform -1 0 1428 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_72
timestamp 1626400951
transform -1 0 1524 0 -1 105
box -2 -3 98 103
use XNOR2X1  XNOR2X1_17
timestamp 1626400951
transform -1 0 1580 0 -1 105
box -2 -3 58 103
use FILL  FILL_0_2_0
timestamp 1626400951
transform -1 0 1588 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_2_1
timestamp 1626400951
transform -1 0 1596 0 -1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_69
timestamp 1626400951
transform -1 0 1692 0 -1 105
box -2 -3 98 103
use OR2X2  OR2X2_10
timestamp 1626400951
transform 1 0 1692 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_71
timestamp 1626400951
transform -1 0 1820 0 -1 105
box -2 -3 98 103
use BUFX2  BUFX2_29
timestamp 1626400951
transform -1 0 1844 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_38
timestamp 1626400951
transform -1 0 1940 0 -1 105
box -2 -3 98 103
use INVX1  INVX1_4
timestamp 1626400951
transform 1 0 1940 0 -1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_5
timestamp 1626400951
transform 1 0 1956 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_19
timestamp 1626400951
transform 1 0 1980 0 -1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_10
timestamp 1626400951
transform -1 0 2028 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_10
timestamp 1626400951
transform -1 0 2044 0 -1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_28
timestamp 1626400951
transform 1 0 2044 0 -1 105
box -2 -3 98 103
use FILL  FILL_0_3_0
timestamp 1626400951
transform -1 0 2148 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_3_1
timestamp 1626400951
transform -1 0 2156 0 -1 105
box -2 -3 10 103
use INVX2  INVX2_16
timestamp 1626400951
transform -1 0 2172 0 -1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_146
timestamp 1626400951
transform -1 0 2268 0 -1 105
box -2 -3 98 103
use INVX1  INVX1_204
timestamp 1626400951
transform 1 0 2268 0 -1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_5
timestamp 1626400951
transform -1 0 2332 0 -1 105
box -2 -3 50 103
use INVX1  INVX1_206
timestamp 1626400951
transform 1 0 2332 0 -1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_196
timestamp 1626400951
transform -1 0 2372 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_207
timestamp 1626400951
transform -1 0 2388 0 -1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_195
timestamp 1626400951
transform -1 0 2412 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_214
timestamp 1626400951
transform 1 0 2412 0 -1 105
box -2 -3 18 103
use OAI22X1  OAI22X1_9
timestamp 1626400951
transform -1 0 2468 0 -1 105
box -2 -3 42 103
use NAND2X1  NAND2X1_145
timestamp 1626400951
transform -1 0 2492 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_213
timestamp 1626400951
transform 1 0 2492 0 -1 105
box -2 -3 18 103
use AOI21X1  AOI21X1_105
timestamp 1626400951
transform 1 0 2508 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_201
timestamp 1626400951
transform -1 0 2564 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_209
timestamp 1626400951
transform -1 0 2580 0 -1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_200
timestamp 1626400951
transform 1 0 2580 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_143
timestamp 1626400951
transform 1 0 2604 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_106
timestamp 1626400951
transform 1 0 2628 0 -1 105
box -2 -3 34 103
use BUFX2  BUFX2_17
timestamp 1626400951
transform -1 0 2684 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_154
timestamp 1626400951
transform 1 0 2684 0 -1 105
box -2 -3 18 103
use FILL  FILL_1_1
timestamp 1626400951
transform -1 0 2708 0 -1 105
box -2 -3 10 103
<< labels >>
flabel metal6 s 576 -30 592 -22 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal6 s 1080 -30 1096 -22 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal2 s 838 -22 842 -18 7 FreeSans 24 270 0 0 clk
port 2 nsew
flabel metal2 s 742 1828 746 1832 3 FreeSans 24 90 0 0 reset
port 3 nsew
flabel metal3 s 2734 678 2738 682 3 FreeSans 24 0 0 0 block0[0]
port 4 nsew
flabel metal2 s 254 1828 258 1832 3 FreeSans 24 90 0 0 block0[1]
port 5 nsew
flabel metal2 s 598 -22 602 -18 7 FreeSans 24 270 0 0 block0[2]
port 6 nsew
flabel metal3 s 2734 1728 2738 1732 3 FreeSans 24 0 0 0 block0[3]
port 7 nsew
flabel metal3 s 2734 1248 2738 1252 3 FreeSans 24 0 0 0 block0[4]
port 8 nsew
flabel metal3 s 2734 868 2738 872 3 FreeSans 24 0 0 0 block0[5]
port 9 nsew
flabel metal3 s -26 1678 -22 1682 7 FreeSans 24 0 0 0 block0[6]
port 10 nsew
flabel metal3 s -26 528 -22 532 7 FreeSans 24 0 0 0 block0[7]
port 11 nsew
flabel metal3 s 2734 468 2738 472 3 FreeSans 24 0 0 0 block1[0]
port 12 nsew
flabel metal2 s 2518 -22 2522 -18 7 FreeSans 24 270 0 0 block1[1]
port 13 nsew
flabel metal2 s 2382 1828 2386 1832 3 FreeSans 24 90 0 0 block1[2]
port 14 nsew
flabel metal3 s 2734 978 2738 982 3 FreeSans 24 0 0 0 block1[3]
port 15 nsew
flabel metal2 s 1566 -22 1570 -18 7 FreeSans 24 270 0 0 block1[4]
port 16 nsew
flabel metal3 s -26 718 -22 722 7 FreeSans 24 0 0 0 block1[5]
port 17 nsew
flabel metal3 s -26 1508 -22 1512 7 FreeSans 24 0 0 0 block1[6]
port 18 nsew
flabel metal3 s -26 468 -22 472 7 FreeSans 24 0 0 0 block1[7]
port 19 nsew
flabel metal3 s 2734 588 2738 592 3 FreeSans 24 0 0 0 block2[0]
port 20 nsew
flabel metal2 s 46 -22 50 -18 7 FreeSans 24 270 0 0 block2[1]
port 21 nsew
flabel metal2 s 2182 -22 2186 -18 7 FreeSans 24 270 0 0 block2[2]
port 22 nsew
flabel metal2 s 758 -22 762 -18 7 FreeSans 24 270 0 0 block2[3]
port 23 nsew
flabel metal3 s -26 818 -22 822 7 FreeSans 24 0 0 0 block2[4]
port 24 nsew
flabel metal2 s 1766 1828 1770 1832 3 FreeSans 24 90 0 0 block2[5]
port 25 nsew
flabel metal3 s 2734 1668 2738 1672 3 FreeSans 24 0 0 0 block2[6]
port 26 nsew
flabel metal3 s -26 28 -22 32 7 FreeSans 24 270 0 0 block2[7]
port 27 nsew
flabel metal3 s 2734 748 2738 752 3 FreeSans 24 0 0 0 block3[0]
port 28 nsew
flabel metal2 s 1726 1828 1730 1832 3 FreeSans 24 90 0 0 block3[1]
port 29 nsew
flabel metal3 s -26 988 -22 992 7 FreeSans 24 0 0 0 block3[2]
port 30 nsew
flabel metal3 s 2734 78 2738 82 3 FreeSans 24 0 0 0 block3[3]
port 31 nsew
flabel metal2 s 1958 1828 1962 1832 3 FreeSans 24 90 0 0 block3[4]
port 32 nsew
flabel metal2 s 734 -22 738 -18 7 FreeSans 24 270 0 0 block3[5]
port 33 nsew
flabel metal2 s 1830 1828 1834 1832 3 FreeSans 24 90 0 0 block3[6]
port 34 nsew
flabel metal3 s 2734 918 2738 922 3 FreeSans 24 0 0 0 block3[7]
port 35 nsew
flabel metal3 s 2734 938 2738 942 3 FreeSans 24 0 0 0 block4[0]
port 36 nsew
flabel metal2 s 822 1828 826 1832 3 FreeSans 24 90 0 0 block4[1]
port 37 nsew
flabel metal2 s 1486 -22 1490 -18 7 FreeSans 24 270 0 0 block4[2]
port 38 nsew
flabel metal2 s 102 1828 106 1832 3 FreeSans 24 90 0 0 block4[3]
port 39 nsew
flabel metal3 s 2734 1108 2738 1112 3 FreeSans 24 0 0 0 block4[4]
port 40 nsew
flabel metal3 s -26 128 -22 132 7 FreeSans 24 0 0 0 block4[5]
port 41 nsew
flabel metal3 s 2734 618 2738 622 3 FreeSans 24 0 0 0 block4[6]
port 42 nsew
flabel metal3 s 2734 498 2738 502 3 FreeSans 24 0 0 0 block4[7]
port 43 nsew
flabel metal3 s 2734 888 2738 892 3 FreeSans 24 0 0 0 block5[0]
port 44 nsew
flabel metal3 s 2734 568 2738 572 3 FreeSans 24 0 0 0 block5[1]
port 45 nsew
flabel metal2 s 534 -22 538 -18 7 FreeSans 24 270 0 0 block5[2]
port 46 nsew
flabel metal2 s 294 1828 298 1832 3 FreeSans 24 90 0 0 block5[3]
port 47 nsew
flabel metal3 s -26 1658 -22 1662 7 FreeSans 24 0 0 0 block5[4]
port 48 nsew
flabel metal2 s 2334 -22 2338 -18 7 FreeSans 24 270 0 0 block5[5]
port 49 nsew
flabel metal3 s -26 1288 -22 1292 7 FreeSans 24 0 0 0 block5[6]
port 50 nsew
flabel metal3 s -26 298 -22 302 7 FreeSans 24 0 0 0 block5[7]
port 51 nsew
flabel metal3 s 2734 1148 2738 1152 3 FreeSans 24 0 0 0 block6[0]
port 52 nsew
flabel metal3 s -26 778 -22 782 7 FreeSans 24 0 0 0 block6[1]
port 53 nsew
flabel metal3 s -26 1458 -22 1462 7 FreeSans 24 0 0 0 block6[2]
port 54 nsew
flabel metal2 s 1350 1828 1354 1832 3 FreeSans 24 90 0 0 block6[3]
port 55 nsew
flabel metal3 s 2734 1068 2738 1072 3 FreeSans 24 0 0 0 block6[4]
port 56 nsew
flabel metal3 s -26 168 -22 172 7 FreeSans 24 0 0 0 block6[5]
port 57 nsew
flabel metal3 s -26 908 -22 912 7 FreeSans 24 0 0 0 block6[6]
port 58 nsew
flabel metal2 s 1942 1828 1946 1832 3 FreeSans 24 90 0 0 block6[7]
port 59 nsew
flabel metal3 s 2734 548 2738 552 3 FreeSans 24 0 0 0 block7[0]
port 60 nsew
flabel metal3 s 2734 268 2738 272 3 FreeSans 24 0 0 0 block7[1]
port 61 nsew
flabel metal2 s 78 1828 82 1832 3 FreeSans 24 90 0 0 block7[2]
port 62 nsew
flabel metal3 s 2734 1128 2738 1132 3 FreeSans 24 0 0 0 block7[3]
port 63 nsew
flabel metal3 s 2734 1338 2738 1342 3 FreeSans 24 0 0 0 block7[4]
port 64 nsew
flabel metal3 s -26 648 -22 652 7 FreeSans 24 0 0 0 block7[5]
port 65 nsew
flabel metal3 s -26 928 -22 932 7 FreeSans 24 0 0 0 block7[6]
port 66 nsew
flabel metal3 s 2734 248 2738 252 3 FreeSans 24 0 0 0 block7[7]
port 67 nsew
flabel metal3 s 2734 1268 2738 1272 3 FreeSans 24 0 0 0 block8[0]
port 68 nsew
flabel metal3 s -26 508 -22 512 7 FreeSans 24 0 0 0 block8[1]
port 69 nsew
flabel metal3 s 2734 448 2738 452 3 FreeSans 24 0 0 0 block8[2]
port 70 nsew
flabel metal3 s -26 1568 -22 1572 7 FreeSans 24 0 0 0 block8[3]
port 71 nsew
flabel metal2 s 2406 -22 2410 -18 7 FreeSans 24 270 0 0 block8[4]
port 72 nsew
flabel metal3 s -26 1748 -22 1752 7 FreeSans 24 90 0 0 block8[5]
port 73 nsew
flabel metal3 s 2734 1638 2738 1642 3 FreeSans 24 0 0 0 block8[6]
port 74 nsew
flabel metal2 s 46 1828 50 1832 7 FreeSans 24 90 0 0 block8[7]
port 75 nsew
flabel metal3 s 2734 958 2738 962 3 FreeSans 24 0 0 0 block9[0]
port 76 nsew
flabel metal2 s 2086 1828 2090 1832 3 FreeSans 24 90 0 0 block9[1]
port 77 nsew
flabel metal3 s -26 98 -22 102 7 FreeSans 24 0 0 0 block9[2]
port 78 nsew
flabel metal2 s 614 -22 618 -18 7 FreeSans 24 270 0 0 block9[3]
port 79 nsew
flabel metal2 s 1750 1828 1754 1832 3 FreeSans 24 90 0 0 block9[4]
port 80 nsew
flabel metal3 s -26 1698 -22 1702 7 FreeSans 24 0 0 0 block9[5]
port 81 nsew
flabel metal3 s -26 1638 -22 1642 7 FreeSans 24 0 0 0 block9[6]
port 82 nsew
flabel metal3 s -26 1148 -22 1152 7 FreeSans 24 0 0 0 block9[7]
port 83 nsew
flabel metal3 s 2734 1688 2738 1692 3 FreeSans 24 0 0 0 block10[0]
port 84 nsew
flabel metal2 s 2582 1828 2586 1832 3 FreeSans 24 90 0 0 block10[1]
port 85 nsew
flabel metal2 s 1278 1828 1282 1832 3 FreeSans 24 90 0 0 block10[2]
port 86 nsew
flabel metal2 s 1982 1828 1986 1832 3 FreeSans 24 90 0 0 block10[3]
port 87 nsew
flabel metal2 s 638 1828 642 1832 3 FreeSans 24 90 0 0 block10[4]
port 88 nsew
flabel metal3 s -26 1588 -22 1592 7 FreeSans 24 0 0 0 block10[5]
port 89 nsew
flabel metal3 s 2734 28 2738 32 3 FreeSans 24 270 0 0 block10[6]
port 90 nsew
flabel metal2 s 862 1828 866 1832 3 FreeSans 24 90 0 0 block10[7]
port 91 nsew
flabel metal3 s 2734 1088 2738 1092 3 FreeSans 24 0 0 0 block11[0]
port 92 nsew
flabel metal2 s 1838 -22 1842 -18 7 FreeSans 24 270 0 0 block11[1]
port 93 nsew
flabel metal3 s -26 148 -22 152 7 FreeSans 24 0 0 0 block11[2]
port 94 nsew
flabel metal3 s -26 948 -22 952 7 FreeSans 24 0 0 0 block11[3]
port 95 nsew
flabel metal2 s 2054 -22 2058 -18 7 FreeSans 24 270 0 0 block11[4]
port 96 nsew
flabel metal2 s 1934 -22 1938 -18 7 FreeSans 24 270 0 0 block11[5]
port 97 nsew
flabel metal2 s 1238 -22 1242 -18 7 FreeSans 24 270 0 0 block11[6]
port 98 nsew
flabel metal2 s 598 1828 602 1832 3 FreeSans 24 90 0 0 block11[7]
port 99 nsew
flabel metal2 s 934 1828 938 1832 3 FreeSans 24 90 0 0 start
port 100 nsew
flabel metal3 s -26 488 -22 492 7 FreeSans 24 0 0 0 target[0]
port 101 nsew
flabel metal3 s -26 358 -22 362 7 FreeSans 24 0 0 0 target[1]
port 102 nsew
flabel metal3 s -26 278 -22 282 7 FreeSans 24 0 0 0 target[2]
port 103 nsew
flabel metal3 s -26 668 -22 672 7 FreeSans 24 0 0 0 target[3]
port 104 nsew
flabel metal3 s -26 758 -22 762 7 FreeSans 24 0 0 0 target[4]
port 105 nsew
flabel metal3 s -26 968 -22 972 7 FreeSans 24 0 0 0 target[5]
port 106 nsew
flabel metal3 s -26 1168 -22 1172 7 FreeSans 24 0 0 0 target[6]
port 107 nsew
flabel metal3 s -26 1128 -22 1132 7 FreeSans 24 0 0 0 target[7]
port 108 nsew
flabel metal3 s -26 1548 -22 1552 7 FreeSans 24 0 0 0 target[8]
port 109 nsew
flabel metal3 s -26 1728 -22 1732 7 FreeSans 24 0 0 0 target[9]
port 110 nsew
flabel metal3 s -26 1348 -22 1352 7 FreeSans 24 0 0 0 target[10]
port 111 nsew
flabel metal3 s -26 1248 -22 1252 7 FreeSans 24 0 0 0 target[11]
port 112 nsew
flabel metal2 s 182 1828 186 1832 3 FreeSans 24 90 0 0 target[12]
port 113 nsew
flabel metal2 s 222 1828 226 1832 3 FreeSans 24 90 0 0 target[13]
port 114 nsew
flabel metal2 s 406 1828 410 1832 3 FreeSans 24 90 0 0 target[14]
port 115 nsew
flabel metal2 s 366 1828 370 1832 3 FreeSans 24 90 0 0 target[15]
port 116 nsew
flabel metal2 s 1526 1828 1530 1832 3 FreeSans 24 90 0 0 nonce0[0]
port 117 nsew
flabel metal2 s 1558 1828 1562 1832 3 FreeSans 24 90 0 0 nonce0[1]
port 118 nsew
flabel metal2 s 774 1828 778 1832 3 FreeSans 24 90 0 0 nonce0[2]
port 119 nsew
flabel metal2 s 1126 1828 1130 1832 3 FreeSans 24 90 0 0 nonce0[3]
port 120 nsew
flabel metal2 s 838 1828 842 1832 3 FreeSans 24 90 0 0 nonce0[4]
port 121 nsew
flabel metal2 s 758 1828 762 1832 3 FreeSans 24 90 0 0 nonce0[5]
port 122 nsew
flabel metal2 s 1478 1828 1482 1832 3 FreeSans 24 90 0 0 nonce0[6]
port 123 nsew
flabel metal2 s 502 1828 506 1832 3 FreeSans 24 90 0 0 nonce0[7]
port 124 nsew
flabel metal2 s 1102 1828 1106 1832 3 FreeSans 24 90 0 0 nonce1[0]
port 125 nsew
flabel metal2 s 454 1828 458 1832 3 FreeSans 24 90 0 0 nonce1[1]
port 126 nsew
flabel metal2 s 550 -22 554 -18 7 FreeSans 24 270 0 0 nonce1[2]
port 127 nsew
flabel metal2 s 966 1828 970 1832 3 FreeSans 24 90 0 0 nonce1[3]
port 128 nsew
flabel metal2 s 1718 -22 1722 -18 7 FreeSans 24 270 0 0 nonce1[4]
port 129 nsew
flabel metal2 s 2686 1828 2690 1832 3 FreeSans 24 90 0 0 nonce1[5]
port 130 nsew
flabel metal2 s 1886 1828 1890 1832 3 FreeSans 24 90 0 0 nonce1[6]
port 131 nsew
flabel metal2 s 2670 -22 2674 -18 3 FreeSans 24 270 0 0 nonce1[7]
port 132 nsew
flabel metal2 s 1502 1828 1506 1832 3 FreeSans 24 90 0 0 nonce2[0]
port 133 nsew
flabel metal2 s 1990 -22 1994 -18 7 FreeSans 24 270 0 0 nonce2[1]
port 134 nsew
flabel metal2 s 1702 1828 1706 1832 3 FreeSans 24 90 0 0 nonce2[2]
port 135 nsew
flabel metal2 s 1246 1828 1250 1832 3 FreeSans 24 90 0 0 nonce2[3]
port 136 nsew
flabel metal2 s 1310 1828 1314 1832 3 FreeSans 24 90 0 0 nonce2[4]
port 137 nsew
flabel metal3 s -26 68 -22 72 7 FreeSans 24 0 0 0 nonce2[5]
port 138 nsew
flabel metal2 s 950 1828 954 1832 3 FreeSans 24 90 0 0 nonce2[6]
port 139 nsew
flabel metal2 s 1454 1828 1458 1832 3 FreeSans 24 90 0 0 nonce2[7]
port 140 nsew
flabel metal2 s 1430 1828 1434 1832 3 FreeSans 24 90 0 0 nonce3[0]
port 141 nsew
flabel metal2 s 790 1828 794 1832 3 FreeSans 24 90 0 0 nonce3[1]
port 142 nsew
flabel metal2 s 1678 1828 1682 1832 3 FreeSans 24 90 0 0 nonce3[2]
port 143 nsew
flabel metal2 s 1822 -22 1826 -18 7 FreeSans 24 270 0 0 nonce3[3]
port 144 nsew
flabel metal3 s -26 48 -22 52 7 FreeSans 24 270 0 0 nonce3[4]
port 145 nsew
flabel metal2 s 1782 1828 1786 1832 3 FreeSans 24 90 0 0 nonce3[5]
port 146 nsew
flabel metal2 s 358 -22 362 -18 7 FreeSans 24 270 0 0 nonce3[6]
port 147 nsew
flabel metal2 s 198 -22 202 -18 7 FreeSans 24 270 0 0 nonce3[7]
port 148 nsew
flabel metal2 s 1222 1828 1226 1832 3 FreeSans 24 90 0 0 finish
port 149 nsew
<< end >>
