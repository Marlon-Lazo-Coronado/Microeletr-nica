VERSION 5.3 ;
   NAMESCASESENSITIVE ON ;
   NOWIREEXTENSIONATPIN ON ;
   DIVIDERCHAR "/" ;
   BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO area_sys
   CLASS BLOCK ;
   FOREIGN area_sys ;
   ORIGIN 2.6000 3.0000 ;
   SIZE 276.4000 BY 186.2000 ;
   PIN vdd
      PORT
         LAYER metal1 ;
	    RECT 0.2000 180.2000 271.0000 180.8000 ;
	    RECT 0.6000 177.9000 1.0000 180.2000 ;
	    RECT 2.2000 175.9000 2.6000 180.2000 ;
	    RECT 5.4000 175.9000 5.8000 180.2000 ;
	    RECT 6.2000 177.9000 6.6000 180.2000 ;
	    RECT 7.8000 177.9000 8.2000 180.2000 ;
	    RECT 8.6000 177.9000 9.0000 180.2000 ;
	    RECT 10.2000 177.9000 10.6000 180.2000 ;
	    RECT 11.8000 177.9000 12.2000 180.2000 ;
	    RECT 12.6000 177.9000 13.0000 180.2000 ;
	    RECT 14.2000 177.9000 14.6000 180.2000 ;
	    RECT 15.8000 177.9000 16.2000 180.2000 ;
	    RECT 16.6000 177.9000 17.0000 180.2000 ;
	    RECT 20.6000 176.5000 21.0000 180.2000 ;
	    RECT 23.0000 177.9000 23.4000 180.2000 ;
	    RECT 25.4000 175.9000 25.8000 180.2000 ;
	    RECT 26.2000 177.9000 26.6000 180.2000 ;
	    RECT 27.8000 177.9000 28.2000 180.2000 ;
	    RECT 29.4000 177.9000 29.8000 180.2000 ;
	    RECT 31.5000 175.9000 31.9000 180.2000 ;
	    RECT 33.4000 177.9000 33.8000 180.2000 ;
	    RECT 35.0000 177.9000 35.4000 180.2000 ;
	    RECT 36.6000 177.9000 37.0000 180.2000 ;
	    RECT 37.4000 177.9000 37.8000 180.2000 ;
	    RECT 39.0000 177.9000 39.4000 180.2000 ;
	    RECT 40.6000 177.9000 41.0000 180.2000 ;
	    RECT 41.4000 177.9000 41.8000 180.2000 ;
	    RECT 43.0000 177.9000 43.4000 180.2000 ;
	    RECT 44.6000 177.9000 45.0000 180.2000 ;
	    RECT 45.4000 177.9000 45.8000 180.2000 ;
	    RECT 47.0000 177.9000 47.4000 180.2000 ;
	    RECT 48.6000 177.9000 49.0000 180.2000 ;
	    RECT 50.2000 176.5000 50.6000 180.2000 ;
	    RECT 52.6000 175.9000 53.0000 180.2000 ;
	    RECT 55.4000 177.9000 55.8000 180.2000 ;
	    RECT 57.0000 177.9000 57.4000 180.2000 ;
	    RECT 59.8000 176.0000 60.2000 180.2000 ;
	    RECT 63.8000 176.0000 64.2000 180.2000 ;
	    RECT 66.6000 177.9000 67.0000 180.2000 ;
	    RECT 68.2000 177.9000 68.6000 180.2000 ;
	    RECT 71.0000 175.9000 71.4000 180.2000 ;
	    RECT 73.4000 176.5000 73.8000 180.2000 ;
	    RECT 75.8000 176.5000 76.2000 180.2000 ;
	    RECT 78.2000 176.5000 78.6000 180.2000 ;
	    RECT 80.6000 176.0000 81.0000 180.2000 ;
	    RECT 83.4000 177.9000 83.8000 180.2000 ;
	    RECT 85.0000 177.9000 85.4000 180.2000 ;
	    RECT 87.8000 175.9000 88.2000 180.2000 ;
	    RECT 89.4000 177.9000 89.8000 180.2000 ;
	    RECT 91.0000 175.9000 91.4000 180.2000 ;
	    RECT 94.2000 176.5000 94.6000 180.2000 ;
	    RECT 96.6000 176.5000 97.0000 180.2000 ;
	    RECT 99.0000 176.0000 99.4000 180.2000 ;
	    RECT 101.8000 177.9000 102.2000 180.2000 ;
	    RECT 103.4000 177.9000 103.8000 180.2000 ;
	    RECT 106.2000 175.9000 106.6000 180.2000 ;
	    RECT 108.6000 176.5000 109.0000 180.2000 ;
	    RECT 112.6000 176.5000 113.0000 180.2000 ;
	    RECT 115.0000 175.9000 115.4000 180.2000 ;
	    RECT 117.8000 177.9000 118.2000 180.2000 ;
	    RECT 119.4000 177.9000 119.8000 180.2000 ;
	    RECT 122.2000 176.0000 122.6000 180.2000 ;
	    RECT 124.6000 176.5000 125.0000 180.2000 ;
	    RECT 127.8000 175.9000 128.2000 180.2000 ;
	    RECT 129.4000 177.9000 129.8000 180.2000 ;
	    RECT 131.0000 176.5000 131.4000 180.2000 ;
	    RECT 133.4000 176.0000 133.8000 180.2000 ;
	    RECT 136.2000 177.9000 136.6000 180.2000 ;
	    RECT 137.8000 177.9000 138.2000 180.2000 ;
	    RECT 140.6000 175.9000 141.0000 180.2000 ;
	    RECT 143.0000 176.5000 143.4000 180.2000 ;
	    RECT 145.4000 176.5000 145.8000 180.2000 ;
	    RECT 147.8000 176.5000 148.2000 180.2000 ;
	    RECT 150.2000 176.5000 150.6000 180.2000 ;
	    RECT 152.6000 176.5000 153.0000 180.2000 ;
	    RECT 155.0000 175.9000 155.4000 180.2000 ;
	    RECT 157.8000 177.9000 158.2000 180.2000 ;
	    RECT 159.4000 177.9000 159.8000 180.2000 ;
	    RECT 162.2000 176.0000 162.6000 180.2000 ;
	    RECT 165.4000 177.9000 165.8000 180.2000 ;
	    RECT 167.8000 176.5000 168.2000 180.2000 ;
	    RECT 170.2000 176.5000 170.6000 180.2000 ;
	    RECT 172.6000 176.5000 173.0000 180.2000 ;
	    RECT 175.0000 176.0000 175.4000 180.2000 ;
	    RECT 177.8000 177.9000 178.2000 180.2000 ;
	    RECT 179.4000 177.9000 179.8000 180.2000 ;
	    RECT 182.2000 175.9000 182.6000 180.2000 ;
	    RECT 185.4000 175.9000 185.8000 180.2000 ;
	    RECT 187.0000 177.9000 187.4000 180.2000 ;
	    RECT 188.6000 176.5000 189.0000 180.2000 ;
	    RECT 191.0000 176.0000 191.4000 180.2000 ;
	    RECT 193.8000 177.9000 194.2000 180.2000 ;
	    RECT 195.4000 177.9000 195.8000 180.2000 ;
	    RECT 198.2000 175.9000 198.6000 180.2000 ;
	    RECT 199.8000 175.9000 200.2000 180.2000 ;
	    RECT 201.9000 177.9000 202.3000 180.2000 ;
	    RECT 203.8000 176.5000 204.2000 180.2000 ;
	    RECT 207.0000 176.0000 207.4000 180.2000 ;
	    RECT 209.8000 177.9000 210.2000 180.2000 ;
	    RECT 211.4000 177.9000 211.8000 180.2000 ;
	    RECT 214.2000 175.9000 214.6000 180.2000 ;
	    RECT 219.0000 175.9000 219.4000 180.2000 ;
	    RECT 219.8000 175.9000 220.2000 180.2000 ;
	    RECT 221.9000 177.9000 222.3000 180.2000 ;
	    RECT 223.0000 177.9000 223.4000 180.2000 ;
	    RECT 224.6000 177.9000 225.0000 180.2000 ;
	    RECT 226.2000 176.5000 226.6000 180.2000 ;
	    RECT 229.4000 176.0000 229.8000 180.2000 ;
	    RECT 232.2000 177.9000 232.6000 180.2000 ;
	    RECT 233.8000 177.9000 234.2000 180.2000 ;
	    RECT 236.6000 175.9000 237.0000 180.2000 ;
	    RECT 238.2000 177.9000 238.6000 180.2000 ;
	    RECT 239.8000 177.9000 240.2000 180.2000 ;
	    RECT 240.6000 175.9000 241.0000 180.2000 ;
	    RECT 243.0000 177.9000 243.4000 180.2000 ;
	    RECT 246.2000 175.9000 246.6000 180.2000 ;
	    RECT 248.6000 175.9000 249.0000 180.2000 ;
	    RECT 249.4000 177.9000 249.8000 180.2000 ;
	    RECT 251.0000 176.1000 251.4000 180.2000 ;
	    RECT 254.2000 175.9000 254.6000 180.2000 ;
	    RECT 255.0000 177.9000 255.4000 180.2000 ;
	    RECT 257.4000 176.0000 257.8000 180.2000 ;
	    RECT 260.2000 177.9000 260.6000 180.2000 ;
	    RECT 261.8000 177.9000 262.2000 180.2000 ;
	    RECT 264.6000 175.9000 265.0000 180.2000 ;
	    RECT 267.0000 177.9000 267.4000 180.2000 ;
	    RECT 268.6000 176.5000 269.0000 180.2000 ;
	    RECT 1.4000 160.8000 1.8000 164.5000 ;
	    RECT 3.3000 160.8000 3.7000 163.1000 ;
	    RECT 5.4000 160.8000 5.8000 165.1000 ;
	    RECT 6.2000 160.8000 6.6000 163.1000 ;
	    RECT 7.8000 160.8000 8.2000 163.1000 ;
	    RECT 9.4000 160.8000 9.8000 162.9000 ;
	    RECT 11.8000 160.8000 12.2000 164.5000 ;
	    RECT 15.8000 160.8000 16.2000 163.1000 ;
	    RECT 17.4000 160.8000 17.8000 163.1000 ;
	    RECT 18.2000 160.8000 18.6000 163.1000 ;
	    RECT 22.2000 160.8000 22.6000 164.5000 ;
	    RECT 23.8000 160.8000 24.2000 165.1000 ;
	    RECT 27.0000 160.8000 27.4000 163.1000 ;
	    RECT 27.8000 160.8000 28.2000 163.1000 ;
	    RECT 29.4000 160.8000 29.8000 162.9000 ;
	    RECT 31.0000 160.8000 31.4000 163.1000 ;
	    RECT 32.6000 160.8000 33.0000 163.1000 ;
	    RECT 34.2000 160.8000 34.6000 163.1000 ;
	    RECT 35.0000 160.8000 35.4000 165.1000 ;
	    RECT 37.1000 160.8000 37.5000 163.1000 ;
	    RECT 38.2000 160.8000 38.6000 163.1000 ;
	    RECT 39.8000 160.8000 40.2000 165.1000 ;
	    RECT 42.2000 160.8000 42.6000 162.9000 ;
	    RECT 43.8000 160.8000 44.2000 163.1000 ;
	    RECT 44.6000 160.8000 45.0000 163.1000 ;
	    RECT 48.6000 160.8000 49.0000 164.5000 ;
	    RECT 50.2000 160.8000 50.6000 165.1000 ;
	    RECT 53.4000 160.8000 53.8000 164.5000 ;
	    RECT 56.6000 160.8000 57.0000 165.1000 ;
	    RECT 59.0000 160.8000 59.4000 165.1000 ;
	    RECT 61.1000 160.8000 61.5000 163.1000 ;
	    RECT 62.2000 160.8000 62.6000 163.1000 ;
	    RECT 64.6000 160.8000 65.0000 164.5000 ;
	    RECT 68.6000 160.8000 69.0000 164.5000 ;
	    RECT 71.0000 160.8000 71.4000 163.1000 ;
	    RECT 73.4000 160.8000 73.8000 164.5000 ;
	    RECT 75.8000 160.8000 76.2000 163.1000 ;
	    RECT 77.4000 160.8000 77.8000 165.1000 ;
	    RECT 80.2000 160.8000 80.6000 163.1000 ;
	    RECT 81.8000 160.8000 82.2000 163.1000 ;
	    RECT 84.6000 160.8000 85.0000 165.0000 ;
	    RECT 87.0000 160.8000 87.4000 165.0000 ;
	    RECT 89.8000 160.8000 90.2000 163.1000 ;
	    RECT 91.4000 160.8000 91.8000 163.1000 ;
	    RECT 94.2000 160.8000 94.6000 165.1000 ;
	    RECT 95.8000 160.8000 96.2000 163.1000 ;
	    RECT 97.4000 160.8000 97.8000 165.1000 ;
	    RECT 102.2000 160.8000 102.6000 164.5000 ;
	    RECT 104.6000 160.8000 105.0000 163.1000 ;
	    RECT 107.8000 160.8000 108.2000 165.0000 ;
	    RECT 110.6000 160.8000 111.0000 163.1000 ;
	    RECT 112.2000 160.8000 112.6000 163.1000 ;
	    RECT 115.0000 160.8000 115.4000 165.1000 ;
	    RECT 116.6000 160.8000 117.0000 163.1000 ;
	    RECT 119.0000 160.8000 119.4000 164.5000 ;
	    RECT 122.2000 160.8000 122.6000 165.1000 ;
	    RECT 125.0000 160.8000 125.4000 163.1000 ;
	    RECT 126.6000 160.8000 127.0000 163.1000 ;
	    RECT 129.4000 160.8000 129.8000 165.0000 ;
	    RECT 131.0000 160.8000 131.4000 163.1000 ;
	    RECT 132.6000 160.8000 133.0000 165.1000 ;
	    RECT 136.6000 160.8000 137.0000 164.5000 ;
	    RECT 139.0000 160.8000 139.4000 163.1000 ;
	    RECT 141.4000 160.8000 141.8000 165.1000 ;
	    RECT 143.0000 160.8000 143.4000 163.1000 ;
	    RECT 144.6000 160.8000 145.0000 165.1000 ;
	    RECT 147.4000 160.8000 147.8000 163.1000 ;
	    RECT 149.0000 160.8000 149.4000 163.1000 ;
	    RECT 151.8000 160.8000 152.2000 165.0000 ;
	    RECT 153.4000 160.8000 153.8000 163.1000 ;
	    RECT 155.8000 160.8000 156.2000 165.1000 ;
	    RECT 158.6000 160.8000 159.0000 163.1000 ;
	    RECT 160.2000 160.8000 160.6000 163.1000 ;
	    RECT 163.0000 160.8000 163.4000 165.0000 ;
	    RECT 166.2000 160.8000 166.6000 165.1000 ;
	    RECT 170.2000 160.8000 170.6000 165.1000 ;
	    RECT 171.8000 160.8000 172.2000 163.1000 ;
	    RECT 173.4000 160.8000 173.8000 165.0000 ;
	    RECT 176.2000 160.8000 176.6000 163.1000 ;
	    RECT 177.8000 160.8000 178.2000 163.1000 ;
	    RECT 180.6000 160.8000 181.0000 165.1000 ;
	    RECT 183.8000 160.8000 184.2000 165.1000 ;
	    RECT 185.4000 160.8000 185.8000 163.1000 ;
	    RECT 187.0000 160.8000 187.4000 165.1000 ;
	    RECT 189.8000 160.8000 190.2000 163.1000 ;
	    RECT 191.4000 160.8000 191.8000 163.1000 ;
	    RECT 194.2000 160.8000 194.6000 165.0000 ;
	    RECT 196.6000 160.8000 197.0000 165.0000 ;
	    RECT 199.4000 160.8000 199.8000 163.1000 ;
	    RECT 201.0000 160.8000 201.4000 163.1000 ;
	    RECT 203.8000 160.8000 204.2000 165.1000 ;
	    RECT 207.0000 160.8000 207.4000 164.5000 ;
	    RECT 208.6000 160.8000 209.0000 165.1000 ;
	    RECT 212.6000 160.8000 213.0000 163.1000 ;
	    RECT 214.2000 160.8000 214.6000 163.1000 ;
	    RECT 215.3000 160.8000 215.7000 163.1000 ;
	    RECT 217.4000 160.8000 217.8000 165.1000 ;
	    RECT 218.2000 160.8000 218.6000 165.1000 ;
	    RECT 220.6000 160.8000 221.0000 163.1000 ;
	    RECT 222.2000 160.8000 222.6000 163.1000 ;
	    RECT 223.0000 160.8000 223.4000 163.1000 ;
	    RECT 224.6000 160.8000 225.0000 163.1000 ;
	    RECT 225.4000 160.8000 225.8000 163.1000 ;
	    RECT 227.0000 160.8000 227.4000 165.1000 ;
	    RECT 229.4000 160.8000 229.8000 165.1000 ;
	    RECT 231.5000 160.8000 231.9000 163.1000 ;
	    RECT 232.6000 160.8000 233.0000 165.1000 ;
	    RECT 234.7000 160.8000 235.1000 163.1000 ;
	    RECT 235.8000 160.8000 236.2000 165.1000 ;
	    RECT 237.9000 160.8000 238.3000 163.1000 ;
	    RECT 239.0000 160.8000 239.4000 165.1000 ;
	    RECT 242.2000 160.8000 242.6000 165.1000 ;
	    RECT 243.8000 160.8000 244.2000 164.9000 ;
	    RECT 245.4000 160.8000 245.8000 163.1000 ;
	    RECT 246.2000 160.8000 246.6000 165.1000 ;
	    RECT 248.3000 160.8000 248.7000 163.1000 ;
	    RECT 249.4000 160.8000 249.8000 165.1000 ;
	    RECT 251.0000 160.8000 251.4000 164.5000 ;
	    RECT 252.6000 160.8000 253.0000 165.1000 ;
	    RECT 254.7000 160.8000 255.1000 163.1000 ;
	    RECT 257.4000 160.8000 257.8000 164.5000 ;
	    RECT 260.6000 160.8000 261.0000 164.5000 ;
	    RECT 263.0000 160.8000 263.5000 164.4000 ;
	    RECT 266.1000 161.1000 266.6000 164.4000 ;
	    RECT 266.1000 160.8000 266.5000 161.1000 ;
	    RECT 268.6000 160.8000 269.0000 164.5000 ;
	    RECT 270.2000 160.8000 270.6000 165.1000 ;
	    RECT 0.2000 160.2000 271.0000 160.8000 ;
	    RECT 0.6000 157.9000 1.0000 160.2000 ;
	    RECT 4.6000 156.5000 5.0000 160.2000 ;
	    RECT 7.0000 157.9000 7.4000 160.2000 ;
	    RECT 7.8000 157.9000 8.2000 160.2000 ;
	    RECT 9.4000 157.9000 9.8000 160.2000 ;
	    RECT 11.0000 157.9000 11.4000 160.2000 ;
	    RECT 11.8000 157.9000 12.2000 160.2000 ;
	    RECT 13.4000 157.9000 13.8000 160.2000 ;
	    RECT 14.2000 157.9000 14.6000 160.2000 ;
	    RECT 15.8000 158.1000 16.2000 160.2000 ;
	    RECT 19.0000 155.9000 19.4000 160.2000 ;
	    RECT 21.1000 155.9000 21.5000 160.2000 ;
	    RECT 23.0000 155.9000 23.4000 160.2000 ;
	    RECT 25.1000 157.9000 25.5000 160.2000 ;
	    RECT 26.2000 155.9000 26.6000 160.2000 ;
	    RECT 29.4000 158.1000 29.8000 160.2000 ;
	    RECT 31.0000 157.9000 31.4000 160.2000 ;
	    RECT 32.6000 156.5000 33.0000 160.2000 ;
	    RECT 36.6000 156.5000 37.0000 160.2000 ;
	    RECT 40.6000 155.9000 41.0000 160.2000 ;
	    RECT 41.4000 155.9000 41.8000 160.2000 ;
	    RECT 43.5000 157.9000 43.9000 160.2000 ;
	    RECT 45.4000 156.5000 45.8000 160.2000 ;
	    RECT 47.0000 157.9000 47.4000 160.2000 ;
	    RECT 48.6000 155.9000 49.0000 160.2000 ;
	    RECT 51.8000 155.9000 52.2000 160.2000 ;
	    RECT 54.6000 157.9000 55.0000 160.2000 ;
	    RECT 56.2000 157.9000 56.6000 160.2000 ;
	    RECT 59.0000 156.0000 59.4000 160.2000 ;
	    RECT 63.0000 156.0000 63.4000 160.2000 ;
	    RECT 65.8000 157.9000 66.2000 160.2000 ;
	    RECT 67.4000 157.9000 67.8000 160.2000 ;
	    RECT 70.2000 155.9000 70.6000 160.2000 ;
	    RECT 71.8000 155.9000 72.2000 160.2000 ;
	    RECT 73.4000 156.5000 73.8000 160.2000 ;
	    RECT 75.8000 156.5000 76.2000 160.2000 ;
	    RECT 77.4000 157.9000 77.8000 160.2000 ;
	    RECT 79.0000 155.9000 79.4000 160.2000 ;
	    RECT 81.4000 155.9000 81.8000 160.2000 ;
	    RECT 83.0000 156.5000 83.4000 160.2000 ;
	    RECT 84.9000 157.9000 85.3000 160.2000 ;
	    RECT 87.0000 155.9000 87.4000 160.2000 ;
	    RECT 89.4000 155.9000 89.8000 160.2000 ;
	    RECT 90.2000 155.9000 90.6000 160.2000 ;
	    RECT 92.3000 157.9000 92.7000 160.2000 ;
	    RECT 93.4000 157.9000 93.8000 160.2000 ;
	    RECT 95.0000 157.9000 95.4000 160.2000 ;
	    RECT 97.4000 155.9000 97.8000 160.2000 ;
	    RECT 98.2000 157.9000 98.6000 160.2000 ;
	    RECT 99.8000 157.9000 100.2000 160.2000 ;
	    RECT 101.4000 157.9000 101.8000 160.2000 ;
	    RECT 103.8000 155.9000 104.2000 160.2000 ;
	    RECT 104.9000 157.9000 105.3000 160.2000 ;
	    RECT 107.0000 155.9000 107.4000 160.2000 ;
	    RECT 107.8000 157.9000 108.2000 160.2000 ;
	    RECT 109.4000 157.9000 109.8000 160.2000 ;
	    RECT 112.6000 155.9000 113.0000 160.2000 ;
	    RECT 115.4000 157.9000 115.8000 160.2000 ;
	    RECT 117.0000 157.9000 117.4000 160.2000 ;
	    RECT 119.8000 156.0000 120.2000 160.2000 ;
	    RECT 122.2000 156.5000 122.6000 160.2000 ;
	    RECT 124.6000 156.0000 125.0000 160.2000 ;
	    RECT 127.4000 157.9000 127.8000 160.2000 ;
	    RECT 129.0000 157.9000 129.4000 160.2000 ;
	    RECT 131.8000 155.9000 132.2000 160.2000 ;
	    RECT 134.7000 155.9000 135.1000 160.2000 ;
	    RECT 138.2000 156.5000 138.6000 160.2000 ;
	    RECT 140.6000 157.9000 141.0000 160.2000 ;
	    RECT 142.2000 156.0000 142.6000 160.2000 ;
	    RECT 145.0000 157.9000 145.4000 160.2000 ;
	    RECT 146.6000 157.9000 147.0000 160.2000 ;
	    RECT 149.4000 155.9000 149.8000 160.2000 ;
	    RECT 153.4000 156.5000 153.8000 160.2000 ;
	    RECT 155.8000 156.5000 156.2000 160.2000 ;
	    RECT 159.8000 155.9000 160.2000 160.2000 ;
	    RECT 162.6000 157.9000 163.0000 160.2000 ;
	    RECT 164.2000 157.9000 164.6000 160.2000 ;
	    RECT 167.0000 156.0000 167.4000 160.2000 ;
	    RECT 170.2000 156.5000 170.6000 160.2000 ;
	    RECT 172.1000 157.9000 172.5000 160.2000 ;
	    RECT 174.2000 155.9000 174.6000 160.2000 ;
	    RECT 176.6000 155.9000 177.0000 160.2000 ;
	    RECT 177.4000 157.9000 177.8000 160.2000 ;
	    RECT 179.0000 157.9000 179.4000 160.2000 ;
	    RECT 179.8000 157.9000 180.2000 160.2000 ;
	    RECT 181.4000 157.9000 181.8000 160.2000 ;
	    RECT 182.2000 155.9000 182.6000 160.2000 ;
	    RECT 186.2000 156.5000 186.6000 160.2000 ;
	    RECT 188.1000 157.9000 188.5000 160.2000 ;
	    RECT 190.2000 155.9000 190.6000 160.2000 ;
	    RECT 192.6000 155.9000 193.0000 160.2000 ;
	    RECT 193.4000 155.9000 193.8000 160.2000 ;
	    RECT 195.5000 157.9000 195.9000 160.2000 ;
	    RECT 197.4000 156.5000 197.8000 160.2000 ;
	    RECT 199.8000 157.9000 200.2000 160.2000 ;
	    RECT 201.4000 157.9000 201.8000 160.2000 ;
	    RECT 203.0000 156.0000 203.4000 160.2000 ;
	    RECT 205.8000 157.9000 206.2000 160.2000 ;
	    RECT 207.4000 157.9000 207.8000 160.2000 ;
	    RECT 210.2000 155.9000 210.6000 160.2000 ;
	    RECT 214.2000 156.1000 214.6000 160.2000 ;
	    RECT 215.8000 157.9000 216.2000 160.2000 ;
	    RECT 216.6000 155.9000 217.0000 160.2000 ;
	    RECT 219.0000 155.9000 219.4000 160.2000 ;
	    RECT 221.1000 157.9000 221.5000 160.2000 ;
	    RECT 222.2000 155.9000 222.6000 160.2000 ;
	    RECT 224.3000 157.9000 224.7000 160.2000 ;
	    RECT 226.2000 157.9000 226.6000 160.2000 ;
	    RECT 228.6000 155.9000 229.0000 160.2000 ;
	    RECT 230.2000 156.5000 230.6000 160.2000 ;
	    RECT 231.8000 155.9000 232.2000 160.2000 ;
	    RECT 232.6000 155.9000 233.0000 160.2000 ;
	    RECT 235.8000 156.6000 236.3000 160.2000 ;
	    RECT 238.9000 159.9000 239.3000 160.2000 ;
	    RECT 238.9000 156.6000 239.4000 159.9000 ;
	    RECT 242.2000 155.9000 242.6000 160.2000 ;
	    RECT 244.6000 155.9000 245.0000 160.2000 ;
	    RECT 246.2000 156.5000 246.6000 160.2000 ;
	    RECT 248.6000 155.9000 249.0000 160.2000 ;
	    RECT 252.6000 156.5000 253.0000 160.2000 ;
	    RECT 254.2000 155.9000 254.6000 160.2000 ;
	    RECT 256.3000 157.9000 256.7000 160.2000 ;
	    RECT 259.0000 155.9000 259.4000 160.2000 ;
	    RECT 259.8000 155.9000 260.2000 160.2000 ;
	    RECT 263.0000 157.9000 263.4000 160.2000 ;
	    RECT 263.8000 157.9000 264.2000 160.2000 ;
	    RECT 265.4000 157.9000 265.8000 160.2000 ;
	    RECT 267.3000 155.9000 267.7000 160.2000 ;
	    RECT 0.6000 140.8000 1.0000 145.1000 ;
	    RECT 3.0000 140.8000 3.4000 145.1000 ;
	    RECT 5.1000 140.8000 5.5000 143.1000 ;
	    RECT 6.2000 140.8000 6.6000 145.1000 ;
	    RECT 8.3000 140.8000 8.7000 143.1000 ;
	    RECT 9.4000 140.8000 9.8000 145.1000 ;
	    RECT 12.6000 140.8000 13.0000 145.1000 ;
	    RECT 13.4000 140.8000 13.8000 143.1000 ;
	    RECT 15.8000 140.8000 16.2000 142.9000 ;
	    RECT 17.4000 140.8000 17.8000 143.1000 ;
	    RECT 18.2000 140.8000 18.6000 143.1000 ;
	    RECT 19.8000 140.8000 20.2000 143.1000 ;
	    RECT 20.6000 140.8000 21.0000 145.1000 ;
	    RECT 22.7000 140.8000 23.1000 143.1000 ;
	    RECT 24.6000 140.8000 25.0000 144.5000 ;
	    RECT 27.8000 140.8000 28.2000 144.5000 ;
	    RECT 31.0000 140.8000 31.4000 145.0000 ;
	    RECT 33.8000 140.8000 34.2000 143.1000 ;
	    RECT 35.4000 140.8000 35.8000 143.1000 ;
	    RECT 38.2000 140.8000 38.6000 145.1000 ;
	    RECT 39.8000 140.8000 40.2000 143.1000 ;
	    RECT 41.4000 140.8000 41.8000 145.1000 ;
	    RECT 44.6000 140.8000 45.0000 145.1000 ;
	    RECT 46.2000 140.8000 46.6000 143.1000 ;
	    RECT 51.8000 140.8000 52.2000 144.1000 ;
	    RECT 53.7000 140.8000 54.1000 143.1000 ;
	    RECT 55.8000 140.8000 56.2000 145.1000 ;
	    RECT 57.4000 140.8000 57.8000 143.1000 ;
	    RECT 60.6000 140.8000 61.0000 143.1000 ;
	    RECT 62.2000 140.8000 62.6000 144.5000 ;
	    RECT 65.4000 140.8000 65.8000 145.0000 ;
	    RECT 68.2000 140.8000 68.6000 143.1000 ;
	    RECT 69.8000 140.8000 70.2000 143.1000 ;
	    RECT 72.6000 140.8000 73.0000 145.1000 ;
	    RECT 75.0000 140.8000 75.4000 145.1000 ;
	    RECT 77.8000 140.8000 78.2000 143.1000 ;
	    RECT 79.4000 140.8000 79.8000 143.1000 ;
	    RECT 82.2000 140.8000 82.6000 145.0000 ;
	    RECT 83.8000 140.8000 84.2000 143.1000 ;
	    RECT 85.4000 140.8000 85.8000 143.1000 ;
	    RECT 87.0000 140.8000 87.4000 145.0000 ;
	    RECT 89.8000 140.8000 90.2000 143.1000 ;
	    RECT 91.4000 140.8000 91.8000 143.1000 ;
	    RECT 94.2000 140.8000 94.6000 145.1000 ;
	    RECT 95.8000 140.8000 96.2000 145.1000 ;
	    RECT 98.5000 140.8000 98.9000 143.1000 ;
	    RECT 100.6000 140.8000 101.0000 145.1000 ;
	    RECT 102.2000 140.8000 102.6000 143.1000 ;
	    RECT 103.0000 140.8000 103.4000 143.1000 ;
	    RECT 104.6000 140.8000 105.0000 142.9000 ;
	    RECT 106.2000 140.8000 106.6000 143.1000 ;
	    RECT 107.8000 140.8000 108.2000 143.1000 ;
	    RECT 110.2000 140.8000 110.6000 145.1000 ;
	    RECT 112.6000 140.8000 113.0000 145.1000 ;
	    RECT 115.0000 140.8000 115.4000 143.1000 ;
	    RECT 116.6000 140.8000 117.0000 143.1000 ;
	    RECT 117.4000 140.8000 117.8000 143.1000 ;
	    RECT 119.0000 140.8000 119.4000 142.9000 ;
	    RECT 121.4000 140.8000 121.8000 143.1000 ;
	    RECT 123.0000 140.8000 123.4000 145.1000 ;
	    RECT 125.8000 140.8000 126.2000 143.1000 ;
	    RECT 127.4000 140.8000 127.8000 143.1000 ;
	    RECT 130.2000 140.8000 130.6000 145.0000 ;
	    RECT 131.8000 140.8000 132.2000 145.1000 ;
	    RECT 134.2000 140.8000 134.6000 144.5000 ;
	    RECT 136.6000 140.8000 137.0000 143.1000 ;
	    RECT 139.0000 140.8000 139.4000 144.5000 ;
	    RECT 144.6000 140.8000 145.0000 144.5000 ;
	    RECT 147.0000 140.8000 147.4000 143.1000 ;
	    RECT 148.6000 140.8000 149.0000 145.1000 ;
	    RECT 151.4000 140.8000 151.8000 143.1000 ;
	    RECT 153.0000 140.8000 153.4000 143.1000 ;
	    RECT 155.8000 140.8000 156.2000 145.0000 ;
	    RECT 157.4000 140.8000 157.8000 145.1000 ;
	    RECT 159.0000 140.8000 159.4000 144.5000 ;
	    RECT 163.0000 140.8000 163.4000 145.0000 ;
	    RECT 165.8000 140.8000 166.2000 143.1000 ;
	    RECT 167.4000 140.8000 167.8000 143.1000 ;
	    RECT 170.2000 140.8000 170.6000 145.1000 ;
	    RECT 171.8000 140.8000 172.2000 143.1000 ;
	    RECT 173.4000 140.8000 173.8000 145.1000 ;
	    RECT 176.1000 140.8000 176.5000 143.1000 ;
	    RECT 178.2000 140.8000 178.6000 145.1000 ;
	    RECT 179.8000 140.8000 180.2000 144.9000 ;
	    RECT 181.4000 140.8000 181.8000 143.1000 ;
	    RECT 182.2000 140.8000 182.6000 143.1000 ;
	    RECT 185.4000 140.8000 185.8000 145.1000 ;
	    RECT 186.2000 140.8000 186.6000 145.1000 ;
	    RECT 188.6000 140.8000 189.0000 145.1000 ;
	    RECT 190.7000 140.8000 191.1000 143.1000 ;
	    RECT 191.8000 140.8000 192.2000 145.1000 ;
	    RECT 194.2000 140.8000 194.6000 145.1000 ;
	    RECT 196.3000 140.8000 196.7000 143.1000 ;
	    RECT 198.2000 140.8000 198.6000 145.1000 ;
	    RECT 201.0000 140.8000 201.4000 143.1000 ;
	    RECT 202.6000 140.8000 203.0000 143.1000 ;
	    RECT 205.4000 140.8000 205.8000 145.0000 ;
	    RECT 208.6000 140.8000 209.0000 144.5000 ;
	    RECT 210.2000 140.8000 210.6000 143.1000 ;
	    RECT 211.8000 140.8000 212.2000 143.1000 ;
	    RECT 215.0000 140.8000 215.4000 144.5000 ;
	    RECT 218.2000 140.8000 218.6000 144.5000 ;
	    RECT 220.9000 140.8000 221.3000 143.1000 ;
	    RECT 223.0000 140.8000 223.4000 145.1000 ;
	    RECT 225.4000 140.8000 225.8000 145.1000 ;
	    RECT 226.2000 140.8000 226.6000 145.1000 ;
	    RECT 230.2000 140.8000 230.6000 145.1000 ;
	    RECT 231.8000 140.8000 232.2000 144.5000 ;
	    RECT 233.4000 140.8000 233.8000 145.1000 ;
	    RECT 235.0000 140.8000 235.4000 144.5000 ;
	    RECT 236.6000 140.8000 237.0000 145.1000 ;
	    RECT 239.0000 140.8000 239.4000 145.1000 ;
	    RECT 239.8000 140.8000 240.2000 143.1000 ;
	    RECT 243.0000 140.8000 243.4000 145.1000 ;
	    RECT 243.8000 140.8000 244.2000 143.1000 ;
	    RECT 245.4000 140.8000 245.8000 142.9000 ;
	    RECT 248.6000 140.8000 249.0000 145.1000 ;
	    RECT 249.7000 140.8000 250.1000 143.1000 ;
	    RECT 251.8000 140.8000 252.2000 145.1000 ;
	    RECT 252.9000 140.8000 253.3000 143.1000 ;
	    RECT 255.0000 140.8000 255.4000 145.1000 ;
	    RECT 256.6000 140.8000 257.0000 144.9000 ;
	    RECT 258.2000 140.8000 258.6000 143.1000 ;
	    RECT 259.0000 140.8000 259.4000 145.1000 ;
	    RECT 261.7000 140.8000 262.1000 143.1000 ;
	    RECT 263.8000 140.8000 264.2000 145.1000 ;
	    RECT 266.2000 140.8000 266.6000 145.1000 ;
	    RECT 267.0000 140.8000 267.4000 143.1000 ;
	    RECT 268.6000 140.8000 269.0000 143.1000 ;
	    RECT 270.2000 140.8000 270.6000 143.1000 ;
	    RECT 0.2000 140.2000 271.0000 140.8000 ;
	    RECT 1.4000 138.1000 1.8000 140.2000 ;
	    RECT 3.0000 137.9000 3.4000 140.2000 ;
	    RECT 4.9000 135.9000 5.3000 140.2000 ;
	    RECT 7.0000 137.9000 7.4000 140.2000 ;
	    RECT 8.6000 137.9000 9.0000 140.2000 ;
	    RECT 11.0000 135.9000 11.4000 140.2000 ;
	    RECT 12.6000 135.9000 13.0000 140.2000 ;
	    RECT 13.4000 135.9000 13.8000 140.2000 ;
	    RECT 15.0000 137.9000 15.4000 140.2000 ;
	    RECT 16.6000 137.9000 17.0000 140.2000 ;
	    RECT 18.7000 135.9000 19.1000 140.2000 ;
	    RECT 20.6000 137.9000 21.0000 140.2000 ;
	    RECT 22.2000 138.1000 22.6000 140.2000 ;
	    RECT 25.4000 135.9000 25.8000 140.2000 ;
	    RECT 27.0000 136.1000 27.4000 140.2000 ;
	    RECT 28.6000 137.9000 29.0000 140.2000 ;
	    RECT 29.4000 137.9000 29.8000 140.2000 ;
	    RECT 31.0000 137.9000 31.4000 140.2000 ;
	    RECT 31.8000 135.9000 32.2000 140.2000 ;
	    RECT 33.9000 137.9000 34.3000 140.2000 ;
	    RECT 35.3000 137.9000 35.7000 140.2000 ;
	    RECT 37.4000 135.9000 37.8000 140.2000 ;
	    RECT 39.0000 137.9000 39.4000 140.2000 ;
	    RECT 40.6000 136.0000 41.0000 140.2000 ;
	    RECT 43.4000 137.9000 43.8000 140.2000 ;
	    RECT 45.0000 137.9000 45.4000 140.2000 ;
	    RECT 47.8000 135.9000 48.2000 140.2000 ;
	    RECT 49.4000 135.9000 49.8000 140.2000 ;
	    RECT 51.8000 137.9000 52.2000 140.2000 ;
	    RECT 53.4000 136.1000 53.8000 140.2000 ;
	    RECT 55.0000 135.9000 55.4000 140.2000 ;
	    RECT 58.2000 135.9000 58.6000 140.2000 ;
	    RECT 60.6000 137.9000 61.0000 140.2000 ;
	    RECT 63.0000 135.9000 63.4000 140.2000 ;
	    RECT 65.8000 137.9000 66.2000 140.2000 ;
	    RECT 67.4000 137.9000 67.8000 140.2000 ;
	    RECT 70.2000 136.0000 70.6000 140.2000 ;
	    RECT 71.8000 135.9000 72.2000 140.2000 ;
	    RECT 73.4000 136.5000 73.8000 140.2000 ;
	    RECT 75.8000 135.9000 76.2000 140.2000 ;
	    RECT 78.6000 137.9000 79.0000 140.2000 ;
	    RECT 80.2000 137.9000 80.6000 140.2000 ;
	    RECT 83.0000 136.0000 83.4000 140.2000 ;
	    RECT 84.6000 135.9000 85.0000 140.2000 ;
	    RECT 86.2000 136.5000 86.6000 140.2000 ;
	    RECT 87.8000 137.9000 88.2000 140.2000 ;
	    RECT 90.2000 136.5000 90.6000 140.2000 ;
	    RECT 91.8000 135.9000 92.2000 140.2000 ;
	    RECT 93.4000 135.9000 93.8000 140.2000 ;
	    RECT 95.0000 135.9000 95.4000 140.2000 ;
	    RECT 96.6000 135.9000 97.0000 140.2000 ;
	    RECT 98.2000 135.9000 98.6000 140.2000 ;
	    RECT 99.0000 137.9000 99.4000 140.2000 ;
	    RECT 100.6000 137.9000 101.0000 140.2000 ;
	    RECT 102.2000 137.9000 102.6000 140.2000 ;
	    RECT 107.8000 136.9000 108.2000 140.2000 ;
	    RECT 112.6000 135.9000 113.0000 140.2000 ;
	    RECT 113.4000 137.9000 113.8000 140.2000 ;
	    RECT 115.0000 136.1000 115.4000 140.2000 ;
	    RECT 118.2000 135.9000 118.6000 140.2000 ;
	    RECT 119.8000 135.9000 120.2000 140.2000 ;
	    RECT 122.6000 137.9000 123.0000 140.2000 ;
	    RECT 124.2000 137.9000 124.6000 140.2000 ;
	    RECT 127.0000 136.0000 127.4000 140.2000 ;
	    RECT 129.4000 135.9000 129.8000 140.2000 ;
	    RECT 132.2000 137.9000 132.6000 140.2000 ;
	    RECT 133.8000 137.9000 134.2000 140.2000 ;
	    RECT 136.6000 136.0000 137.0000 140.2000 ;
	    RECT 139.0000 135.9000 139.4000 140.2000 ;
	    RECT 141.8000 137.9000 142.2000 140.2000 ;
	    RECT 143.4000 137.9000 143.8000 140.2000 ;
	    RECT 146.2000 136.0000 146.6000 140.2000 ;
	    RECT 148.6000 136.5000 149.0000 140.2000 ;
	    RECT 151.0000 135.9000 151.4000 140.2000 ;
	    RECT 153.8000 137.9000 154.2000 140.2000 ;
	    RECT 155.4000 137.9000 155.8000 140.2000 ;
	    RECT 158.2000 136.0000 158.6000 140.2000 ;
	    RECT 161.4000 135.9000 161.8000 140.2000 ;
	    RECT 163.0000 135.9000 163.4000 140.2000 ;
	    RECT 164.6000 135.9000 165.0000 140.2000 ;
	    RECT 166.2000 135.9000 166.6000 140.2000 ;
	    RECT 167.8000 135.9000 168.2000 140.2000 ;
	    RECT 168.6000 135.9000 169.0000 140.2000 ;
	    RECT 170.2000 135.9000 170.6000 140.2000 ;
	    RECT 171.8000 135.9000 172.2000 140.2000 ;
	    RECT 173.4000 135.9000 173.8000 140.2000 ;
	    RECT 175.0000 135.9000 175.4000 140.2000 ;
	    RECT 175.8000 137.9000 176.2000 140.2000 ;
	    RECT 177.4000 138.1000 177.8000 140.2000 ;
	    RECT 179.8000 136.5000 180.2000 140.2000 ;
	    RECT 181.4000 135.9000 181.8000 140.2000 ;
	    RECT 183.0000 136.5000 183.4000 140.2000 ;
	    RECT 184.6000 135.9000 185.0000 140.2000 ;
	    RECT 186.2000 136.5000 186.6000 140.2000 ;
	    RECT 187.8000 135.9000 188.2000 140.2000 ;
	    RECT 189.4000 136.5000 189.8000 140.2000 ;
	    RECT 191.0000 135.9000 191.4000 140.2000 ;
	    RECT 191.8000 135.9000 192.2000 140.2000 ;
	    RECT 193.4000 135.9000 193.8000 140.2000 ;
	    RECT 194.2000 135.9000 194.6000 140.2000 ;
	    RECT 196.6000 137.9000 197.0000 140.2000 ;
	    RECT 198.2000 138.1000 198.6000 140.2000 ;
	    RECT 200.6000 137.9000 201.0000 140.2000 ;
	    RECT 201.4000 137.9000 201.8000 140.2000 ;
	    RECT 203.0000 137.9000 203.4000 140.2000 ;
	    RECT 203.8000 137.9000 204.2000 140.2000 ;
	    RECT 207.0000 135.9000 207.4000 140.2000 ;
	    RECT 208.1000 137.9000 208.5000 140.2000 ;
	    RECT 210.2000 135.9000 210.6000 140.2000 ;
	    RECT 214.2000 136.5000 214.6000 140.2000 ;
	    RECT 215.8000 137.9000 216.2000 140.2000 ;
	    RECT 217.4000 137.9000 217.8000 140.2000 ;
	    RECT 218.2000 137.9000 218.6000 140.2000 ;
	    RECT 219.8000 137.9000 220.2000 140.2000 ;
	    RECT 220.6000 137.9000 221.0000 140.2000 ;
	    RECT 222.2000 137.9000 222.6000 140.2000 ;
	    RECT 223.8000 137.9000 224.2000 140.2000 ;
	    RECT 224.6000 137.9000 225.0000 140.2000 ;
	    RECT 226.2000 137.9000 226.6000 140.2000 ;
	    RECT 227.0000 137.9000 227.4000 140.2000 ;
	    RECT 228.6000 137.9000 229.0000 140.2000 ;
	    RECT 229.4000 137.9000 229.8000 140.2000 ;
	    RECT 231.0000 137.9000 231.4000 140.2000 ;
	    RECT 231.8000 137.9000 232.2000 140.2000 ;
	    RECT 233.4000 137.9000 233.8000 140.2000 ;
	    RECT 234.2000 137.9000 234.6000 140.2000 ;
	    RECT 235.8000 137.9000 236.2000 140.2000 ;
	    RECT 236.6000 135.9000 237.0000 140.2000 ;
	    RECT 239.0000 135.9000 239.4000 140.2000 ;
	    RECT 243.0000 135.9000 243.4000 140.2000 ;
	    RECT 244.1000 137.9000 244.5000 140.2000 ;
	    RECT 246.2000 135.9000 246.6000 140.2000 ;
	    RECT 247.0000 135.9000 247.4000 140.2000 ;
	    RECT 249.1000 137.9000 249.5000 140.2000 ;
	    RECT 250.2000 135.9000 250.6000 140.2000 ;
	    RECT 253.4000 135.9000 253.8000 140.2000 ;
	    RECT 254.2000 135.9000 254.6000 140.2000 ;
	    RECT 256.3000 137.9000 256.7000 140.2000 ;
	    RECT 257.7000 137.9000 258.1000 140.2000 ;
	    RECT 259.8000 135.9000 260.2000 140.2000 ;
	    RECT 262.2000 135.9000 262.6000 140.2000 ;
	    RECT 263.8000 136.1000 264.2000 140.2000 ;
	    RECT 265.4000 137.9000 265.8000 140.2000 ;
	    RECT 267.0000 136.5000 267.4000 140.2000 ;
	    RECT 268.6000 135.9000 269.0000 140.2000 ;
	    RECT 1.4000 121.1000 1.9000 124.4000 ;
	    RECT 1.5000 120.8000 1.9000 121.1000 ;
	    RECT 4.5000 120.8000 5.0000 124.4000 ;
	    RECT 7.0000 120.8000 7.4000 124.5000 ;
	    RECT 9.4000 120.8000 9.8000 125.1000 ;
	    RECT 12.6000 120.8000 13.0000 123.1000 ;
	    RECT 14.2000 121.1000 14.7000 124.4000 ;
	    RECT 14.3000 120.8000 14.7000 121.1000 ;
	    RECT 17.3000 120.8000 17.8000 124.4000 ;
	    RECT 20.6000 120.8000 21.0000 125.1000 ;
	    RECT 22.2000 120.8000 22.6000 124.5000 ;
	    RECT 24.6000 120.8000 25.0000 123.1000 ;
	    RECT 27.8000 120.8000 28.2000 125.1000 ;
	    RECT 28.6000 120.8000 29.0000 125.1000 ;
	    RECT 30.7000 120.8000 31.1000 123.1000 ;
	    RECT 34.2000 120.8000 34.6000 124.5000 ;
	    RECT 35.8000 120.8000 36.2000 123.1000 ;
	    RECT 37.4000 120.8000 37.8000 123.1000 ;
	    RECT 39.0000 120.8000 39.4000 123.1000 ;
	    RECT 40.1000 120.8000 40.5000 123.1000 ;
	    RECT 42.2000 120.8000 42.6000 125.1000 ;
	    RECT 43.8000 120.8000 44.2000 123.1000 ;
	    RECT 45.4000 120.8000 45.8000 125.0000 ;
	    RECT 48.2000 120.8000 48.6000 123.1000 ;
	    RECT 49.8000 120.8000 50.2000 123.1000 ;
	    RECT 52.6000 120.8000 53.0000 125.1000 ;
	    RECT 54.2000 120.8000 54.6000 123.1000 ;
	    RECT 55.8000 120.8000 56.2000 124.9000 ;
	    RECT 60.1000 120.8000 60.5000 125.1000 ;
	    RECT 63.5000 120.8000 63.9000 125.1000 ;
	    RECT 65.4000 120.8000 65.8000 123.1000 ;
	    RECT 67.0000 120.8000 67.4000 124.9000 ;
	    RECT 69.4000 120.8000 69.8000 125.1000 ;
	    RECT 72.2000 120.8000 72.6000 123.1000 ;
	    RECT 73.8000 120.8000 74.2000 123.1000 ;
	    RECT 76.6000 120.8000 77.0000 125.0000 ;
	    RECT 79.8000 120.8000 80.2000 124.5000 ;
	    RECT 81.7000 120.8000 82.1000 123.1000 ;
	    RECT 83.8000 120.8000 84.2000 125.1000 ;
	    RECT 84.6000 120.8000 85.0000 125.1000 ;
	    RECT 86.2000 120.8000 86.6000 125.1000 ;
	    RECT 87.8000 120.8000 88.2000 125.1000 ;
	    RECT 89.4000 120.8000 89.8000 125.1000 ;
	    RECT 91.0000 120.8000 91.4000 125.1000 ;
	    RECT 91.8000 120.8000 92.2000 125.1000 ;
	    RECT 94.2000 120.8000 94.6000 125.1000 ;
	    RECT 95.8000 120.8000 96.2000 124.5000 ;
	    RECT 97.4000 120.8000 97.8000 123.1000 ;
	    RECT 99.0000 120.8000 99.4000 124.9000 ;
	    RECT 100.6000 120.8000 101.0000 123.1000 ;
	    RECT 102.2000 120.8000 102.6000 123.1000 ;
	    RECT 103.0000 120.8000 103.4000 125.1000 ;
	    RECT 105.1000 120.8000 105.5000 123.1000 ;
	    RECT 107.5000 120.8000 107.9000 125.1000 ;
	    RECT 111.0000 120.8000 111.4000 123.1000 ;
	    RECT 112.6000 120.8000 113.0000 123.1000 ;
	    RECT 113.4000 120.8000 113.8000 123.1000 ;
	    RECT 115.0000 120.8000 115.4000 122.9000 ;
	    RECT 117.4000 120.8000 117.8000 124.9000 ;
	    RECT 119.0000 120.8000 119.4000 123.1000 ;
	    RECT 120.6000 120.8000 121.0000 123.1000 ;
	    RECT 123.0000 120.8000 123.4000 125.1000 ;
	    RECT 123.8000 120.8000 124.2000 125.1000 ;
	    RECT 125.9000 120.8000 126.3000 123.1000 ;
	    RECT 127.0000 120.8000 127.4000 125.1000 ;
	    RECT 130.2000 120.8000 130.6000 125.0000 ;
	    RECT 133.0000 120.8000 133.4000 123.1000 ;
	    RECT 134.6000 120.8000 135.0000 123.1000 ;
	    RECT 137.4000 120.8000 137.8000 125.1000 ;
	    RECT 139.8000 120.8000 140.2000 124.5000 ;
	    RECT 142.5000 120.8000 142.9000 123.1000 ;
	    RECT 144.6000 120.8000 145.0000 125.1000 ;
	    RECT 147.0000 120.8000 147.4000 125.1000 ;
	    RECT 148.6000 120.8000 149.0000 124.5000 ;
	    RECT 151.0000 120.8000 151.4000 123.1000 ;
	    RECT 152.6000 120.8000 153.0000 123.1000 ;
	    RECT 154.2000 120.8000 154.6000 123.1000 ;
	    RECT 155.0000 120.8000 155.4000 125.1000 ;
	    RECT 157.1000 120.8000 157.5000 123.1000 ;
	    RECT 159.8000 120.8000 160.2000 125.1000 ;
	    RECT 163.0000 120.8000 163.4000 124.5000 ;
	    RECT 164.6000 120.8000 165.0000 125.1000 ;
	    RECT 166.2000 120.8000 166.6000 125.0000 ;
	    RECT 169.0000 120.8000 169.4000 123.1000 ;
	    RECT 170.6000 120.8000 171.0000 123.1000 ;
	    RECT 173.4000 120.8000 173.8000 125.1000 ;
	    RECT 175.0000 120.8000 175.4000 123.1000 ;
	    RECT 176.6000 120.8000 177.0000 123.1000 ;
	    RECT 177.4000 120.8000 177.8000 125.1000 ;
	    RECT 179.0000 120.8000 179.4000 124.5000 ;
	    RECT 180.6000 120.8000 181.0000 123.1000 ;
	    RECT 182.2000 120.8000 182.6000 123.1000 ;
	    RECT 183.0000 120.8000 183.4000 125.1000 ;
	    RECT 184.6000 120.8000 185.0000 124.5000 ;
	    RECT 186.2000 120.8000 186.6000 123.1000 ;
	    RECT 187.8000 120.8000 188.2000 123.1000 ;
	    RECT 188.6000 120.8000 189.0000 125.1000 ;
	    RECT 190.2000 120.8000 190.6000 123.1000 ;
	    RECT 191.8000 120.8000 192.2000 123.1000 ;
	    RECT 193.4000 120.8000 193.8000 122.9000 ;
	    RECT 195.0000 120.8000 195.4000 123.1000 ;
	    RECT 196.6000 120.8000 197.0000 125.1000 ;
	    RECT 199.4000 120.8000 199.8000 123.1000 ;
	    RECT 201.0000 120.8000 201.4000 123.1000 ;
	    RECT 203.8000 120.8000 204.2000 125.0000 ;
	    RECT 205.4000 120.8000 205.8000 125.1000 ;
	    RECT 207.8000 120.8000 208.2000 125.1000 ;
	    RECT 209.4000 120.8000 209.8000 125.1000 ;
	    RECT 212.6000 120.8000 213.0000 125.1000 ;
	    RECT 215.0000 120.8000 215.4000 125.1000 ;
	    RECT 219.0000 120.8000 219.4000 124.5000 ;
	    RECT 220.6000 120.8000 221.0000 125.1000 ;
	    RECT 223.0000 120.8000 223.4000 125.1000 ;
	    RECT 225.4000 120.8000 225.8000 123.1000 ;
	    RECT 227.0000 120.8000 227.4000 123.1000 ;
	    RECT 227.8000 120.8000 228.2000 125.1000 ;
	    RECT 229.4000 120.8000 229.8000 125.1000 ;
	    RECT 231.0000 120.8000 231.4000 125.1000 ;
	    RECT 232.6000 120.8000 233.0000 125.1000 ;
	    RECT 235.0000 120.8000 235.4000 125.1000 ;
	    RECT 235.8000 120.8000 236.2000 125.1000 ;
	    RECT 238.2000 120.8000 238.6000 123.1000 ;
	    RECT 239.8000 120.8000 240.2000 125.1000 ;
	    RECT 241.9000 120.8000 242.3000 123.1000 ;
	    RECT 243.0000 120.8000 243.4000 123.1000 ;
	    RECT 246.2000 120.8000 246.6000 125.1000 ;
	    RECT 247.8000 120.8000 248.2000 123.1000 ;
	    RECT 250.2000 120.8000 250.6000 125.1000 ;
	    RECT 251.0000 120.8000 251.4000 125.1000 ;
	    RECT 253.1000 120.8000 253.5000 123.1000 ;
	    RECT 255.0000 120.8000 255.4000 123.1000 ;
	    RECT 257.4000 120.8000 257.8000 124.5000 ;
	    RECT 259.0000 120.8000 259.4000 123.1000 ;
	    RECT 261.4000 120.8000 261.8000 124.5000 ;
	    RECT 265.4000 120.8000 265.8000 124.5000 ;
	    RECT 267.0000 120.8000 267.4000 123.1000 ;
	    RECT 268.6000 120.8000 269.0000 123.1000 ;
	    RECT 0.2000 120.2000 271.0000 120.8000 ;
	    RECT 0.6000 117.9000 1.0000 120.2000 ;
	    RECT 3.8000 115.9000 4.2000 120.2000 ;
	    RECT 5.4000 116.5000 5.8000 120.2000 ;
	    RECT 7.8000 115.9000 8.2000 120.2000 ;
	    RECT 11.0000 117.9000 11.4000 120.2000 ;
	    RECT 12.6000 116.6000 13.1000 120.2000 ;
	    RECT 15.7000 119.9000 16.1000 120.2000 ;
	    RECT 15.7000 116.6000 16.2000 119.9000 ;
	    RECT 17.4000 115.9000 17.8000 120.2000 ;
	    RECT 19.5000 117.9000 19.9000 120.2000 ;
	    RECT 20.6000 117.9000 21.0000 120.2000 ;
	    RECT 22.2000 117.9000 22.6000 120.2000 ;
	    RECT 23.0000 117.9000 23.4000 120.2000 ;
	    RECT 24.6000 116.1000 25.0000 120.2000 ;
	    RECT 26.2000 115.9000 26.6000 120.2000 ;
	    RECT 28.3000 117.9000 28.7000 120.2000 ;
	    RECT 29.4000 115.9000 29.8000 120.2000 ;
	    RECT 31.5000 117.9000 31.9000 120.2000 ;
	    RECT 35.0000 116.5000 35.4000 120.2000 ;
	    RECT 37.4000 116.0000 37.8000 120.2000 ;
	    RECT 40.2000 117.9000 40.6000 120.2000 ;
	    RECT 41.8000 117.9000 42.2000 120.2000 ;
	    RECT 44.6000 115.9000 45.0000 120.2000 ;
	    RECT 46.2000 117.9000 46.6000 120.2000 ;
	    RECT 47.8000 117.9000 48.2000 120.2000 ;
	    RECT 49.4000 117.9000 49.8000 120.2000 ;
	    RECT 51.0000 116.0000 51.4000 120.2000 ;
	    RECT 53.8000 117.9000 54.2000 120.2000 ;
	    RECT 55.4000 117.9000 55.8000 120.2000 ;
	    RECT 58.2000 115.9000 58.6000 120.2000 ;
	    RECT 62.5000 115.9000 62.9000 120.2000 ;
	    RECT 65.4000 116.0000 65.8000 120.2000 ;
	    RECT 68.2000 117.9000 68.6000 120.2000 ;
	    RECT 69.8000 117.9000 70.2000 120.2000 ;
	    RECT 72.6000 115.9000 73.0000 120.2000 ;
	    RECT 74.2000 117.9000 74.6000 120.2000 ;
	    RECT 75.8000 118.1000 76.2000 120.2000 ;
	    RECT 78.2000 115.9000 78.6000 120.2000 ;
	    RECT 81.0000 117.9000 81.4000 120.2000 ;
	    RECT 82.6000 117.9000 83.0000 120.2000 ;
	    RECT 85.4000 116.0000 85.8000 120.2000 ;
	    RECT 88.6000 115.9000 89.0000 120.2000 ;
	    RECT 90.2000 116.0000 90.6000 120.2000 ;
	    RECT 93.0000 117.9000 93.4000 120.2000 ;
	    RECT 94.6000 117.9000 95.0000 120.2000 ;
	    RECT 97.4000 115.9000 97.8000 120.2000 ;
	    RECT 99.8000 117.9000 100.2000 120.2000 ;
	    RECT 100.6000 117.9000 101.0000 120.2000 ;
	    RECT 104.6000 116.5000 105.0000 120.2000 ;
	    RECT 107.8000 115.9000 108.2000 120.2000 ;
	    RECT 111.0000 117.9000 111.4000 120.2000 ;
	    RECT 112.6000 117.9000 113.0000 120.2000 ;
	    RECT 113.4000 117.9000 113.8000 120.2000 ;
	    RECT 115.0000 117.9000 115.4000 120.2000 ;
	    RECT 116.6000 117.9000 117.0000 120.2000 ;
	    RECT 117.4000 117.9000 117.8000 120.2000 ;
	    RECT 119.0000 117.9000 119.4000 120.2000 ;
	    RECT 120.6000 117.9000 121.0000 120.2000 ;
	    RECT 122.2000 116.5000 122.6000 120.2000 ;
	    RECT 123.8000 115.9000 124.2000 120.2000 ;
	    RECT 126.2000 117.9000 126.6000 120.2000 ;
	    RECT 127.8000 117.9000 128.2000 120.2000 ;
	    RECT 129.4000 118.1000 129.8000 120.2000 ;
	    RECT 131.8000 117.9000 132.2000 120.2000 ;
	    RECT 132.9000 117.9000 133.3000 120.2000 ;
	    RECT 135.0000 115.9000 135.4000 120.2000 ;
	    RECT 136.6000 116.5000 137.0000 120.2000 ;
	    RECT 139.3000 117.9000 139.7000 120.2000 ;
	    RECT 141.4000 115.9000 141.8000 120.2000 ;
	    RECT 143.8000 116.5000 144.2000 120.2000 ;
	    RECT 146.2000 117.9000 146.6000 120.2000 ;
	    RECT 148.6000 116.5000 149.0000 120.2000 ;
	    RECT 150.2000 117.9000 150.6000 120.2000 ;
	    RECT 151.8000 117.9000 152.2000 120.2000 ;
	    RECT 152.6000 115.9000 153.0000 120.2000 ;
	    RECT 154.7000 117.9000 155.1000 120.2000 ;
	    RECT 155.8000 115.9000 156.2000 120.2000 ;
	    RECT 157.4000 116.5000 157.8000 120.2000 ;
	    RECT 161.4000 116.0000 161.8000 120.2000 ;
	    RECT 164.2000 117.9000 164.6000 120.2000 ;
	    RECT 165.8000 117.9000 166.2000 120.2000 ;
	    RECT 168.6000 115.9000 169.0000 120.2000 ;
	    RECT 170.2000 115.9000 170.6000 120.2000 ;
	    RECT 172.6000 116.9000 173.0000 120.2000 ;
	    RECT 179.0000 116.1000 179.4000 120.2000 ;
	    RECT 180.6000 117.9000 181.0000 120.2000 ;
	    RECT 182.2000 116.0000 182.6000 120.2000 ;
	    RECT 185.0000 117.9000 185.4000 120.2000 ;
	    RECT 186.6000 117.9000 187.0000 120.2000 ;
	    RECT 189.4000 115.9000 189.8000 120.2000 ;
	    RECT 191.8000 116.0000 192.2000 120.2000 ;
	    RECT 194.6000 117.9000 195.0000 120.2000 ;
	    RECT 196.2000 117.9000 196.6000 120.2000 ;
	    RECT 199.0000 115.9000 199.4000 120.2000 ;
	    RECT 200.6000 115.9000 201.0000 120.2000 ;
	    RECT 202.2000 115.9000 202.6000 120.2000 ;
	    RECT 203.8000 115.9000 204.2000 120.2000 ;
	    RECT 206.2000 115.9000 206.6000 120.2000 ;
	    RECT 207.0000 117.9000 207.4000 120.2000 ;
	    RECT 208.6000 117.9000 209.0000 120.2000 ;
	    RECT 209.4000 117.9000 209.8000 120.2000 ;
	    RECT 212.6000 115.9000 213.0000 120.2000 ;
	    RECT 214.7000 117.9000 215.1000 120.2000 ;
	    RECT 215.8000 117.9000 216.2000 120.2000 ;
	    RECT 219.0000 115.9000 219.4000 120.2000 ;
	    RECT 219.8000 115.9000 220.2000 120.2000 ;
	    RECT 222.5000 117.9000 222.9000 120.2000 ;
	    RECT 224.6000 115.9000 225.0000 120.2000 ;
	    RECT 225.4000 117.9000 225.8000 120.2000 ;
	    RECT 227.0000 116.1000 227.4000 120.2000 ;
	    RECT 228.6000 117.9000 229.0000 120.2000 ;
	    RECT 230.2000 117.9000 230.6000 120.2000 ;
	    RECT 232.6000 115.9000 233.0000 120.2000 ;
	    RECT 233.4000 115.9000 233.8000 120.2000 ;
	    RECT 235.8000 117.9000 236.2000 120.2000 ;
	    RECT 237.4000 117.9000 237.8000 120.2000 ;
	    RECT 238.2000 117.9000 238.6000 120.2000 ;
	    RECT 239.8000 116.1000 240.2000 120.2000 ;
	    RECT 241.4000 117.9000 241.8000 120.2000 ;
	    RECT 243.0000 117.9000 243.4000 120.2000 ;
	    RECT 243.8000 117.9000 244.2000 120.2000 ;
	    RECT 245.4000 117.9000 245.8000 120.2000 ;
	    RECT 246.2000 117.9000 246.6000 120.2000 ;
	    RECT 247.8000 117.9000 248.2000 120.2000 ;
	    RECT 248.6000 117.9000 249.0000 120.2000 ;
	    RECT 250.2000 117.9000 250.6000 120.2000 ;
	    RECT 252.6000 115.9000 253.0000 120.2000 ;
	    RECT 255.0000 115.9000 255.4000 120.2000 ;
	    RECT 257.4000 115.9000 257.8000 120.2000 ;
	    RECT 259.8000 115.9000 260.2000 120.2000 ;
	    RECT 260.6000 115.9000 261.0000 120.2000 ;
	    RECT 262.7000 117.9000 263.1000 120.2000 ;
	    RECT 263.8000 115.9000 264.2000 120.2000 ;
	    RECT 265.9000 117.9000 266.3000 120.2000 ;
	    RECT 267.0000 117.9000 267.4000 120.2000 ;
	    RECT 268.6000 117.9000 269.0000 120.2000 ;
	    RECT 0.6000 100.8000 1.0000 105.1000 ;
	    RECT 2.7000 100.8000 3.1000 103.1000 ;
	    RECT 3.8000 100.8000 4.2000 103.1000 ;
	    RECT 5.4000 100.8000 5.8000 103.1000 ;
	    RECT 7.8000 100.8000 8.2000 105.1000 ;
	    RECT 9.4000 100.8000 9.8000 104.5000 ;
	    RECT 11.8000 100.8000 12.2000 103.1000 ;
	    RECT 13.4000 100.8000 13.8000 103.1000 ;
	    RECT 15.0000 100.8000 15.5000 104.4000 ;
	    RECT 18.1000 101.1000 18.6000 104.4000 ;
	    RECT 18.1000 100.8000 18.5000 101.1000 ;
	    RECT 19.8000 100.8000 20.2000 103.1000 ;
	    RECT 21.4000 100.8000 21.8000 105.1000 ;
	    RECT 24.6000 100.8000 25.0000 105.1000 ;
	    RECT 27.4000 100.8000 27.8000 103.1000 ;
	    RECT 29.0000 100.8000 29.4000 103.1000 ;
	    RECT 31.8000 100.8000 32.2000 105.0000 ;
	    RECT 33.4000 100.8000 33.8000 103.1000 ;
	    RECT 35.0000 100.8000 35.4000 105.1000 ;
	    RECT 42.2000 100.8000 42.6000 104.1000 ;
	    RECT 44.6000 100.8000 45.0000 103.1000 ;
	    RECT 45.4000 100.8000 45.8000 105.1000 ;
	    RECT 47.8000 100.8000 48.2000 105.1000 ;
	    RECT 49.9000 100.8000 50.3000 103.1000 ;
	    RECT 52.6000 100.8000 53.0000 105.1000 ;
	    RECT 53.7000 100.8000 54.1000 103.1000 ;
	    RECT 55.8000 100.8000 56.2000 105.1000 ;
	    RECT 59.8000 100.8000 60.2000 104.5000 ;
	    RECT 62.2000 100.8000 62.6000 104.5000 ;
	    RECT 65.4000 100.8000 65.8000 102.9000 ;
	    RECT 67.0000 100.8000 67.4000 103.1000 ;
	    RECT 68.6000 100.8000 69.0000 105.1000 ;
	    RECT 71.4000 100.8000 71.8000 103.1000 ;
	    RECT 73.0000 100.8000 73.4000 103.1000 ;
	    RECT 75.8000 100.8000 76.2000 105.0000 ;
	    RECT 79.0000 100.8000 79.4000 104.5000 ;
	    RECT 80.9000 100.8000 81.3000 103.1000 ;
	    RECT 83.0000 100.8000 83.4000 105.1000 ;
	    RECT 85.4000 100.8000 85.8000 104.5000 ;
	    RECT 87.3000 100.8000 87.7000 103.1000 ;
	    RECT 89.4000 100.8000 89.8000 105.1000 ;
	    RECT 90.2000 100.8000 90.6000 103.1000 ;
	    RECT 91.8000 100.8000 92.2000 103.1000 ;
	    RECT 93.4000 100.8000 93.8000 103.1000 ;
	    RECT 95.0000 100.8000 95.4000 102.9000 ;
	    RECT 96.6000 100.8000 97.0000 103.1000 ;
	    RECT 99.0000 100.8000 99.4000 105.1000 ;
	    RECT 101.1000 100.8000 101.5000 105.1000 ;
	    RECT 103.0000 100.8000 103.4000 105.1000 ;
	    RECT 105.1000 100.8000 105.5000 103.1000 ;
	    RECT 107.0000 100.8000 107.4000 102.9000 ;
	    RECT 108.6000 100.8000 109.0000 103.1000 ;
	    RECT 113.4000 100.8000 113.8000 104.5000 ;
	    RECT 115.8000 100.8000 116.2000 104.5000 ;
	    RECT 119.8000 100.8000 120.2000 105.1000 ;
	    RECT 120.9000 100.8000 121.3000 103.1000 ;
	    RECT 123.0000 100.8000 123.4000 105.1000 ;
	    RECT 124.6000 100.8000 125.0000 105.1000 ;
	    RECT 127.4000 100.8000 127.8000 103.1000 ;
	    RECT 129.0000 100.8000 129.4000 103.1000 ;
	    RECT 131.8000 100.8000 132.2000 105.0000 ;
	    RECT 134.2000 100.8000 134.6000 105.1000 ;
	    RECT 137.0000 100.8000 137.4000 103.1000 ;
	    RECT 138.6000 100.8000 139.0000 103.1000 ;
	    RECT 141.4000 100.8000 141.8000 105.0000 ;
	    RECT 144.6000 100.8000 145.0000 105.1000 ;
	    RECT 150.2000 100.8000 150.6000 104.1000 ;
	    RECT 152.6000 100.8000 153.0000 104.9000 ;
	    RECT 154.2000 100.8000 154.6000 103.1000 ;
	    RECT 156.3000 100.8000 156.7000 105.1000 ;
	    RECT 159.0000 100.8000 159.4000 104.5000 ;
	    RECT 163.8000 100.8000 164.2000 103.1000 ;
	    RECT 165.4000 100.8000 165.8000 102.9000 ;
	    RECT 167.0000 100.8000 167.4000 103.1000 ;
	    RECT 167.8000 100.8000 168.2000 103.1000 ;
	    RECT 169.4000 100.8000 169.8000 104.9000 ;
	    RECT 171.0000 100.8000 171.4000 103.1000 ;
	    RECT 172.6000 100.8000 173.0000 102.9000 ;
	    RECT 174.2000 100.8000 174.6000 105.1000 ;
	    RECT 176.6000 100.8000 177.0000 102.9000 ;
	    RECT 178.2000 100.8000 178.6000 103.1000 ;
	    RECT 180.6000 100.8000 181.0000 104.5000 ;
	    RECT 182.2000 100.8000 182.6000 105.1000 ;
	    RECT 184.3000 100.8000 184.7000 103.1000 ;
	    RECT 186.2000 100.8000 186.7000 104.4000 ;
	    RECT 189.3000 101.1000 189.8000 104.4000 ;
	    RECT 189.3000 100.8000 189.7000 101.1000 ;
	    RECT 192.6000 100.8000 193.0000 104.5000 ;
	    RECT 194.2000 100.8000 194.6000 105.1000 ;
	    RECT 196.3000 100.8000 196.7000 103.1000 ;
	    RECT 198.2000 100.8000 198.7000 104.4000 ;
	    RECT 201.3000 101.1000 201.8000 104.4000 ;
	    RECT 201.3000 100.8000 201.7000 101.1000 ;
	    RECT 203.0000 100.8000 203.4000 103.1000 ;
	    RECT 204.6000 100.8000 205.0000 103.1000 ;
	    RECT 205.4000 100.8000 205.8000 105.1000 ;
	    RECT 207.5000 100.8000 207.9000 103.1000 ;
	    RECT 210.2000 100.8000 210.6000 104.5000 ;
	    RECT 213.7000 100.8000 214.1000 103.1000 ;
	    RECT 215.8000 100.8000 216.2000 105.1000 ;
	    RECT 217.4000 100.8000 217.8000 104.9000 ;
	    RECT 220.0000 100.8000 220.4000 105.1000 ;
	    RECT 222.2000 100.8000 222.6000 103.1000 ;
	    RECT 223.3000 100.8000 223.7000 103.1000 ;
	    RECT 225.4000 100.8000 225.8000 105.1000 ;
	    RECT 226.2000 100.8000 226.6000 103.1000 ;
	    RECT 227.8000 100.8000 228.2000 104.9000 ;
	    RECT 229.4000 100.8000 229.8000 105.1000 ;
	    RECT 231.0000 100.8000 231.4000 104.5000 ;
	    RECT 232.6000 100.8000 233.0000 105.1000 ;
	    RECT 235.0000 100.8000 235.4000 105.1000 ;
	    RECT 239.0000 100.8000 239.4000 105.1000 ;
	    RECT 239.8000 100.8000 240.2000 103.1000 ;
	    RECT 242.2000 101.1000 242.7000 104.4000 ;
	    RECT 242.3000 100.8000 242.7000 101.1000 ;
	    RECT 245.3000 100.8000 245.8000 104.4000 ;
	    RECT 248.6000 100.8000 249.0000 105.1000 ;
	    RECT 251.0000 100.8000 251.4000 104.5000 ;
	    RECT 252.6000 100.8000 253.0000 105.1000 ;
	    RECT 254.7000 100.8000 255.1000 103.1000 ;
	    RECT 256.6000 101.1000 257.1000 104.4000 ;
	    RECT 256.7000 100.8000 257.1000 101.1000 ;
	    RECT 259.7000 100.8000 260.2000 104.4000 ;
	    RECT 261.7000 100.8000 262.1000 103.1000 ;
	    RECT 263.8000 100.8000 264.2000 105.1000 ;
	    RECT 264.9000 100.8000 265.3000 103.1000 ;
	    RECT 267.0000 100.8000 267.4000 105.1000 ;
	    RECT 268.6000 100.8000 269.0000 103.1000 ;
	    RECT 0.2000 100.2000 271.0000 100.8000 ;
	    RECT 0.6000 97.9000 1.0000 100.2000 ;
	    RECT 2.2000 95.9000 2.6000 100.2000 ;
	    RECT 5.4000 95.9000 5.8000 100.2000 ;
	    RECT 6.2000 97.9000 6.6000 100.2000 ;
	    RECT 10.2000 96.5000 10.6000 100.2000 ;
	    RECT 11.8000 97.9000 12.2000 100.2000 ;
	    RECT 13.4000 97.9000 13.8000 100.2000 ;
	    RECT 14.2000 97.9000 14.6000 100.2000 ;
	    RECT 15.8000 96.1000 16.2000 100.2000 ;
	    RECT 18.2000 96.6000 18.7000 100.2000 ;
	    RECT 21.3000 99.9000 21.7000 100.2000 ;
	    RECT 21.3000 96.6000 21.8000 99.9000 ;
	    RECT 23.0000 95.9000 23.4000 100.2000 ;
	    RECT 25.1000 97.9000 25.5000 100.2000 ;
	    RECT 26.2000 97.9000 26.6000 100.2000 ;
	    RECT 27.8000 97.9000 28.2000 100.2000 ;
	    RECT 29.4000 96.5000 29.8000 100.2000 ;
	    RECT 31.8000 95.9000 32.2000 100.2000 ;
	    RECT 35.0000 97.9000 35.4000 100.2000 ;
	    RECT 35.8000 97.9000 36.2000 100.2000 ;
	    RECT 38.2000 96.6000 38.7000 100.2000 ;
	    RECT 41.3000 99.9000 41.7000 100.2000 ;
	    RECT 41.3000 96.6000 41.8000 99.9000 ;
	    RECT 44.6000 95.9000 45.0000 100.2000 ;
	    RECT 46.2000 97.9000 46.6000 100.2000 ;
	    RECT 48.6000 96.5000 49.0000 100.2000 ;
	    RECT 50.2000 95.9000 50.6000 100.2000 ;
	    RECT 52.9000 97.9000 53.3000 100.2000 ;
	    RECT 55.0000 95.9000 55.4000 100.2000 ;
	    RECT 55.8000 97.9000 56.2000 100.2000 ;
	    RECT 60.6000 96.5000 61.0000 100.2000 ;
	    RECT 63.0000 96.0000 63.4000 100.2000 ;
	    RECT 65.8000 97.9000 66.2000 100.2000 ;
	    RECT 67.4000 97.9000 67.8000 100.2000 ;
	    RECT 70.2000 95.9000 70.6000 100.2000 ;
	    RECT 71.8000 97.9000 72.2000 100.2000 ;
	    RECT 73.4000 98.1000 73.8000 100.2000 ;
	    RECT 75.0000 95.9000 75.4000 100.2000 ;
	    RECT 77.4000 97.9000 77.8000 100.2000 ;
	    RECT 79.0000 97.9000 79.4000 100.2000 ;
	    RECT 80.6000 98.1000 81.0000 100.2000 ;
	    RECT 82.2000 97.9000 82.6000 100.2000 ;
	    RECT 83.8000 98.1000 84.2000 100.2000 ;
	    RECT 85.4000 97.9000 85.8000 100.2000 ;
	    RECT 86.2000 95.9000 86.6000 100.2000 ;
	    RECT 87.8000 96.5000 88.2000 100.2000 ;
	    RECT 89.4000 95.9000 89.8000 100.2000 ;
	    RECT 91.0000 96.5000 91.4000 100.2000 ;
	    RECT 92.6000 95.9000 93.0000 100.2000 ;
	    RECT 94.2000 96.5000 94.6000 100.2000 ;
	    RECT 96.1000 97.9000 96.5000 100.2000 ;
	    RECT 98.2000 95.9000 98.6000 100.2000 ;
	    RECT 100.6000 96.5000 101.0000 100.2000 ;
	    RECT 103.0000 97.9000 103.4000 100.2000 ;
	    RECT 104.6000 96.0000 105.0000 100.2000 ;
	    RECT 107.4000 97.9000 107.8000 100.2000 ;
	    RECT 109.0000 97.9000 109.4000 100.2000 ;
	    RECT 111.8000 95.9000 112.2000 100.2000 ;
	    RECT 115.8000 96.0000 116.2000 100.2000 ;
	    RECT 118.6000 97.9000 119.0000 100.2000 ;
	    RECT 120.2000 97.9000 120.6000 100.2000 ;
	    RECT 123.0000 95.9000 123.4000 100.2000 ;
	    RECT 125.4000 95.9000 125.8000 100.2000 ;
	    RECT 126.2000 97.9000 126.6000 100.2000 ;
	    RECT 128.6000 95.9000 129.0000 100.2000 ;
	    RECT 131.4000 97.9000 131.8000 100.2000 ;
	    RECT 133.0000 97.9000 133.4000 100.2000 ;
	    RECT 135.8000 96.0000 136.2000 100.2000 ;
	    RECT 138.2000 96.5000 138.6000 100.2000 ;
	    RECT 140.9000 97.9000 141.3000 100.2000 ;
	    RECT 143.0000 95.9000 143.4000 100.2000 ;
	    RECT 143.8000 95.9000 144.2000 100.2000 ;
	    RECT 145.9000 97.9000 146.3000 100.2000 ;
	    RECT 147.0000 95.9000 147.4000 100.2000 ;
	    RECT 148.6000 95.9000 149.0000 100.2000 ;
	    RECT 150.2000 95.9000 150.6000 100.2000 ;
	    RECT 151.8000 95.9000 152.2000 100.2000 ;
	    RECT 153.4000 95.9000 153.8000 100.2000 ;
	    RECT 155.0000 96.0000 155.4000 100.2000 ;
	    RECT 157.8000 97.9000 158.2000 100.2000 ;
	    RECT 159.4000 97.9000 159.8000 100.2000 ;
	    RECT 162.2000 95.9000 162.6000 100.2000 ;
	    RECT 167.0000 96.5000 167.4000 100.2000 ;
	    RECT 168.6000 97.9000 169.0000 100.2000 ;
	    RECT 170.2000 97.9000 170.6000 100.2000 ;
	    RECT 171.8000 96.5000 172.2000 100.2000 ;
	    RECT 175.0000 96.0000 175.4000 100.2000 ;
	    RECT 177.8000 97.9000 178.2000 100.2000 ;
	    RECT 179.4000 97.9000 179.8000 100.2000 ;
	    RECT 182.2000 95.9000 182.6000 100.2000 ;
	    RECT 183.8000 97.9000 184.2000 100.2000 ;
	    RECT 185.4000 97.9000 185.8000 100.2000 ;
	    RECT 186.2000 95.9000 186.6000 100.2000 ;
	    RECT 188.3000 97.9000 188.7000 100.2000 ;
	    RECT 190.2000 97.9000 190.6000 100.2000 ;
	    RECT 191.8000 96.0000 192.2000 100.2000 ;
	    RECT 194.6000 97.9000 195.0000 100.2000 ;
	    RECT 196.2000 97.9000 196.6000 100.2000 ;
	    RECT 199.0000 95.9000 199.4000 100.2000 ;
	    RECT 202.2000 96.5000 202.6000 100.2000 ;
	    RECT 204.1000 97.9000 204.5000 100.2000 ;
	    RECT 206.2000 95.9000 206.6000 100.2000 ;
	    RECT 207.0000 97.9000 207.4000 100.2000 ;
	    RECT 208.6000 97.9000 209.0000 100.2000 ;
	    RECT 211.0000 95.9000 211.4000 100.2000 ;
	    RECT 213.4000 97.9000 213.8000 100.2000 ;
	    RECT 215.0000 97.9000 215.4000 100.2000 ;
	    RECT 216.7000 99.9000 217.1000 100.2000 ;
	    RECT 216.6000 96.6000 217.1000 99.9000 ;
	    RECT 219.7000 96.6000 220.2000 100.2000 ;
	    RECT 223.0000 95.9000 223.4000 100.2000 ;
	    RECT 224.6000 96.5000 225.0000 100.2000 ;
	    RECT 226.2000 95.9000 226.6000 100.2000 ;
	    RECT 227.8000 97.9000 228.2000 100.2000 ;
	    RECT 228.6000 97.9000 229.0000 100.2000 ;
	    RECT 230.2000 97.9000 230.6000 100.2000 ;
	    RECT 231.0000 97.9000 231.4000 100.2000 ;
	    RECT 232.6000 97.9000 233.0000 100.2000 ;
	    RECT 234.2000 96.5000 234.6000 100.2000 ;
	    RECT 235.8000 95.9000 236.2000 100.2000 ;
	    RECT 237.7000 95.9000 238.1000 100.2000 ;
	    RECT 239.8000 97.9000 240.2000 100.2000 ;
	    RECT 241.4000 97.9000 241.8000 100.2000 ;
	    RECT 242.2000 95.9000 242.6000 100.2000 ;
	    RECT 246.2000 95.9000 246.6000 100.2000 ;
	    RECT 247.0000 95.9000 247.4000 100.2000 ;
	    RECT 250.2000 96.1000 250.6000 100.2000 ;
	    RECT 252.8000 95.9000 253.2000 100.2000 ;
	    RECT 254.2000 95.9000 254.6000 100.2000 ;
	    RECT 257.5000 99.9000 257.9000 100.2000 ;
	    RECT 257.4000 96.6000 257.9000 99.9000 ;
	    RECT 260.5000 96.6000 261.0000 100.2000 ;
	    RECT 263.0000 96.6000 263.5000 100.2000 ;
	    RECT 266.1000 99.9000 266.5000 100.2000 ;
	    RECT 266.1000 96.6000 266.6000 99.9000 ;
	    RECT 269.4000 95.9000 269.8000 100.2000 ;
	    RECT 0.9000 80.8000 1.3000 83.1000 ;
	    RECT 3.0000 80.8000 3.4000 85.1000 ;
	    RECT 4.6000 80.8000 5.0000 83.1000 ;
	    RECT 6.2000 80.8000 6.6000 84.5000 ;
	    RECT 10.2000 80.8000 10.6000 83.1000 ;
	    RECT 11.8000 81.1000 12.3000 84.4000 ;
	    RECT 11.9000 80.8000 12.3000 81.1000 ;
	    RECT 14.9000 80.8000 15.4000 84.4000 ;
	    RECT 16.6000 80.8000 17.0000 83.1000 ;
	    RECT 18.2000 80.8000 18.6000 83.1000 ;
	    RECT 19.0000 80.8000 19.4000 85.1000 ;
	    RECT 22.2000 81.1000 22.7000 84.4000 ;
	    RECT 22.3000 80.8000 22.7000 81.1000 ;
	    RECT 25.3000 80.8000 25.8000 84.4000 ;
	    RECT 27.8000 80.8000 28.3000 84.4000 ;
	    RECT 30.9000 81.1000 31.4000 84.4000 ;
	    RECT 33.4000 81.1000 33.9000 84.4000 ;
	    RECT 30.9000 80.8000 31.3000 81.1000 ;
	    RECT 33.5000 80.8000 33.9000 81.1000 ;
	    RECT 36.5000 80.8000 37.0000 84.4000 ;
	    RECT 39.0000 80.8000 39.4000 85.1000 ;
	    RECT 41.8000 80.8000 42.2000 83.1000 ;
	    RECT 43.4000 80.8000 43.8000 83.1000 ;
	    RECT 46.2000 80.8000 46.6000 85.0000 ;
	    RECT 49.4000 80.8000 49.8000 85.1000 ;
	    RECT 51.0000 80.8000 51.4000 82.9000 ;
	    RECT 52.6000 80.8000 53.0000 83.1000 ;
	    RECT 54.5000 80.8000 54.9000 85.1000 ;
	    RECT 56.6000 80.8000 57.0000 83.1000 ;
	    RECT 58.2000 80.8000 58.6000 83.1000 ;
	    RECT 60.9000 80.8000 61.3000 83.1000 ;
	    RECT 63.0000 80.8000 63.4000 85.1000 ;
	    RECT 64.6000 80.8000 65.0000 82.9000 ;
	    RECT 66.2000 80.8000 66.6000 83.1000 ;
	    RECT 67.8000 80.8000 68.2000 85.1000 ;
	    RECT 70.6000 80.8000 71.0000 83.1000 ;
	    RECT 72.2000 80.8000 72.6000 83.1000 ;
	    RECT 75.0000 80.8000 75.4000 85.0000 ;
	    RECT 76.6000 80.8000 77.0000 85.1000 ;
	    RECT 79.8000 80.8000 80.2000 85.0000 ;
	    RECT 82.6000 80.8000 83.0000 83.1000 ;
	    RECT 84.2000 80.8000 84.6000 83.1000 ;
	    RECT 87.0000 80.8000 87.4000 85.1000 ;
	    RECT 89.4000 80.8000 89.8000 85.1000 ;
	    RECT 92.2000 80.8000 92.6000 83.1000 ;
	    RECT 93.8000 80.8000 94.2000 83.1000 ;
	    RECT 96.6000 80.8000 97.0000 85.0000 ;
	    RECT 98.2000 80.8000 98.6000 85.1000 ;
	    RECT 100.3000 80.8000 100.7000 83.1000 ;
	    RECT 101.4000 80.8000 101.8000 85.1000 ;
	    RECT 103.0000 80.8000 103.4000 84.5000 ;
	    RECT 104.6000 80.8000 105.0000 85.1000 ;
	    RECT 106.2000 80.8000 106.6000 85.1000 ;
	    RECT 107.8000 80.8000 108.2000 85.1000 ;
	    RECT 111.8000 80.8000 112.2000 84.5000 ;
	    RECT 113.4000 80.8000 113.8000 83.1000 ;
	    RECT 115.0000 80.8000 115.4000 82.9000 ;
	    RECT 116.6000 80.8000 117.0000 83.1000 ;
	    RECT 118.2000 80.8000 118.6000 83.1000 ;
	    RECT 119.8000 80.8000 120.2000 83.1000 ;
	    RECT 121.4000 80.8000 121.8000 85.1000 ;
	    RECT 124.2000 80.8000 124.6000 83.1000 ;
	    RECT 125.8000 80.8000 126.2000 83.1000 ;
	    RECT 128.6000 80.8000 129.0000 85.0000 ;
	    RECT 130.2000 80.8000 130.6000 85.1000 ;
	    RECT 132.6000 80.8000 133.0000 83.1000 ;
	    RECT 134.2000 80.8000 134.6000 85.1000 ;
	    RECT 137.4000 80.8000 137.8000 85.0000 ;
	    RECT 140.2000 80.8000 140.6000 83.1000 ;
	    RECT 141.8000 80.8000 142.2000 83.1000 ;
	    RECT 144.6000 80.8000 145.0000 85.1000 ;
	    RECT 147.0000 80.8000 147.4000 85.1000 ;
	    RECT 149.8000 80.8000 150.2000 83.1000 ;
	    RECT 151.4000 80.8000 151.8000 83.1000 ;
	    RECT 154.2000 80.8000 154.6000 85.0000 ;
	    RECT 155.8000 80.8000 156.2000 83.1000 ;
	    RECT 157.4000 80.8000 157.8000 83.1000 ;
	    RECT 158.5000 80.8000 158.9000 83.1000 ;
	    RECT 160.6000 80.8000 161.0000 85.1000 ;
	    RECT 164.6000 80.8000 165.0000 84.5000 ;
	    RECT 166.2000 80.8000 166.6000 83.1000 ;
	    RECT 167.8000 80.8000 168.2000 83.1000 ;
	    RECT 169.4000 80.8000 169.8000 83.1000 ;
	    RECT 170.2000 80.8000 170.6000 83.1000 ;
	    RECT 171.8000 80.8000 172.2000 83.1000 ;
	    RECT 173.4000 80.8000 173.8000 85.0000 ;
	    RECT 176.2000 80.8000 176.6000 83.1000 ;
	    RECT 177.8000 80.8000 178.2000 83.1000 ;
	    RECT 180.6000 80.8000 181.0000 85.1000 ;
	    RECT 183.0000 80.8000 183.4000 83.1000 ;
	    RECT 183.8000 80.8000 184.2000 85.1000 ;
	    RECT 186.2000 80.8000 186.6000 83.1000 ;
	    RECT 187.8000 80.8000 188.2000 83.1000 ;
	    RECT 190.2000 80.8000 190.6000 84.5000 ;
	    RECT 193.4000 80.8000 193.8000 85.1000 ;
	    RECT 195.0000 80.8000 195.4000 82.9000 ;
	    RECT 196.6000 80.8000 197.0000 83.1000 ;
	    RECT 197.4000 80.8000 197.8000 83.1000 ;
	    RECT 200.6000 80.8000 201.0000 85.1000 ;
	    RECT 201.4000 80.8000 201.8000 85.1000 ;
	    RECT 203.5000 80.8000 203.9000 83.1000 ;
	    RECT 204.6000 80.8000 205.0000 83.1000 ;
	    RECT 206.2000 80.8000 206.6000 83.1000 ;
	    RECT 207.0000 80.8000 207.4000 85.1000 ;
	    RECT 209.4000 80.8000 209.8000 83.1000 ;
	    RECT 212.6000 80.8000 213.0000 85.1000 ;
	    RECT 214.7000 80.8000 215.1000 83.1000 ;
	    RECT 216.1000 80.8000 216.5000 83.1000 ;
	    RECT 218.2000 80.8000 218.6000 85.1000 ;
	    RECT 220.6000 80.8000 221.0000 84.5000 ;
	    RECT 222.2000 80.8000 222.6000 85.1000 ;
	    RECT 224.3000 80.8000 224.7000 83.1000 ;
	    RECT 225.4000 80.8000 225.8000 85.1000 ;
	    RECT 227.5000 80.8000 227.9000 83.1000 ;
	    RECT 229.4000 80.8000 229.8000 83.1000 ;
	    RECT 231.0000 80.8000 231.4000 83.1000 ;
	    RECT 232.6000 81.1000 233.1000 84.4000 ;
	    RECT 232.7000 80.8000 233.1000 81.1000 ;
	    RECT 235.7000 80.8000 236.2000 84.4000 ;
	    RECT 237.4000 80.8000 237.8000 83.1000 ;
	    RECT 239.0000 80.8000 239.4000 85.1000 ;
	    RECT 240.6000 80.8000 241.0000 85.1000 ;
	    RECT 241.4000 80.8000 241.8000 83.1000 ;
	    RECT 243.0000 80.8000 243.4000 85.1000 ;
	    RECT 245.1000 80.8000 245.5000 83.1000 ;
	    RECT 246.2000 80.8000 246.6000 85.1000 ;
	    RECT 248.3000 80.8000 248.7000 83.1000 ;
	    RECT 251.0000 80.8000 251.4000 85.1000 ;
	    RECT 251.8000 80.8000 252.2000 85.1000 ;
	    RECT 253.9000 80.8000 254.3000 83.1000 ;
	    RECT 255.0000 80.8000 255.4000 85.1000 ;
	    RECT 257.1000 80.8000 257.5000 83.1000 ;
	    RECT 259.0000 81.1000 259.5000 84.4000 ;
	    RECT 259.1000 80.8000 259.5000 81.1000 ;
	    RECT 262.1000 80.8000 262.6000 84.4000 ;
	    RECT 264.6000 80.8000 265.1000 84.4000 ;
	    RECT 267.7000 81.1000 268.2000 84.4000 ;
	    RECT 267.7000 80.8000 268.1000 81.1000 ;
	    RECT 0.2000 80.2000 271.0000 80.8000 ;
	    RECT 0.6000 77.9000 1.0000 80.2000 ;
	    RECT 4.6000 76.5000 5.0000 80.2000 ;
	    RECT 6.2000 75.9000 6.6000 80.2000 ;
	    RECT 9.4000 75.9000 9.8000 80.2000 ;
	    RECT 11.0000 77.9000 11.4000 80.2000 ;
	    RECT 11.8000 77.9000 12.2000 80.2000 ;
	    RECT 15.8000 76.5000 16.2000 80.2000 ;
	    RECT 17.7000 77.9000 18.1000 80.2000 ;
	    RECT 19.8000 75.9000 20.2000 80.2000 ;
	    RECT 21.4000 77.9000 21.8000 80.2000 ;
	    RECT 22.2000 77.9000 22.6000 80.2000 ;
	    RECT 23.8000 77.9000 24.2000 80.2000 ;
	    RECT 24.6000 77.9000 25.0000 80.2000 ;
	    RECT 26.2000 76.1000 26.6000 80.2000 ;
	    RECT 27.8000 75.9000 28.2000 80.2000 ;
	    RECT 29.9000 77.9000 30.3000 80.2000 ;
	    RECT 31.0000 77.9000 31.4000 80.2000 ;
	    RECT 32.6000 77.9000 33.0000 80.2000 ;
	    RECT 33.4000 75.9000 33.8000 80.2000 ;
	    RECT 36.6000 76.6000 37.1000 80.2000 ;
	    RECT 39.7000 79.9000 40.1000 80.2000 ;
	    RECT 39.7000 76.6000 40.2000 79.9000 ;
	    RECT 41.4000 77.9000 41.8000 80.2000 ;
	    RECT 43.3000 77.9000 43.7000 80.2000 ;
	    RECT 45.4000 75.9000 45.8000 80.2000 ;
	    RECT 47.0000 76.5000 47.4000 80.2000 ;
	    RECT 51.0000 77.9000 51.4000 80.2000 ;
	    RECT 51.8000 75.9000 52.2000 80.2000 ;
	    RECT 53.9000 77.9000 54.3000 80.2000 ;
	    RECT 55.0000 77.9000 55.4000 80.2000 ;
	    RECT 56.6000 78.1000 57.0000 80.2000 ;
	    RECT 60.6000 75.9000 61.0000 80.2000 ;
	    RECT 63.4000 77.9000 63.8000 80.2000 ;
	    RECT 65.0000 77.9000 65.4000 80.2000 ;
	    RECT 67.8000 76.0000 68.2000 80.2000 ;
	    RECT 71.0000 76.5000 71.4000 80.2000 ;
	    RECT 72.9000 77.9000 73.3000 80.2000 ;
	    RECT 75.0000 75.9000 75.4000 80.2000 ;
	    RECT 76.1000 77.9000 76.5000 80.2000 ;
	    RECT 78.2000 75.9000 78.6000 80.2000 ;
	    RECT 79.8000 75.9000 80.2000 80.2000 ;
	    RECT 82.6000 77.9000 83.0000 80.2000 ;
	    RECT 84.2000 77.9000 84.6000 80.2000 ;
	    RECT 87.0000 76.0000 87.4000 80.2000 ;
	    RECT 89.4000 77.9000 89.8000 80.2000 ;
	    RECT 90.2000 77.9000 90.6000 80.2000 ;
	    RECT 91.8000 77.9000 92.2000 80.2000 ;
	    RECT 92.6000 75.9000 93.0000 80.2000 ;
	    RECT 94.7000 77.9000 95.1000 80.2000 ;
	    RECT 97.4000 75.9000 97.8000 80.2000 ;
	    RECT 98.2000 75.9000 98.6000 80.2000 ;
	    RECT 99.8000 76.5000 100.2000 80.2000 ;
	    RECT 102.2000 76.5000 102.6000 80.2000 ;
	    RECT 107.0000 76.0000 107.4000 80.2000 ;
	    RECT 109.8000 77.9000 110.2000 80.2000 ;
	    RECT 111.4000 77.9000 111.8000 80.2000 ;
	    RECT 114.2000 75.9000 114.6000 80.2000 ;
	    RECT 116.6000 76.5000 117.0000 80.2000 ;
	    RECT 118.2000 75.9000 118.6000 80.2000 ;
	    RECT 119.8000 76.0000 120.2000 80.2000 ;
	    RECT 122.6000 77.9000 123.0000 80.2000 ;
	    RECT 124.2000 77.9000 124.6000 80.2000 ;
	    RECT 127.0000 75.9000 127.4000 80.2000 ;
	    RECT 129.4000 75.9000 129.8000 80.2000 ;
	    RECT 132.2000 77.9000 132.6000 80.2000 ;
	    RECT 133.8000 77.9000 134.2000 80.2000 ;
	    RECT 136.6000 76.0000 137.0000 80.2000 ;
	    RECT 139.0000 76.5000 139.4000 80.2000 ;
	    RECT 140.6000 75.9000 141.0000 80.2000 ;
	    RECT 141.4000 75.9000 141.8000 80.2000 ;
	    RECT 143.5000 77.9000 143.9000 80.2000 ;
	    RECT 144.6000 75.9000 145.0000 80.2000 ;
	    RECT 146.2000 75.9000 146.6000 80.2000 ;
	    RECT 147.8000 75.9000 148.2000 80.2000 ;
	    RECT 149.4000 75.9000 149.8000 80.2000 ;
	    RECT 151.0000 75.9000 151.4000 80.2000 ;
	    RECT 151.8000 75.9000 152.2000 80.2000 ;
	    RECT 153.4000 75.9000 153.8000 80.2000 ;
	    RECT 155.0000 75.9000 155.4000 80.2000 ;
	    RECT 156.6000 75.9000 157.0000 80.2000 ;
	    RECT 158.2000 75.9000 158.6000 80.2000 ;
	    RECT 160.6000 77.9000 161.0000 80.2000 ;
	    RECT 162.2000 76.1000 162.6000 80.2000 ;
	    RECT 163.8000 77.9000 164.2000 80.2000 ;
	    RECT 165.4000 77.9000 165.8000 80.2000 ;
	    RECT 167.0000 77.9000 167.4000 80.2000 ;
	    RECT 168.6000 76.0000 169.0000 80.2000 ;
	    RECT 171.4000 77.9000 171.8000 80.2000 ;
	    RECT 173.0000 77.9000 173.4000 80.2000 ;
	    RECT 175.8000 75.9000 176.2000 80.2000 ;
	    RECT 177.4000 77.9000 177.8000 80.2000 ;
	    RECT 179.0000 77.9000 179.4000 80.2000 ;
	    RECT 181.4000 76.5000 181.8000 80.2000 ;
	    RECT 183.8000 78.1000 184.2000 80.2000 ;
	    RECT 185.4000 77.9000 185.8000 80.2000 ;
	    RECT 187.8000 75.9000 188.2000 80.2000 ;
	    RECT 188.6000 77.9000 189.0000 80.2000 ;
	    RECT 190.2000 77.9000 190.6000 80.2000 ;
	    RECT 192.3000 75.9000 192.7000 80.2000 ;
	    RECT 194.5000 77.9000 194.9000 80.2000 ;
	    RECT 196.6000 75.9000 197.0000 80.2000 ;
	    RECT 198.5000 75.9000 198.9000 80.2000 ;
	    RECT 202.2000 75.9000 202.6000 80.2000 ;
	    RECT 203.0000 77.9000 203.4000 80.2000 ;
	    RECT 204.6000 77.9000 205.0000 80.2000 ;
	    RECT 207.0000 76.5000 207.4000 80.2000 ;
	    RECT 211.0000 76.0000 211.4000 80.2000 ;
	    RECT 213.8000 77.9000 214.2000 80.2000 ;
	    RECT 215.4000 77.9000 215.8000 80.2000 ;
	    RECT 218.2000 75.9000 218.6000 80.2000 ;
	    RECT 220.6000 77.9000 221.0000 80.2000 ;
	    RECT 221.4000 77.9000 221.8000 80.2000 ;
	    RECT 223.8000 77.9000 224.2000 80.2000 ;
	    RECT 224.6000 75.9000 225.0000 80.2000 ;
	    RECT 226.7000 77.9000 227.1000 80.2000 ;
	    RECT 227.8000 77.9000 228.2000 80.2000 ;
	    RECT 229.4000 78.1000 229.8000 80.2000 ;
	    RECT 231.0000 75.9000 231.4000 80.2000 ;
	    RECT 233.1000 77.9000 233.5000 80.2000 ;
	    RECT 234.5000 77.9000 234.9000 80.2000 ;
	    RECT 236.6000 75.9000 237.0000 80.2000 ;
	    RECT 237.4000 75.9000 237.8000 80.2000 ;
	    RECT 240.6000 77.9000 241.0000 80.2000 ;
	    RECT 241.4000 77.9000 241.8000 80.2000 ;
	    RECT 243.0000 77.9000 243.4000 80.2000 ;
	    RECT 243.8000 75.9000 244.2000 80.2000 ;
	    RECT 247.1000 79.9000 247.5000 80.2000 ;
	    RECT 247.0000 76.6000 247.5000 79.9000 ;
	    RECT 250.1000 76.6000 250.6000 80.2000 ;
	    RECT 252.6000 78.1000 253.0000 80.2000 ;
	    RECT 254.2000 77.9000 254.6000 80.2000 ;
	    RECT 255.0000 77.9000 255.4000 80.2000 ;
	    RECT 256.6000 77.9000 257.0000 80.2000 ;
	    RECT 257.7000 77.9000 258.1000 80.2000 ;
	    RECT 259.8000 75.9000 260.2000 80.2000 ;
	    RECT 260.9000 77.9000 261.3000 80.2000 ;
	    RECT 263.0000 75.9000 263.4000 80.2000 ;
	    RECT 263.8000 75.9000 264.2000 80.2000 ;
	    RECT 266.2000 77.9000 266.6000 80.2000 ;
	    RECT 267.8000 77.9000 268.2000 80.2000 ;
	    RECT 269.4000 77.9000 269.8000 80.2000 ;
	    RECT 0.6000 60.8000 1.0000 63.1000 ;
	    RECT 2.2000 60.8000 2.6000 63.1000 ;
	    RECT 3.8000 60.8000 4.2000 63.1000 ;
	    RECT 6.2000 60.8000 6.6000 65.1000 ;
	    RECT 8.6000 60.8000 9.0000 64.5000 ;
	    RECT 10.5000 60.8000 10.9000 63.1000 ;
	    RECT 12.6000 60.8000 13.0000 65.1000 ;
	    RECT 15.0000 60.8000 15.4000 65.1000 ;
	    RECT 16.6000 60.8000 17.0000 64.5000 ;
	    RECT 19.0000 60.8000 19.4000 63.1000 ;
	    RECT 20.6000 60.8000 21.0000 63.1000 ;
	    RECT 22.2000 60.8000 22.6000 64.5000 ;
	    RECT 24.6000 60.8000 25.0000 65.1000 ;
	    RECT 28.6000 60.8000 29.0000 64.5000 ;
	    RECT 30.2000 60.8000 30.6000 63.1000 ;
	    RECT 31.8000 60.8000 32.2000 63.1000 ;
	    RECT 33.4000 60.8000 33.8000 63.1000 ;
	    RECT 34.2000 60.8000 34.6000 63.1000 ;
	    RECT 35.8000 60.8000 36.2000 63.1000 ;
	    RECT 36.6000 60.8000 37.0000 65.1000 ;
	    RECT 39.8000 60.8000 40.2000 65.1000 ;
	    RECT 41.4000 60.8000 41.8000 62.9000 ;
	    RECT 43.0000 60.8000 43.4000 63.1000 ;
	    RECT 43.8000 60.8000 44.2000 63.1000 ;
	    RECT 45.4000 60.8000 45.8000 63.1000 ;
	    RECT 47.0000 60.8000 47.4000 63.1000 ;
	    RECT 47.8000 60.8000 48.2000 65.1000 ;
	    RECT 51.0000 60.8000 51.4000 65.0000 ;
	    RECT 53.8000 60.8000 54.2000 63.1000 ;
	    RECT 55.4000 60.8000 55.8000 63.1000 ;
	    RECT 58.2000 60.8000 58.6000 65.1000 ;
	    RECT 61.4000 60.8000 61.8000 65.1000 ;
	    RECT 63.8000 60.8000 64.2000 63.1000 ;
	    RECT 65.4000 60.8000 65.8000 62.9000 ;
	    RECT 67.0000 60.8000 67.4000 65.1000 ;
	    RECT 69.1000 60.8000 69.5000 63.1000 ;
	    RECT 71.8000 60.8000 72.2000 65.1000 ;
	    RECT 73.4000 60.8000 73.8000 65.0000 ;
	    RECT 76.2000 60.8000 76.6000 63.1000 ;
	    RECT 77.8000 60.8000 78.2000 63.1000 ;
	    RECT 80.6000 60.8000 81.0000 65.1000 ;
	    RECT 82.5000 60.8000 82.9000 63.1000 ;
	    RECT 84.6000 60.8000 85.0000 65.1000 ;
	    RECT 87.0000 60.8000 87.4000 64.5000 ;
	    RECT 88.6000 60.8000 89.0000 63.1000 ;
	    RECT 90.2000 60.8000 90.6000 62.9000 ;
	    RECT 91.8000 60.8000 92.2000 65.1000 ;
	    RECT 93.4000 60.8000 93.8000 64.5000 ;
	    RECT 95.0000 60.8000 95.4000 65.1000 ;
	    RECT 96.6000 60.8000 97.0000 64.5000 ;
	    RECT 98.2000 60.8000 98.6000 65.1000 ;
	    RECT 99.8000 60.8000 100.2000 64.5000 ;
	    RECT 101.4000 60.8000 101.8000 65.1000 ;
	    RECT 103.0000 60.8000 103.4000 64.5000 ;
	    RECT 104.6000 60.8000 105.0000 65.1000 ;
	    RECT 106.2000 60.8000 106.6000 64.5000 ;
	    RECT 110.2000 60.8000 110.6000 64.5000 ;
	    RECT 111.8000 60.8000 112.2000 65.1000 ;
	    RECT 113.4000 60.8000 113.8000 64.5000 ;
	    RECT 115.0000 60.8000 115.4000 65.1000 ;
	    RECT 115.8000 60.8000 116.2000 63.1000 ;
	    RECT 117.4000 60.8000 117.8000 62.9000 ;
	    RECT 120.6000 60.8000 121.0000 64.5000 ;
	    RECT 122.5000 60.8000 122.9000 63.1000 ;
	    RECT 124.6000 60.8000 125.0000 65.1000 ;
	    RECT 125.7000 60.8000 126.1000 63.1000 ;
	    RECT 127.8000 60.8000 128.2000 65.1000 ;
	    RECT 129.4000 60.8000 129.8000 64.5000 ;
	    RECT 131.0000 60.8000 131.4000 65.1000 ;
	    RECT 132.6000 60.8000 133.0000 64.5000 ;
	    RECT 134.2000 60.8000 134.6000 65.1000 ;
	    RECT 135.0000 60.8000 135.4000 65.1000 ;
	    RECT 136.6000 60.8000 137.0000 65.1000 ;
	    RECT 138.2000 60.8000 138.6000 65.1000 ;
	    RECT 139.3000 60.8000 139.7000 63.1000 ;
	    RECT 141.4000 60.8000 141.8000 65.1000 ;
	    RECT 143.0000 60.8000 143.4000 64.5000 ;
	    RECT 145.4000 60.8000 145.8000 65.1000 ;
	    RECT 147.5000 60.8000 147.9000 63.1000 ;
	    RECT 149.4000 60.8000 149.8000 64.5000 ;
	    RECT 152.6000 60.8000 153.0000 65.1000 ;
	    RECT 155.4000 60.8000 155.8000 63.1000 ;
	    RECT 157.0000 60.8000 157.4000 63.1000 ;
	    RECT 159.8000 60.8000 160.2000 65.0000 ;
	    RECT 163.0000 60.8000 163.4000 63.1000 ;
	    RECT 164.6000 60.8000 165.0000 63.1000 ;
	    RECT 166.2000 60.8000 166.6000 63.1000 ;
	    RECT 167.0000 60.8000 167.4000 65.1000 ;
	    RECT 168.6000 60.8000 169.0000 64.5000 ;
	    RECT 171.0000 60.8000 171.4000 64.5000 ;
	    RECT 172.6000 60.8000 173.0000 65.1000 ;
	    RECT 174.2000 60.8000 174.6000 63.1000 ;
	    RECT 175.0000 60.8000 175.4000 63.1000 ;
	    RECT 176.6000 60.8000 177.0000 63.1000 ;
	    RECT 178.2000 60.8000 178.6000 63.1000 ;
	    RECT 179.8000 60.8000 180.2000 64.9000 ;
	    RECT 182.4000 60.8000 182.8000 65.1000 ;
	    RECT 183.8000 60.8000 184.2000 65.1000 ;
	    RECT 187.5000 60.8000 187.9000 65.1000 ;
	    RECT 190.0000 60.8000 190.4000 65.1000 ;
	    RECT 192.6000 60.8000 193.0000 64.9000 ;
	    RECT 195.0000 60.8000 195.5000 64.4000 ;
	    RECT 198.1000 61.1000 198.6000 64.4000 ;
	    RECT 198.1000 60.8000 198.5000 61.1000 ;
	    RECT 200.6000 60.8000 201.0000 64.5000 ;
	    RECT 202.2000 60.8000 202.6000 63.1000 ;
	    RECT 203.8000 60.8000 204.2000 63.1000 ;
	    RECT 205.4000 60.8000 205.8000 63.1000 ;
	    RECT 206.2000 60.8000 206.6000 65.1000 ;
	    RECT 207.8000 60.8000 208.2000 65.1000 ;
	    RECT 208.6000 60.8000 209.0000 65.1000 ;
	    RECT 214.2000 60.8000 214.6000 65.1000 ;
	    RECT 215.8000 60.8000 216.2000 62.9000 ;
	    RECT 217.4000 60.8000 217.8000 63.1000 ;
	    RECT 218.2000 60.8000 218.6000 63.1000 ;
	    RECT 219.8000 60.8000 220.2000 63.1000 ;
	    RECT 222.2000 60.8000 222.6000 64.5000 ;
	    RECT 223.8000 60.8000 224.2000 65.1000 ;
	    RECT 225.9000 60.8000 226.3000 63.1000 ;
	    RECT 227.0000 60.8000 227.4000 63.1000 ;
	    RECT 228.6000 60.8000 229.0000 63.1000 ;
	    RECT 229.7000 60.8000 230.1000 63.1000 ;
	    RECT 231.8000 60.8000 232.2000 65.1000 ;
	    RECT 232.6000 60.8000 233.0000 63.1000 ;
	    RECT 234.5000 60.8000 234.9000 63.1000 ;
	    RECT 236.6000 60.8000 237.0000 65.1000 ;
	    RECT 237.4000 60.8000 237.8000 65.1000 ;
	    RECT 239.5000 60.8000 239.9000 63.1000 ;
	    RECT 241.4000 60.8000 241.8000 64.5000 ;
	    RECT 243.8000 60.8000 244.2000 63.1000 ;
	    RECT 245.4000 60.8000 245.8000 63.1000 ;
	    RECT 247.0000 60.8000 247.4000 63.1000 ;
	    RECT 248.6000 60.8000 249.0000 62.9000 ;
	    RECT 251.8000 60.8000 252.2000 65.1000 ;
	    RECT 252.6000 60.8000 253.0000 65.1000 ;
	    RECT 254.7000 60.8000 255.1000 63.1000 ;
	    RECT 256.6000 60.8000 257.0000 63.1000 ;
	    RECT 258.2000 61.1000 258.7000 64.4000 ;
	    RECT 258.3000 60.8000 258.7000 61.1000 ;
	    RECT 261.3000 60.8000 261.8000 64.4000 ;
	    RECT 263.0000 60.8000 263.4000 65.1000 ;
	    RECT 264.6000 60.8000 265.0000 64.5000 ;
	    RECT 267.0000 60.8000 267.4000 64.5000 ;
	    RECT 268.6000 60.8000 269.0000 65.1000 ;
	    RECT 0.2000 60.2000 271.0000 60.8000 ;
	    RECT 1.5000 59.9000 1.9000 60.2000 ;
	    RECT 1.4000 56.6000 1.9000 59.9000 ;
	    RECT 4.5000 56.6000 5.0000 60.2000 ;
	    RECT 6.2000 57.9000 6.6000 60.2000 ;
	    RECT 9.4000 55.9000 9.8000 60.2000 ;
	    RECT 10.2000 57.9000 10.6000 60.2000 ;
	    RECT 12.1000 57.9000 12.5000 60.2000 ;
	    RECT 14.2000 55.9000 14.6000 60.2000 ;
	    RECT 15.0000 57.9000 15.4000 60.2000 ;
	    RECT 16.6000 55.9000 17.0000 60.2000 ;
	    RECT 20.6000 56.5000 21.0000 60.2000 ;
	    RECT 22.2000 57.9000 22.6000 60.2000 ;
	    RECT 23.8000 57.9000 24.2000 60.2000 ;
	    RECT 25.5000 59.9000 25.9000 60.2000 ;
	    RECT 25.4000 56.6000 25.9000 59.9000 ;
	    RECT 28.5000 56.6000 29.0000 60.2000 ;
	    RECT 30.5000 57.9000 30.9000 60.2000 ;
	    RECT 32.6000 55.9000 33.0000 60.2000 ;
	    RECT 33.4000 57.9000 33.8000 60.2000 ;
	    RECT 35.0000 57.9000 35.4000 60.2000 ;
	    RECT 36.6000 57.9000 37.0000 60.2000 ;
	    RECT 38.2000 56.5000 38.6000 60.2000 ;
	    RECT 42.2000 55.9000 42.6000 60.2000 ;
	    RECT 43.8000 55.9000 44.2000 60.2000 ;
	    RECT 46.6000 57.9000 47.0000 60.2000 ;
	    RECT 48.2000 57.9000 48.6000 60.2000 ;
	    RECT 51.0000 56.0000 51.4000 60.2000 ;
	    RECT 53.7000 55.9000 54.1000 60.2000 ;
	    RECT 58.2000 55.9000 58.6000 60.2000 ;
	    RECT 61.0000 57.9000 61.4000 60.2000 ;
	    RECT 62.6000 57.9000 63.0000 60.2000 ;
	    RECT 65.4000 56.0000 65.8000 60.2000 ;
	    RECT 68.6000 56.5000 69.0000 60.2000 ;
	    RECT 70.5000 57.9000 70.9000 60.2000 ;
	    RECT 72.6000 55.9000 73.0000 60.2000 ;
	    RECT 73.7000 57.9000 74.1000 60.2000 ;
	    RECT 75.8000 55.9000 76.2000 60.2000 ;
	    RECT 77.4000 56.5000 77.8000 60.2000 ;
	    RECT 80.6000 58.1000 81.0000 60.2000 ;
	    RECT 82.2000 57.9000 82.6000 60.2000 ;
	    RECT 83.8000 55.9000 84.2000 60.2000 ;
	    RECT 86.6000 57.9000 87.0000 60.2000 ;
	    RECT 88.2000 57.9000 88.6000 60.2000 ;
	    RECT 91.0000 56.0000 91.4000 60.2000 ;
	    RECT 92.6000 55.9000 93.0000 60.2000 ;
	    RECT 94.2000 56.5000 94.6000 60.2000 ;
	    RECT 95.8000 55.9000 96.2000 60.2000 ;
	    RECT 97.4000 56.5000 97.8000 60.2000 ;
	    RECT 99.0000 57.9000 99.4000 60.2000 ;
	    RECT 100.6000 56.1000 101.0000 60.2000 ;
	    RECT 102.2000 57.9000 102.6000 60.2000 ;
	    RECT 103.8000 57.9000 104.2000 60.2000 ;
	    RECT 104.6000 55.9000 105.0000 60.2000 ;
	    RECT 106.2000 56.5000 106.6000 60.2000 ;
	    RECT 110.2000 55.9000 110.6000 60.2000 ;
	    RECT 113.0000 57.9000 113.4000 60.2000 ;
	    RECT 114.6000 57.9000 115.0000 60.2000 ;
	    RECT 117.4000 56.0000 117.8000 60.2000 ;
	    RECT 120.6000 56.5000 121.0000 60.2000 ;
	    RECT 122.2000 57.9000 122.6000 60.2000 ;
	    RECT 123.8000 58.1000 124.2000 60.2000 ;
	    RECT 125.4000 55.9000 125.8000 60.2000 ;
	    RECT 127.0000 57.9000 127.4000 60.2000 ;
	    RECT 128.6000 55.9000 129.0000 60.2000 ;
	    RECT 130.7000 57.9000 131.1000 60.2000 ;
	    RECT 132.6000 56.5000 133.0000 60.2000 ;
	    RECT 135.8000 56.0000 136.2000 60.2000 ;
	    RECT 138.6000 57.9000 139.0000 60.2000 ;
	    RECT 140.2000 57.9000 140.6000 60.2000 ;
	    RECT 143.0000 55.9000 143.4000 60.2000 ;
	    RECT 145.4000 58.1000 145.8000 60.2000 ;
	    RECT 147.0000 57.9000 147.4000 60.2000 ;
	    RECT 147.8000 57.9000 148.2000 60.2000 ;
	    RECT 149.4000 58.1000 149.8000 60.2000 ;
	    RECT 151.8000 56.5000 152.2000 60.2000 ;
	    RECT 154.2000 56.5000 154.6000 60.2000 ;
	    RECT 156.6000 55.9000 157.0000 60.2000 ;
	    RECT 158.7000 57.9000 159.1000 60.2000 ;
	    RECT 162.2000 56.0000 162.6000 60.2000 ;
	    RECT 165.0000 57.9000 165.4000 60.2000 ;
	    RECT 166.6000 57.9000 167.0000 60.2000 ;
	    RECT 169.4000 55.9000 169.8000 60.2000 ;
	    RECT 171.0000 57.9000 171.4000 60.2000 ;
	    RECT 172.6000 57.9000 173.0000 60.2000 ;
	    RECT 175.0000 56.5000 175.4000 60.2000 ;
	    RECT 176.6000 57.9000 177.0000 60.2000 ;
	    RECT 178.2000 57.9000 178.6000 60.2000 ;
	    RECT 179.8000 57.9000 180.2000 60.2000 ;
	    RECT 182.2000 56.5000 182.6000 60.2000 ;
	    RECT 184.6000 56.0000 185.0000 60.2000 ;
	    RECT 187.4000 57.9000 187.8000 60.2000 ;
	    RECT 189.0000 57.9000 189.4000 60.2000 ;
	    RECT 191.8000 55.9000 192.2000 60.2000 ;
	    RECT 194.2000 57.9000 194.6000 60.2000 ;
	    RECT 195.8000 55.9000 196.2000 60.2000 ;
	    RECT 198.6000 57.9000 199.0000 60.2000 ;
	    RECT 200.2000 57.9000 200.6000 60.2000 ;
	    RECT 203.0000 56.0000 203.4000 60.2000 ;
	    RECT 206.2000 56.5000 206.6000 60.2000 ;
	    RECT 210.2000 56.0000 210.6000 60.2000 ;
	    RECT 213.0000 57.9000 213.4000 60.2000 ;
	    RECT 214.6000 57.9000 215.0000 60.2000 ;
	    RECT 217.4000 55.9000 217.8000 60.2000 ;
	    RECT 219.8000 56.0000 220.2000 60.2000 ;
	    RECT 222.6000 57.9000 223.0000 60.2000 ;
	    RECT 224.2000 57.9000 224.6000 60.2000 ;
	    RECT 227.0000 55.9000 227.4000 60.2000 ;
	    RECT 230.2000 55.9000 230.6000 60.2000 ;
	    RECT 231.0000 57.9000 231.4000 60.2000 ;
	    RECT 232.6000 56.1000 233.0000 60.2000 ;
	    RECT 235.0000 55.9000 235.4000 60.2000 ;
	    RECT 237.8000 57.9000 238.2000 60.2000 ;
	    RECT 239.4000 57.9000 239.8000 60.2000 ;
	    RECT 242.2000 56.0000 242.6000 60.2000 ;
	    RECT 243.8000 57.9000 244.2000 60.2000 ;
	    RECT 245.4000 57.9000 245.8000 60.2000 ;
	    RECT 247.0000 56.1000 247.4000 60.2000 ;
	    RECT 249.4000 56.9000 249.8000 60.2000 ;
	    RECT 256.6000 55.9000 257.0000 60.2000 ;
	    RECT 259.0000 56.5000 259.4000 60.2000 ;
	    RECT 260.6000 55.9000 261.0000 60.2000 ;
	    RECT 262.7000 57.9000 263.1000 60.2000 ;
	    RECT 263.8000 57.9000 264.2000 60.2000 ;
	    RECT 265.4000 57.9000 265.8000 60.2000 ;
	    RECT 267.0000 57.9000 267.4000 60.2000 ;
	    RECT 267.8000 55.9000 268.2000 60.2000 ;
	    RECT 1.4000 40.8000 1.9000 44.4000 ;
	    RECT 4.5000 41.1000 5.0000 44.4000 ;
	    RECT 4.5000 40.8000 4.9000 41.1000 ;
	    RECT 6.2000 40.8000 6.6000 43.1000 ;
	    RECT 7.8000 40.8000 8.2000 43.1000 ;
	    RECT 10.2000 40.8000 10.6000 44.5000 ;
	    RECT 12.6000 40.8000 13.0000 43.1000 ;
	    RECT 15.0000 40.8000 15.4000 45.1000 ;
	    RECT 15.8000 40.8000 16.2000 43.1000 ;
	    RECT 17.4000 40.8000 17.8000 43.1000 ;
	    RECT 19.0000 41.1000 19.5000 44.4000 ;
	    RECT 19.1000 40.8000 19.5000 41.1000 ;
	    RECT 22.1000 40.8000 22.6000 44.4000 ;
	    RECT 23.8000 40.8000 24.2000 43.1000 ;
	    RECT 25.4000 40.8000 25.8000 43.1000 ;
	    RECT 27.0000 40.8000 27.4000 43.1000 ;
	    RECT 27.8000 40.8000 28.2000 45.1000 ;
	    RECT 31.0000 40.8000 31.4000 43.1000 ;
	    RECT 32.6000 41.1000 33.1000 44.4000 ;
	    RECT 32.7000 40.8000 33.1000 41.1000 ;
	    RECT 35.7000 40.8000 36.2000 44.4000 ;
	    RECT 38.2000 40.8000 38.6000 43.1000 ;
	    RECT 39.0000 40.8000 39.4000 43.1000 ;
	    RECT 40.6000 40.8000 41.0000 43.1000 ;
	    RECT 41.4000 40.8000 41.8000 43.1000 ;
	    RECT 43.8000 40.8000 44.2000 45.1000 ;
	    RECT 46.6000 40.8000 47.0000 43.1000 ;
	    RECT 48.2000 40.8000 48.6000 43.1000 ;
	    RECT 51.0000 40.8000 51.4000 45.0000 ;
	    RECT 53.7000 40.8000 54.1000 45.1000 ;
	    RECT 56.6000 40.8000 57.0000 44.5000 ;
	    RECT 58.2000 40.8000 58.6000 45.1000 ;
	    RECT 60.6000 40.8000 61.0000 43.1000 ;
	    RECT 67.0000 40.8000 67.4000 44.1000 ;
	    RECT 68.6000 40.8000 69.0000 45.1000 ;
	    RECT 71.8000 40.8000 72.2000 43.1000 ;
	    RECT 72.6000 40.8000 73.0000 43.1000 ;
	    RECT 74.2000 40.8000 74.6000 45.1000 ;
	    RECT 76.9000 40.8000 77.3000 43.1000 ;
	    RECT 79.0000 40.8000 79.4000 45.1000 ;
	    RECT 80.6000 40.8000 81.0000 45.0000 ;
	    RECT 83.4000 40.8000 83.8000 43.1000 ;
	    RECT 85.0000 40.8000 85.4000 43.1000 ;
	    RECT 87.8000 40.8000 88.2000 45.1000 ;
	    RECT 89.7000 40.8000 90.1000 43.1000 ;
	    RECT 91.8000 40.8000 92.2000 45.1000 ;
	    RECT 93.4000 40.8000 93.8000 44.5000 ;
	    RECT 96.6000 40.8000 97.0000 44.5000 ;
	    RECT 99.3000 40.8000 99.7000 43.1000 ;
	    RECT 101.4000 40.8000 101.8000 45.1000 ;
	    RECT 102.2000 40.8000 102.6000 45.1000 ;
	    RECT 104.3000 40.8000 104.7000 43.1000 ;
	    RECT 106.2000 40.8000 106.6000 44.5000 ;
	    RECT 111.0000 40.8000 111.4000 42.9000 ;
	    RECT 112.6000 40.8000 113.0000 43.1000 ;
	    RECT 114.2000 40.8000 114.6000 45.1000 ;
	    RECT 117.0000 40.8000 117.4000 43.1000 ;
	    RECT 118.6000 40.8000 119.0000 43.1000 ;
	    RECT 121.4000 40.8000 121.8000 45.0000 ;
	    RECT 123.0000 40.8000 123.4000 43.1000 ;
	    RECT 124.6000 40.8000 125.0000 43.1000 ;
	    RECT 127.0000 40.8000 127.4000 45.1000 ;
	    RECT 129.4000 40.8000 129.8000 44.5000 ;
	    RECT 131.0000 40.8000 131.4000 43.1000 ;
	    RECT 132.6000 40.8000 133.0000 44.9000 ;
	    RECT 134.2000 40.8000 134.6000 45.1000 ;
	    RECT 135.8000 40.8000 136.2000 45.1000 ;
	    RECT 137.4000 40.8000 137.8000 45.1000 ;
	    RECT 139.0000 40.8000 139.4000 45.1000 ;
	    RECT 140.6000 40.8000 141.0000 45.1000 ;
	    RECT 142.2000 40.8000 142.6000 45.0000 ;
	    RECT 145.0000 40.8000 145.4000 43.1000 ;
	    RECT 146.6000 40.8000 147.0000 43.1000 ;
	    RECT 149.4000 40.8000 149.8000 45.1000 ;
	    RECT 151.8000 40.8000 152.2000 45.0000 ;
	    RECT 154.6000 40.8000 155.0000 43.1000 ;
	    RECT 156.2000 40.8000 156.6000 43.1000 ;
	    RECT 159.0000 40.8000 159.4000 45.1000 ;
	    RECT 162.2000 40.8000 162.6000 45.1000 ;
	    RECT 165.4000 40.8000 165.8000 43.1000 ;
	    RECT 167.0000 40.8000 167.4000 45.1000 ;
	    RECT 169.8000 40.8000 170.2000 43.1000 ;
	    RECT 171.4000 40.8000 171.8000 43.1000 ;
	    RECT 174.2000 40.8000 174.6000 45.0000 ;
	    RECT 175.8000 40.8000 176.2000 43.1000 ;
	    RECT 178.2000 40.8000 178.6000 45.1000 ;
	    RECT 181.0000 40.8000 181.4000 43.1000 ;
	    RECT 182.6000 40.8000 183.0000 43.1000 ;
	    RECT 185.4000 40.8000 185.8000 45.0000 ;
	    RECT 187.0000 40.8000 187.4000 43.1000 ;
	    RECT 188.6000 40.8000 189.0000 44.9000 ;
	    RECT 191.0000 40.8000 191.4000 45.0000 ;
	    RECT 193.8000 40.8000 194.2000 43.1000 ;
	    RECT 195.4000 40.8000 195.8000 43.1000 ;
	    RECT 198.2000 40.8000 198.6000 45.1000 ;
	    RECT 200.6000 40.8000 201.0000 44.9000 ;
	    RECT 202.2000 40.8000 202.6000 43.1000 ;
	    RECT 203.0000 40.8000 203.4000 45.1000 ;
	    RECT 205.1000 40.8000 205.5000 43.1000 ;
	    RECT 207.0000 40.8000 207.4000 44.5000 ;
	    RECT 211.0000 40.8000 211.4000 45.0000 ;
	    RECT 213.8000 40.8000 214.2000 43.1000 ;
	    RECT 215.4000 40.8000 215.8000 43.1000 ;
	    RECT 218.2000 40.8000 218.6000 45.1000 ;
	    RECT 220.6000 40.8000 221.0000 45.0000 ;
	    RECT 223.4000 40.8000 223.8000 43.1000 ;
	    RECT 225.0000 40.8000 225.4000 43.1000 ;
	    RECT 227.8000 40.8000 228.2000 45.1000 ;
	    RECT 230.2000 40.8000 230.6000 45.1000 ;
	    RECT 233.0000 40.8000 233.4000 43.1000 ;
	    RECT 234.6000 40.8000 235.0000 43.1000 ;
	    RECT 237.4000 40.8000 237.8000 45.0000 ;
	    RECT 239.8000 40.8000 240.2000 45.1000 ;
	    RECT 242.6000 40.8000 243.0000 43.1000 ;
	    RECT 244.2000 40.8000 244.6000 43.1000 ;
	    RECT 247.0000 40.8000 247.4000 45.0000 ;
	    RECT 248.6000 40.8000 249.0000 45.1000 ;
	    RECT 250.7000 40.8000 251.1000 43.1000 ;
	    RECT 252.1000 40.8000 252.5000 43.1000 ;
	    RECT 254.2000 40.8000 254.6000 45.1000 ;
	    RECT 255.8000 40.8000 256.2000 44.5000 ;
	    RECT 259.0000 40.8000 259.4000 45.1000 ;
	    RECT 261.8000 40.8000 262.2000 43.1000 ;
	    RECT 263.4000 40.8000 263.8000 43.1000 ;
	    RECT 266.2000 40.8000 266.6000 45.0000 ;
	    RECT 267.8000 40.8000 268.2000 43.1000 ;
	    RECT 269.4000 40.8000 269.8000 43.1000 ;
	    RECT 0.2000 40.2000 271.0000 40.8000 ;
	    RECT 1.5000 39.9000 1.9000 40.2000 ;
	    RECT 1.4000 36.6000 1.9000 39.9000 ;
	    RECT 4.5000 36.6000 5.0000 40.2000 ;
	    RECT 7.1000 39.9000 7.5000 40.2000 ;
	    RECT 7.0000 36.6000 7.5000 39.9000 ;
	    RECT 10.1000 36.6000 10.6000 40.2000 ;
	    RECT 11.8000 37.9000 12.2000 40.2000 ;
	    RECT 13.4000 37.9000 13.8000 40.2000 ;
	    RECT 15.0000 37.9000 15.4000 40.2000 ;
	    RECT 17.4000 35.9000 17.8000 40.2000 ;
	    RECT 18.5000 37.9000 18.9000 40.2000 ;
	    RECT 20.6000 35.9000 21.0000 40.2000 ;
	    RECT 21.4000 35.9000 21.8000 40.2000 ;
	    RECT 23.8000 37.9000 24.2000 40.2000 ;
	    RECT 25.4000 35.9000 25.8000 40.2000 ;
	    RECT 27.5000 37.9000 27.9000 40.2000 ;
	    RECT 28.6000 35.9000 29.0000 40.2000 ;
	    RECT 32.6000 35.9000 33.0000 40.2000 ;
	    RECT 33.4000 37.9000 33.8000 40.2000 ;
	    RECT 35.0000 37.9000 35.4000 40.2000 ;
	    RECT 36.6000 36.6000 37.1000 40.2000 ;
	    RECT 39.7000 39.9000 40.1000 40.2000 ;
	    RECT 39.7000 36.6000 40.2000 39.9000 ;
	    RECT 41.4000 37.9000 41.8000 40.2000 ;
	    RECT 43.0000 35.9000 43.4000 40.2000 ;
	    RECT 45.4000 35.9000 45.8000 40.2000 ;
	    RECT 47.0000 35.9000 47.4000 40.2000 ;
	    RECT 48.6000 36.5000 49.0000 40.2000 ;
	    RECT 51.0000 35.9000 51.4000 40.2000 ;
	    RECT 53.8000 37.9000 54.2000 40.2000 ;
	    RECT 55.4000 37.9000 55.8000 40.2000 ;
	    RECT 58.2000 36.0000 58.6000 40.2000 ;
	    RECT 62.2000 38.1000 62.6000 40.2000 ;
	    RECT 63.8000 37.9000 64.2000 40.2000 ;
	    RECT 64.6000 37.9000 65.0000 40.2000 ;
	    RECT 66.2000 37.9000 66.6000 40.2000 ;
	    RECT 67.0000 37.9000 67.4000 40.2000 ;
	    RECT 68.6000 35.9000 69.0000 40.2000 ;
	    RECT 70.7000 37.9000 71.1000 40.2000 ;
	    RECT 72.6000 35.9000 73.0000 40.2000 ;
	    RECT 75.4000 37.9000 75.8000 40.2000 ;
	    RECT 77.0000 37.9000 77.4000 40.2000 ;
	    RECT 79.8000 36.0000 80.2000 40.2000 ;
	    RECT 81.4000 37.9000 81.8000 40.2000 ;
	    RECT 83.0000 38.1000 83.4000 40.2000 ;
	    RECT 84.6000 37.9000 85.0000 40.2000 ;
	    RECT 86.2000 38.1000 86.6000 40.2000 ;
	    RECT 92.6000 36.9000 93.0000 40.2000 ;
	    RECT 95.0000 37.9000 95.4000 40.2000 ;
	    RECT 96.1000 37.9000 96.5000 40.2000 ;
	    RECT 98.2000 35.9000 98.6000 40.2000 ;
	    RECT 99.0000 35.9000 99.4000 40.2000 ;
	    RECT 101.1000 37.9000 101.5000 40.2000 ;
	    RECT 102.2000 35.9000 102.6000 40.2000 ;
	    RECT 104.3000 37.9000 104.7000 40.2000 ;
	    RECT 107.8000 36.0000 108.2000 40.2000 ;
	    RECT 110.6000 37.9000 111.0000 40.2000 ;
	    RECT 112.2000 37.9000 112.6000 40.2000 ;
	    RECT 115.0000 35.9000 115.4000 40.2000 ;
	    RECT 116.6000 35.9000 117.0000 40.2000 ;
	    RECT 118.7000 37.9000 119.1000 40.2000 ;
	    RECT 122.2000 36.5000 122.6000 40.2000 ;
	    RECT 123.8000 37.9000 124.2000 40.2000 ;
	    RECT 125.4000 38.1000 125.8000 40.2000 ;
	    RECT 127.8000 36.0000 128.2000 40.2000 ;
	    RECT 130.6000 37.9000 131.0000 40.2000 ;
	    RECT 132.2000 37.9000 132.6000 40.2000 ;
	    RECT 135.0000 35.9000 135.4000 40.2000 ;
	    RECT 136.6000 37.9000 137.0000 40.2000 ;
	    RECT 138.2000 36.1000 138.6000 40.2000 ;
	    RECT 140.9000 35.9000 141.3000 40.2000 ;
	    RECT 143.8000 36.0000 144.2000 40.2000 ;
	    RECT 146.6000 37.9000 147.0000 40.2000 ;
	    RECT 148.2000 37.9000 148.6000 40.2000 ;
	    RECT 151.0000 35.9000 151.4000 40.2000 ;
	    RECT 152.6000 37.9000 153.0000 40.2000 ;
	    RECT 154.2000 37.9000 154.6000 40.2000 ;
	    RECT 155.0000 37.9000 155.4000 40.2000 ;
	    RECT 156.6000 37.9000 157.0000 40.2000 ;
	    RECT 158.2000 37.9000 158.6000 40.2000 ;
	    RECT 161.4000 35.9000 161.8000 40.2000 ;
	    RECT 164.2000 37.9000 164.6000 40.2000 ;
	    RECT 165.8000 37.9000 166.2000 40.2000 ;
	    RECT 168.6000 36.0000 169.0000 40.2000 ;
	    RECT 170.2000 37.9000 170.6000 40.2000 ;
	    RECT 171.8000 35.9000 172.2000 40.2000 ;
	    RECT 175.0000 37.9000 175.4000 40.2000 ;
	    RECT 176.6000 36.5000 177.0000 40.2000 ;
	    RECT 178.2000 35.9000 178.6000 40.2000 ;
	    RECT 179.8000 36.0000 180.2000 40.2000 ;
	    RECT 182.6000 37.9000 183.0000 40.2000 ;
	    RECT 184.2000 37.9000 184.6000 40.2000 ;
	    RECT 187.0000 35.9000 187.4000 40.2000 ;
	    RECT 189.4000 36.5000 189.8000 40.2000 ;
	    RECT 191.8000 35.9000 192.2000 40.2000 ;
	    RECT 193.9000 37.9000 194.3000 40.2000 ;
	    RECT 195.8000 36.0000 196.2000 40.2000 ;
	    RECT 198.6000 37.9000 199.0000 40.2000 ;
	    RECT 200.2000 37.9000 200.6000 40.2000 ;
	    RECT 203.0000 35.9000 203.4000 40.2000 ;
	    RECT 204.6000 37.9000 205.0000 40.2000 ;
	    RECT 206.2000 36.1000 206.6000 40.2000 ;
	    RECT 210.2000 36.0000 210.6000 40.2000 ;
	    RECT 213.0000 37.9000 213.4000 40.2000 ;
	    RECT 214.6000 37.9000 215.0000 40.2000 ;
	    RECT 217.4000 35.9000 217.8000 40.2000 ;
	    RECT 219.0000 37.9000 219.4000 40.2000 ;
	    RECT 220.6000 36.1000 221.0000 40.2000 ;
	    RECT 223.0000 36.0000 223.4000 40.2000 ;
	    RECT 225.8000 37.9000 226.2000 40.2000 ;
	    RECT 227.4000 37.9000 227.8000 40.2000 ;
	    RECT 230.2000 35.9000 230.6000 40.2000 ;
	    RECT 232.1000 37.9000 232.5000 40.2000 ;
	    RECT 234.2000 35.9000 234.6000 40.2000 ;
	    RECT 235.8000 36.5000 236.2000 40.2000 ;
	    RECT 238.5000 37.9000 238.9000 40.2000 ;
	    RECT 240.6000 35.9000 241.0000 40.2000 ;
	    RECT 241.4000 35.9000 241.8000 40.2000 ;
	    RECT 245.4000 36.5000 245.8000 40.2000 ;
	    RECT 247.0000 35.9000 247.4000 40.2000 ;
	    RECT 248.6000 35.9000 249.0000 40.2000 ;
	    RECT 249.4000 35.9000 249.8000 40.2000 ;
	    RECT 251.8000 37.9000 252.2000 40.2000 ;
	    RECT 253.4000 35.9000 253.8000 40.2000 ;
	    RECT 255.5000 37.9000 255.9000 40.2000 ;
	    RECT 257.4000 36.1000 257.8000 40.2000 ;
	    RECT 259.0000 37.9000 259.4000 40.2000 ;
	    RECT 259.8000 35.9000 260.2000 40.2000 ;
	    RECT 261.9000 37.9000 262.3000 40.2000 ;
	    RECT 263.8000 37.9000 264.2000 40.2000 ;
	    RECT 266.2000 36.5000 266.6000 40.2000 ;
	    RECT 267.8000 37.9000 268.2000 40.2000 ;
	    RECT 0.6000 20.8000 1.0000 23.1000 ;
	    RECT 3.8000 20.8000 4.2000 25.1000 ;
	    RECT 4.6000 20.8000 5.0000 23.1000 ;
	    RECT 6.2000 20.8000 6.6000 23.1000 ;
	    RECT 7.8000 20.8000 8.2000 24.5000 ;
	    RECT 11.8000 20.8000 12.2000 25.1000 ;
	    RECT 13.4000 20.8000 13.8000 23.1000 ;
	    RECT 14.2000 20.8000 14.6000 23.1000 ;
	    RECT 15.8000 20.8000 16.2000 23.1000 ;
	    RECT 18.2000 20.8000 18.6000 24.5000 ;
	    RECT 20.6000 20.8000 21.0000 23.1000 ;
	    RECT 21.4000 20.8000 21.8000 23.1000 ;
	    RECT 23.0000 20.8000 23.4000 23.1000 ;
	    RECT 24.1000 20.8000 24.5000 23.1000 ;
	    RECT 26.2000 20.8000 26.6000 25.1000 ;
	    RECT 28.6000 20.8000 29.0000 25.1000 ;
	    RECT 29.4000 20.8000 29.8000 23.1000 ;
	    RECT 31.0000 20.8000 31.4000 23.1000 ;
	    RECT 32.6000 20.8000 33.0000 23.1000 ;
	    RECT 34.2000 20.8000 34.6000 25.0000 ;
	    RECT 37.0000 20.8000 37.4000 23.1000 ;
	    RECT 38.6000 20.8000 39.0000 23.1000 ;
	    RECT 41.4000 20.8000 41.8000 25.1000 ;
	    RECT 43.8000 20.8000 44.2000 25.0000 ;
	    RECT 46.6000 20.8000 47.0000 23.1000 ;
	    RECT 48.2000 20.8000 48.6000 23.1000 ;
	    RECT 51.0000 20.8000 51.4000 25.1000 ;
	    RECT 54.2000 20.8000 54.6000 25.1000 ;
	    RECT 55.8000 20.8000 56.2000 23.1000 ;
	    RECT 59.0000 20.8000 59.4000 25.0000 ;
	    RECT 61.8000 20.8000 62.2000 23.1000 ;
	    RECT 63.4000 20.8000 63.8000 23.1000 ;
	    RECT 66.2000 20.8000 66.6000 25.1000 ;
	    RECT 67.8000 20.8000 68.2000 25.1000 ;
	    RECT 69.9000 20.8000 70.3000 23.1000 ;
	    RECT 72.6000 20.8000 73.0000 25.1000 ;
	    RECT 74.2000 20.8000 74.6000 25.0000 ;
	    RECT 77.0000 20.8000 77.4000 23.1000 ;
	    RECT 78.6000 20.8000 79.0000 23.1000 ;
	    RECT 81.4000 20.8000 81.8000 25.1000 ;
	    RECT 83.8000 20.8000 84.2000 25.1000 ;
	    RECT 86.6000 20.8000 87.0000 23.1000 ;
	    RECT 88.2000 20.8000 88.6000 23.1000 ;
	    RECT 91.0000 20.8000 91.4000 25.0000 ;
	    RECT 92.6000 20.8000 93.0000 25.1000 ;
	    RECT 95.0000 20.8000 95.4000 23.1000 ;
	    RECT 96.6000 20.8000 97.0000 23.1000 ;
	    RECT 98.2000 20.8000 98.6000 24.5000 ;
	    RECT 100.6000 20.8000 101.0000 23.1000 ;
	    RECT 102.2000 20.8000 102.6000 23.1000 ;
	    RECT 103.8000 20.8000 104.2000 25.1000 ;
	    RECT 104.6000 20.8000 105.0000 25.1000 ;
	    RECT 106.7000 20.8000 107.1000 23.1000 ;
	    RECT 110.2000 20.8000 110.6000 24.5000 ;
	    RECT 113.4000 20.8000 113.8000 25.0000 ;
	    RECT 116.2000 20.8000 116.6000 23.1000 ;
	    RECT 117.8000 20.8000 118.2000 23.1000 ;
	    RECT 120.6000 20.8000 121.0000 25.1000 ;
	    RECT 122.2000 20.8000 122.6000 23.1000 ;
	    RECT 123.8000 20.8000 124.2000 23.1000 ;
	    RECT 125.4000 20.8000 125.8000 23.1000 ;
	    RECT 126.2000 20.8000 126.6000 25.1000 ;
	    RECT 129.7000 20.8000 130.1000 25.1000 ;
	    RECT 131.8000 20.8000 132.2000 25.1000 ;
	    RECT 134.2000 20.8000 134.6000 23.1000 ;
	    RECT 135.8000 20.8000 136.2000 23.1000 ;
	    RECT 136.9000 20.8000 137.3000 23.1000 ;
	    RECT 139.0000 20.8000 139.4000 25.1000 ;
	    RECT 140.6000 20.8000 141.0000 23.1000 ;
	    RECT 142.2000 20.8000 142.6000 25.1000 ;
	    RECT 145.0000 20.8000 145.4000 23.1000 ;
	    RECT 146.6000 20.8000 147.0000 23.1000 ;
	    RECT 149.4000 20.8000 149.8000 25.0000 ;
	    RECT 151.8000 20.8000 152.2000 24.5000 ;
	    RECT 155.0000 20.8000 155.4000 25.0000 ;
	    RECT 157.8000 20.8000 158.2000 23.1000 ;
	    RECT 159.4000 20.8000 159.8000 23.1000 ;
	    RECT 162.2000 20.8000 162.6000 25.1000 ;
	    RECT 165.4000 20.8000 165.8000 25.1000 ;
	    RECT 167.5000 20.8000 167.9000 23.1000 ;
	    RECT 169.4000 20.8000 169.8000 25.0000 ;
	    RECT 172.2000 20.8000 172.6000 23.1000 ;
	    RECT 173.8000 20.8000 174.2000 23.1000 ;
	    RECT 176.6000 20.8000 177.0000 25.1000 ;
	    RECT 178.2000 20.8000 178.6000 25.1000 ;
	    RECT 181.4000 20.8000 181.8000 23.1000 ;
	    RECT 182.2000 20.8000 182.6000 25.1000 ;
	    RECT 183.8000 20.8000 184.2000 25.1000 ;
	    RECT 185.4000 20.8000 185.8000 25.1000 ;
	    RECT 187.0000 20.8000 187.4000 25.1000 ;
	    RECT 188.6000 20.8000 189.0000 25.1000 ;
	    RECT 190.2000 20.8000 190.6000 25.0000 ;
	    RECT 193.0000 20.8000 193.4000 23.1000 ;
	    RECT 194.6000 20.8000 195.0000 23.1000 ;
	    RECT 197.4000 20.8000 197.8000 25.1000 ;
	    RECT 199.0000 20.8000 199.4000 25.1000 ;
	    RECT 201.2000 20.8000 201.6000 25.1000 ;
	    RECT 203.8000 20.8000 204.2000 24.9000 ;
	    RECT 206.2000 20.8000 206.6000 24.9000 ;
	    RECT 207.8000 20.8000 208.2000 23.1000 ;
	    RECT 208.6000 20.8000 209.0000 25.1000 ;
	    RECT 210.7000 20.8000 211.1000 23.1000 ;
	    RECT 214.2000 20.8000 214.6000 23.1000 ;
	    RECT 215.0000 20.8000 215.4000 23.1000 ;
	    RECT 216.6000 20.8000 217.0000 23.1000 ;
	    RECT 217.4000 20.8000 217.8000 23.1000 ;
	    RECT 219.0000 20.8000 219.4000 23.1000 ;
	    RECT 220.6000 20.8000 221.0000 25.1000 ;
	    RECT 221.4000 20.8000 221.8000 23.1000 ;
	    RECT 223.0000 20.8000 223.4000 23.1000 ;
	    RECT 223.8000 20.8000 224.2000 25.1000 ;
	    RECT 226.2000 20.8000 226.6000 25.1000 ;
	    RECT 228.3000 20.8000 228.7000 23.1000 ;
	    RECT 230.2000 20.8000 230.6000 24.5000 ;
	    RECT 232.6000 20.8000 233.0000 23.1000 ;
	    RECT 234.2000 20.8000 234.6000 23.1000 ;
	    RECT 235.3000 20.8000 235.7000 23.1000 ;
	    RECT 237.4000 20.8000 237.8000 25.1000 ;
	    RECT 239.0000 20.8000 239.4000 24.5000 ;
	    RECT 241.4000 20.8000 241.8000 25.1000 ;
	    RECT 243.0000 20.8000 243.4000 25.1000 ;
	    RECT 244.6000 21.1000 245.1000 24.4000 ;
	    RECT 244.7000 20.8000 245.1000 21.1000 ;
	    RECT 247.7000 20.8000 248.2000 24.4000 ;
	    RECT 250.2000 20.8000 250.6000 25.0000 ;
	    RECT 253.0000 20.8000 253.4000 23.1000 ;
	    RECT 254.6000 20.8000 255.0000 23.1000 ;
	    RECT 257.4000 20.8000 257.8000 25.1000 ;
	    RECT 259.0000 20.8000 259.4000 23.1000 ;
	    RECT 261.4000 20.8000 261.8000 25.0000 ;
	    RECT 264.2000 20.8000 264.6000 23.1000 ;
	    RECT 265.8000 20.8000 266.2000 23.1000 ;
	    RECT 268.6000 20.8000 269.0000 25.1000 ;
	    RECT 0.2000 20.2000 271.0000 20.8000 ;
	    RECT 1.4000 17.9000 1.8000 20.2000 ;
	    RECT 2.2000 15.9000 2.6000 20.2000 ;
	    RECT 5.4000 15.9000 5.8000 20.2000 ;
	    RECT 8.2000 17.9000 8.6000 20.2000 ;
	    RECT 9.8000 17.9000 10.2000 20.2000 ;
	    RECT 12.6000 16.0000 13.0000 20.2000 ;
	    RECT 15.8000 15.9000 16.2000 20.2000 ;
	    RECT 17.4000 17.9000 17.8000 20.2000 ;
	    RECT 19.0000 15.9000 19.4000 20.2000 ;
	    RECT 21.8000 17.9000 22.2000 20.2000 ;
	    RECT 23.4000 17.9000 23.8000 20.2000 ;
	    RECT 26.2000 16.0000 26.6000 20.2000 ;
	    RECT 28.6000 16.5000 29.0000 20.2000 ;
	    RECT 31.0000 16.0000 31.4000 20.2000 ;
	    RECT 33.8000 17.9000 34.2000 20.2000 ;
	    RECT 35.4000 17.9000 35.8000 20.2000 ;
	    RECT 38.2000 15.9000 38.6000 20.2000 ;
	    RECT 40.9000 15.9000 41.3000 20.2000 ;
	    RECT 44.6000 15.9000 45.0000 20.2000 ;
	    RECT 46.2000 17.9000 46.6000 20.2000 ;
	    RECT 47.0000 17.9000 47.4000 20.2000 ;
	    RECT 50.2000 15.9000 50.6000 20.2000 ;
	    RECT 51.8000 16.6000 52.3000 20.2000 ;
	    RECT 54.9000 19.9000 55.3000 20.2000 ;
	    RECT 54.9000 16.6000 55.4000 19.9000 ;
	    RECT 59.8000 16.5000 60.2000 20.2000 ;
	    RECT 61.4000 17.9000 61.8000 20.2000 ;
	    RECT 63.0000 17.9000 63.4000 20.2000 ;
	    RECT 64.1000 17.9000 64.5000 20.2000 ;
	    RECT 66.2000 15.9000 66.6000 20.2000 ;
	    RECT 67.0000 17.9000 67.4000 20.2000 ;
	    RECT 68.6000 15.9000 69.0000 20.2000 ;
	    RECT 70.7000 17.9000 71.1000 20.2000 ;
	    RECT 72.6000 16.5000 73.0000 20.2000 ;
	    RECT 76.6000 17.9000 77.0000 20.2000 ;
	    RECT 77.4000 15.9000 77.8000 20.2000 ;
	    RECT 79.0000 15.9000 79.4000 20.2000 ;
	    RECT 80.6000 15.9000 81.0000 20.2000 ;
	    RECT 82.2000 15.9000 82.6000 20.2000 ;
	    RECT 83.8000 15.9000 84.2000 20.2000 ;
	    RECT 86.2000 15.9000 86.6000 20.2000 ;
	    RECT 87.8000 16.5000 88.2000 20.2000 ;
	    RECT 90.5000 17.9000 90.9000 20.2000 ;
	    RECT 92.6000 15.9000 93.0000 20.2000 ;
	    RECT 95.0000 15.9000 95.4000 20.2000 ;
	    RECT 96.1000 17.9000 96.5000 20.2000 ;
	    RECT 98.2000 15.9000 98.6000 20.2000 ;
	    RECT 99.8000 17.9000 100.2000 20.2000 ;
	    RECT 100.6000 17.9000 101.0000 20.2000 ;
	    RECT 103.0000 16.5000 103.4000 20.2000 ;
	    RECT 105.4000 17.9000 105.8000 20.2000 ;
	    RECT 107.0000 17.9000 107.4000 20.2000 ;
	    RECT 109.7000 17.9000 110.1000 20.2000 ;
	    RECT 111.8000 15.9000 112.2000 20.2000 ;
	    RECT 112.6000 15.9000 113.0000 20.2000 ;
	    RECT 115.8000 17.9000 116.2000 20.2000 ;
	    RECT 116.6000 15.9000 117.0000 20.2000 ;
	    RECT 119.0000 17.9000 119.4000 20.2000 ;
	    RECT 120.6000 17.9000 121.0000 20.2000 ;
	    RECT 122.2000 17.9000 122.6000 20.2000 ;
	    RECT 123.8000 17.9000 124.2000 20.2000 ;
	    RECT 125.4000 15.9000 125.8000 20.2000 ;
	    RECT 128.2000 17.9000 128.6000 20.2000 ;
	    RECT 129.8000 17.9000 130.2000 20.2000 ;
	    RECT 132.6000 16.0000 133.0000 20.2000 ;
	    RECT 134.2000 17.9000 134.6000 20.2000 ;
	    RECT 135.8000 15.9000 136.2000 20.2000 ;
	    RECT 139.0000 16.6000 139.5000 20.2000 ;
	    RECT 142.1000 19.9000 142.5000 20.2000 ;
	    RECT 142.1000 16.6000 142.6000 19.9000 ;
	    RECT 143.8000 17.9000 144.2000 20.2000 ;
	    RECT 145.4000 15.9000 145.8000 20.2000 ;
	    RECT 147.8000 15.9000 148.2000 20.2000 ;
	    RECT 149.4000 15.9000 149.8000 20.2000 ;
	    RECT 151.0000 15.9000 151.4000 20.2000 ;
	    RECT 152.6000 15.9000 153.0000 20.2000 ;
	    RECT 154.2000 15.9000 154.6000 20.2000 ;
	    RECT 155.0000 15.9000 155.4000 20.2000 ;
	    RECT 156.6000 16.5000 157.0000 20.2000 ;
	    RECT 158.2000 17.9000 158.6000 20.2000 ;
	    RECT 161.4000 15.9000 161.8000 20.2000 ;
	    RECT 163.8000 15.9000 164.2000 20.2000 ;
	    RECT 165.4000 15.9000 165.8000 20.2000 ;
	    RECT 167.0000 15.9000 167.4000 20.2000 ;
	    RECT 168.6000 15.9000 169.0000 20.2000 ;
	    RECT 170.2000 15.9000 170.6000 20.2000 ;
	    RECT 171.8000 16.5000 172.2000 20.2000 ;
	    RECT 174.2000 15.9000 174.6000 20.2000 ;
	    RECT 177.0000 17.9000 177.4000 20.2000 ;
	    RECT 178.6000 17.9000 179.0000 20.2000 ;
	    RECT 181.4000 16.0000 181.8000 20.2000 ;
	    RECT 183.0000 17.9000 183.4000 20.2000 ;
	    RECT 184.6000 15.9000 185.0000 20.2000 ;
	    RECT 188.6000 15.9000 189.0000 20.2000 ;
	    RECT 189.4000 17.9000 189.8000 20.2000 ;
	    RECT 191.0000 16.1000 191.4000 20.2000 ;
	    RECT 192.6000 15.9000 193.0000 20.2000 ;
	    RECT 194.7000 17.9000 195.1000 20.2000 ;
	    RECT 196.6000 16.0000 197.0000 20.2000 ;
	    RECT 199.4000 17.9000 199.8000 20.2000 ;
	    RECT 201.0000 17.9000 201.4000 20.2000 ;
	    RECT 203.8000 15.9000 204.2000 20.2000 ;
	    RECT 206.0000 15.9000 206.4000 20.2000 ;
	    RECT 208.6000 16.1000 209.0000 20.2000 ;
	    RECT 210.2000 15.9000 210.6000 20.2000 ;
	    RECT 213.7000 17.9000 214.1000 20.2000 ;
	    RECT 215.8000 15.9000 216.2000 20.2000 ;
	    RECT 216.6000 17.9000 217.0000 20.2000 ;
	    RECT 218.2000 17.9000 218.6000 20.2000 ;
	    RECT 219.0000 17.9000 219.4000 20.2000 ;
	    RECT 220.6000 16.1000 221.0000 20.2000 ;
	    RECT 223.8000 15.9000 224.2000 20.2000 ;
	    RECT 224.6000 17.9000 225.0000 20.2000 ;
	    RECT 226.2000 17.9000 226.6000 20.2000 ;
	    RECT 227.0000 15.9000 227.4000 20.2000 ;
	    RECT 229.4000 17.9000 229.8000 20.2000 ;
	    RECT 231.0000 17.9000 231.4000 20.2000 ;
	    RECT 231.8000 17.9000 232.2000 20.2000 ;
	    RECT 235.8000 16.5000 236.2000 20.2000 ;
	    RECT 237.7000 17.9000 238.1000 20.2000 ;
	    RECT 239.8000 15.9000 240.2000 20.2000 ;
	    RECT 242.2000 15.9000 242.6000 20.2000 ;
	    RECT 243.0000 17.9000 243.4000 20.2000 ;
	    RECT 244.6000 17.9000 245.0000 20.2000 ;
	    RECT 245.4000 15.9000 245.8000 20.2000 ;
	    RECT 247.5000 17.9000 247.9000 20.2000 ;
	    RECT 249.4000 15.9000 249.8000 20.2000 ;
	    RECT 250.2000 15.9000 250.6000 20.2000 ;
	    RECT 253.4000 15.9000 253.8000 20.2000 ;
	    RECT 255.0000 17.9000 255.4000 20.2000 ;
	    RECT 256.6000 17.9000 257.0000 20.2000 ;
	    RECT 259.0000 16.5000 259.4000 20.2000 ;
	    RECT 261.4000 16.0000 261.8000 20.2000 ;
	    RECT 264.2000 17.9000 264.6000 20.2000 ;
	    RECT 265.8000 17.9000 266.2000 20.2000 ;
	    RECT 268.6000 15.9000 269.0000 20.2000 ;
	    RECT 1.4000 0.8000 1.8000 4.5000 ;
	    RECT 3.8000 0.8000 4.2000 4.5000 ;
	    RECT 5.4000 0.8000 5.8000 3.1000 ;
	    RECT 7.0000 0.8000 7.4000 5.1000 ;
	    RECT 10.2000 0.8000 10.6000 5.1000 ;
	    RECT 13.0000 0.8000 13.4000 3.1000 ;
	    RECT 14.6000 0.8000 15.0000 3.1000 ;
	    RECT 17.4000 0.8000 17.8000 5.0000 ;
	    RECT 19.8000 0.8000 20.2000 4.5000 ;
	    RECT 23.0000 0.8000 23.4000 5.1000 ;
	    RECT 24.6000 0.8000 25.0000 3.1000 ;
	    RECT 26.2000 0.8000 26.6000 5.0000 ;
	    RECT 29.0000 0.8000 29.4000 3.1000 ;
	    RECT 30.6000 0.8000 31.0000 3.1000 ;
	    RECT 33.4000 0.8000 33.8000 5.1000 ;
	    RECT 35.8000 0.8000 36.2000 4.5000 ;
	    RECT 39.0000 0.8000 39.4000 5.1000 ;
	    RECT 40.6000 0.8000 41.0000 3.1000 ;
	    RECT 42.2000 0.8000 42.6000 5.0000 ;
	    RECT 45.0000 0.8000 45.4000 3.1000 ;
	    RECT 46.6000 0.8000 47.0000 3.1000 ;
	    RECT 49.4000 0.8000 49.8000 5.1000 ;
	    RECT 51.8000 0.8000 52.2000 4.5000 ;
	    RECT 54.2000 1.1000 54.7000 4.4000 ;
	    RECT 54.3000 0.8000 54.7000 1.1000 ;
	    RECT 57.3000 0.8000 57.8000 4.4000 ;
	    RECT 60.6000 0.8000 61.0000 5.1000 ;
	    RECT 63.8000 0.8000 64.2000 3.1000 ;
	    RECT 65.4000 0.8000 65.9000 4.4000 ;
	    RECT 68.5000 1.1000 69.0000 4.4000 ;
	    RECT 71.0000 1.1000 71.5000 4.4000 ;
	    RECT 68.5000 0.8000 68.9000 1.1000 ;
	    RECT 71.1000 0.8000 71.5000 1.1000 ;
	    RECT 74.1000 0.8000 74.6000 4.4000 ;
	    RECT 77.4000 0.8000 77.8000 5.1000 ;
	    RECT 78.2000 0.8000 78.6000 3.1000 ;
	    RECT 79.8000 0.8000 80.2000 5.1000 ;
	    RECT 83.0000 0.8000 83.4000 5.1000 ;
	    RECT 84.6000 0.8000 85.0000 4.5000 ;
	    RECT 88.6000 0.8000 89.0000 3.1000 ;
	    RECT 89.4000 0.8000 89.8000 3.1000 ;
	    RECT 91.0000 0.8000 91.4000 3.1000 ;
	    RECT 91.8000 0.8000 92.2000 3.1000 ;
	    RECT 93.4000 0.8000 93.8000 3.1000 ;
	    RECT 94.2000 0.8000 94.6000 3.1000 ;
	    RECT 95.8000 0.8000 96.2000 4.9000 ;
	    RECT 99.0000 0.8000 99.4000 4.5000 ;
	    RECT 102.2000 0.8000 102.6000 5.1000 ;
	    RECT 103.0000 0.8000 103.4000 3.1000 ;
	    RECT 104.6000 0.8000 105.0000 3.1000 ;
	    RECT 105.4000 0.8000 105.8000 5.1000 ;
	    RECT 108.6000 0.8000 109.0000 3.1000 ;
	    RECT 111.8000 0.8000 112.3000 4.4000 ;
	    RECT 114.9000 1.1000 115.4000 4.4000 ;
	    RECT 114.9000 0.8000 115.3000 1.1000 ;
	    RECT 116.6000 0.8000 117.0000 3.1000 ;
	    RECT 118.2000 0.8000 118.6000 3.1000 ;
	    RECT 119.8000 0.8000 120.2000 3.1000 ;
	    RECT 120.6000 0.8000 121.0000 5.1000 ;
	    RECT 123.0000 0.8000 123.4000 3.1000 ;
	    RECT 124.6000 0.8000 125.0000 3.1000 ;
	    RECT 126.2000 0.8000 126.7000 4.4000 ;
	    RECT 129.3000 1.1000 129.8000 4.4000 ;
	    RECT 129.3000 0.8000 129.7000 1.1000 ;
	    RECT 131.8000 0.8000 132.2000 4.5000 ;
	    RECT 134.2000 0.8000 134.6000 5.1000 ;
	    RECT 136.6000 0.8000 137.0000 3.1000 ;
	    RECT 138.2000 0.8000 138.6000 3.1000 ;
	    RECT 139.8000 0.8000 140.2000 3.1000 ;
	    RECT 140.6000 0.8000 141.0000 3.1000 ;
	    RECT 142.2000 0.8000 142.6000 3.1000 ;
	    RECT 143.8000 0.8000 144.2000 5.1000 ;
	    RECT 146.6000 0.8000 147.0000 3.1000 ;
	    RECT 148.2000 0.8000 148.6000 3.1000 ;
	    RECT 151.0000 0.8000 151.4000 5.0000 ;
	    RECT 153.4000 0.8000 153.9000 4.4000 ;
	    RECT 156.5000 1.1000 157.0000 4.4000 ;
	    RECT 156.5000 0.8000 156.9000 1.1000 ;
	    RECT 160.6000 0.8000 161.0000 5.1000 ;
	    RECT 163.4000 0.8000 163.8000 3.1000 ;
	    RECT 165.0000 0.8000 165.4000 3.1000 ;
	    RECT 167.8000 0.8000 168.2000 5.0000 ;
	    RECT 170.7000 0.8000 171.1000 5.1000 ;
	    RECT 173.4000 0.8000 173.8000 5.1000 ;
	    RECT 176.2000 0.8000 176.6000 3.1000 ;
	    RECT 177.8000 0.8000 178.2000 3.1000 ;
	    RECT 180.6000 0.8000 181.0000 5.0000 ;
	    RECT 183.0000 0.8000 183.4000 4.5000 ;
	    RECT 185.4000 0.8000 185.8000 5.1000 ;
	    RECT 188.2000 0.8000 188.6000 3.1000 ;
	    RECT 189.8000 0.8000 190.2000 3.1000 ;
	    RECT 192.6000 0.8000 193.0000 5.0000 ;
	    RECT 194.2000 0.8000 194.6000 3.1000 ;
	    RECT 195.8000 0.8000 196.2000 5.1000 ;
	    RECT 199.0000 0.8000 199.4000 4.5000 ;
	    RECT 202.2000 0.8000 202.6000 5.1000 ;
	    RECT 203.8000 0.8000 204.2000 3.1000 ;
	    RECT 205.4000 0.8000 205.8000 5.0000 ;
	    RECT 208.2000 0.8000 208.6000 3.1000 ;
	    RECT 209.8000 0.8000 210.2000 3.1000 ;
	    RECT 212.6000 0.8000 213.0000 5.1000 ;
	    RECT 216.6000 0.8000 217.0000 5.1000 ;
	    RECT 218.2000 0.8000 218.6000 5.1000 ;
	    RECT 221.0000 0.8000 221.4000 3.1000 ;
	    RECT 222.6000 0.8000 223.0000 3.1000 ;
	    RECT 225.4000 0.8000 225.8000 5.0000 ;
	    RECT 227.0000 0.8000 227.4000 3.1000 ;
	    RECT 229.2000 0.8000 229.6000 5.1000 ;
	    RECT 231.8000 0.8000 232.2000 4.9000 ;
	    RECT 233.4000 0.8000 233.8000 3.1000 ;
	    RECT 236.6000 0.8000 237.0000 5.1000 ;
	    RECT 238.2000 0.8000 238.6000 3.1000 ;
	    RECT 240.6000 0.8000 241.0000 5.1000 ;
	    RECT 241.4000 0.8000 241.8000 3.1000 ;
	    RECT 243.0000 0.8000 243.4000 5.1000 ;
	    RECT 246.2000 0.8000 246.6000 5.1000 ;
	    RECT 247.0000 0.8000 247.4000 3.1000 ;
	    RECT 248.6000 0.8000 249.0000 3.1000 ;
	    RECT 249.4000 0.8000 249.8000 3.1000 ;
	    RECT 251.8000 0.8000 252.2000 4.5000 ;
	    RECT 255.8000 0.8000 256.2000 5.1000 ;
	    RECT 257.4000 0.8000 257.8000 3.1000 ;
	    RECT 258.2000 0.8000 258.6000 5.1000 ;
	    RECT 260.6000 0.8000 261.0000 3.1000 ;
	    RECT 262.2000 0.8000 262.6000 3.1000 ;
	    RECT 263.8000 0.8000 264.2000 4.5000 ;
	    RECT 267.0000 0.8000 267.4000 4.5000 ;
	    RECT 268.6000 0.8000 269.0000 3.1000 ;
	    RECT 0.2000 0.2000 271.0000 0.8000 ;
         LAYER metal2 ;
	    RECT 57.6000 180.3000 59.2000 180.7000 ;
	    RECT 160.0000 180.3000 161.6000 180.7000 ;
	    RECT 57.6000 160.3000 59.2000 160.7000 ;
	    RECT 160.0000 160.3000 161.6000 160.7000 ;
	    RECT 57.6000 140.3000 59.2000 140.7000 ;
	    RECT 160.0000 140.3000 161.6000 140.7000 ;
	    RECT 57.6000 120.3000 59.2000 120.7000 ;
	    RECT 160.0000 120.3000 161.6000 120.7000 ;
	    RECT 57.6000 100.3000 59.2000 100.7000 ;
	    RECT 160.0000 100.3000 161.6000 100.7000 ;
	    RECT 57.6000 80.3000 59.2000 80.7000 ;
	    RECT 160.0000 80.3000 161.6000 80.7000 ;
	    RECT 57.6000 60.3000 59.2000 60.7000 ;
	    RECT 160.0000 60.3000 161.6000 60.7000 ;
	    RECT 57.6000 40.3000 59.2000 40.7000 ;
	    RECT 160.0000 40.3000 161.6000 40.7000 ;
	    RECT 57.6000 20.3000 59.2000 20.7000 ;
	    RECT 160.0000 20.3000 161.6000 20.7000 ;
	    RECT 57.6000 0.3000 59.2000 0.7000 ;
	    RECT 160.0000 0.3000 161.6000 0.7000 ;
         LAYER metal3 ;
	    RECT 57.6000 180.3000 59.2000 180.7000 ;
	    RECT 160.0000 180.3000 161.6000 180.7000 ;
	    RECT 57.6000 160.3000 59.2000 160.7000 ;
	    RECT 160.0000 160.3000 161.6000 160.7000 ;
	    RECT 57.6000 140.3000 59.2000 140.7000 ;
	    RECT 160.0000 140.3000 161.6000 140.7000 ;
	    RECT 57.6000 120.3000 59.2000 120.7000 ;
	    RECT 160.0000 120.3000 161.6000 120.7000 ;
	    RECT 57.6000 100.3000 59.2000 100.7000 ;
	    RECT 160.0000 100.3000 161.6000 100.7000 ;
	    RECT 57.6000 80.3000 59.2000 80.7000 ;
	    RECT 160.0000 80.3000 161.6000 80.7000 ;
	    RECT 57.6000 60.3000 59.2000 60.7000 ;
	    RECT 160.0000 60.3000 161.6000 60.7000 ;
	    RECT 57.6000 40.3000 59.2000 40.7000 ;
	    RECT 160.0000 40.3000 161.6000 40.7000 ;
	    RECT 57.6000 20.3000 59.2000 20.7000 ;
	    RECT 160.0000 20.3000 161.6000 20.7000 ;
	    RECT 57.6000 0.3000 59.2000 0.7000 ;
	    RECT 160.0000 0.3000 161.6000 0.7000 ;
         LAYER metal4 ;
	    RECT 57.6000 180.3000 59.2000 180.7000 ;
	    RECT 160.0000 180.3000 161.6000 180.7000 ;
	    RECT 57.6000 160.3000 59.2000 160.7000 ;
	    RECT 160.0000 160.3000 161.6000 160.7000 ;
	    RECT 57.6000 140.3000 59.2000 140.7000 ;
	    RECT 160.0000 140.3000 161.6000 140.7000 ;
	    RECT 57.6000 120.3000 59.2000 120.7000 ;
	    RECT 160.0000 120.3000 161.6000 120.7000 ;
	    RECT 57.6000 100.3000 59.2000 100.7000 ;
	    RECT 160.0000 100.3000 161.6000 100.7000 ;
	    RECT 57.6000 80.3000 59.2000 80.7000 ;
	    RECT 160.0000 80.3000 161.6000 80.7000 ;
	    RECT 57.6000 60.3000 59.2000 60.7000 ;
	    RECT 160.0000 60.3000 161.6000 60.7000 ;
	    RECT 57.6000 40.3000 59.2000 40.7000 ;
	    RECT 160.0000 40.3000 161.6000 40.7000 ;
	    RECT 57.6000 20.3000 59.2000 20.7000 ;
	    RECT 160.0000 20.3000 161.6000 20.7000 ;
	    RECT 57.6000 0.3000 59.2000 0.7000 ;
	    RECT 160.0000 0.3000 161.6000 0.7000 ;
         LAYER metal5 ;
	    RECT 57.6000 180.7000 58.2000 180.8000 ;
	    RECT 58.6000 180.7000 59.2000 180.8000 ;
	    RECT 57.6000 180.2000 59.2000 180.7000 ;
	    RECT 160.0000 180.7000 160.6000 180.8000 ;
	    RECT 161.0000 180.7000 161.6000 180.8000 ;
	    RECT 160.0000 180.2000 161.6000 180.7000 ;
	    RECT 57.6000 160.7000 58.2000 160.8000 ;
	    RECT 58.6000 160.7000 59.2000 160.8000 ;
	    RECT 57.6000 160.2000 59.2000 160.7000 ;
	    RECT 160.0000 160.7000 160.6000 160.8000 ;
	    RECT 161.0000 160.7000 161.6000 160.8000 ;
	    RECT 160.0000 160.2000 161.6000 160.7000 ;
	    RECT 57.6000 140.7000 58.2000 140.8000 ;
	    RECT 58.6000 140.7000 59.2000 140.8000 ;
	    RECT 57.6000 140.2000 59.2000 140.7000 ;
	    RECT 160.0000 140.7000 160.6000 140.8000 ;
	    RECT 161.0000 140.7000 161.6000 140.8000 ;
	    RECT 160.0000 140.2000 161.6000 140.7000 ;
	    RECT 57.6000 120.7000 58.2000 120.8000 ;
	    RECT 58.6000 120.7000 59.2000 120.8000 ;
	    RECT 57.6000 120.2000 59.2000 120.7000 ;
	    RECT 160.0000 120.7000 160.6000 120.8000 ;
	    RECT 161.0000 120.7000 161.6000 120.8000 ;
	    RECT 160.0000 120.2000 161.6000 120.7000 ;
	    RECT 57.6000 100.7000 58.2000 100.8000 ;
	    RECT 58.6000 100.7000 59.2000 100.8000 ;
	    RECT 57.6000 100.2000 59.2000 100.7000 ;
	    RECT 160.0000 100.7000 160.6000 100.8000 ;
	    RECT 161.0000 100.7000 161.6000 100.8000 ;
	    RECT 160.0000 100.2000 161.6000 100.7000 ;
	    RECT 57.6000 80.7000 58.2000 80.8000 ;
	    RECT 58.6000 80.7000 59.2000 80.8000 ;
	    RECT 57.6000 80.2000 59.2000 80.7000 ;
	    RECT 160.0000 80.7000 160.6000 80.8000 ;
	    RECT 161.0000 80.7000 161.6000 80.8000 ;
	    RECT 160.0000 80.2000 161.6000 80.7000 ;
	    RECT 57.6000 60.7000 58.2000 60.8000 ;
	    RECT 58.6000 60.7000 59.2000 60.8000 ;
	    RECT 57.6000 60.2000 59.2000 60.7000 ;
	    RECT 160.0000 60.7000 160.6000 60.8000 ;
	    RECT 161.0000 60.7000 161.6000 60.8000 ;
	    RECT 160.0000 60.2000 161.6000 60.7000 ;
	    RECT 57.6000 40.7000 58.2000 40.8000 ;
	    RECT 58.6000 40.7000 59.2000 40.8000 ;
	    RECT 57.6000 40.2000 59.2000 40.7000 ;
	    RECT 160.0000 40.7000 160.6000 40.8000 ;
	    RECT 161.0000 40.7000 161.6000 40.8000 ;
	    RECT 160.0000 40.2000 161.6000 40.7000 ;
	    RECT 57.6000 20.7000 58.2000 20.8000 ;
	    RECT 58.6000 20.7000 59.2000 20.8000 ;
	    RECT 57.6000 20.2000 59.2000 20.7000 ;
	    RECT 160.0000 20.7000 160.6000 20.8000 ;
	    RECT 161.0000 20.7000 161.6000 20.8000 ;
	    RECT 160.0000 20.2000 161.6000 20.7000 ;
	    RECT 57.6000 0.7000 58.2000 0.8000 ;
	    RECT 58.6000 0.7000 59.2000 0.8000 ;
	    RECT 57.6000 0.2000 59.2000 0.7000 ;
	    RECT 160.0000 0.7000 160.6000 0.8000 ;
	    RECT 161.0000 0.7000 161.6000 0.8000 ;
	    RECT 160.0000 0.2000 161.6000 0.7000 ;
         LAYER metal6 ;
	    RECT 57.6000 -3.0000 59.2000 183.0000 ;
	    RECT 160.0000 -3.0000 161.6000 183.0000 ;
      END
   END vdd
   PIN gnd
      PORT
         LAYER metal1 ;
	    RECT 3.0000 174.4000 3.4000 175.2000 ;
	    RECT 4.6000 174.4000 5.0000 175.2000 ;
	    RECT 7.8000 173.4000 8.2000 174.2000 ;
	    RECT 10.2000 173.4000 10.6000 174.2000 ;
	    RECT 12.6000 173.4000 13.0000 174.2000 ;
	    RECT 29.4000 173.4000 29.8000 174.2000 ;
	    RECT 0.6000 170.8000 1.0000 172.1000 ;
	    RECT 3.0000 170.8000 3.4000 172.7000 ;
	    RECT 7.8000 170.8000 8.2000 173.1000 ;
	    RECT 10.2000 170.8000 10.6000 173.1000 ;
	    RECT 11.8000 170.8000 12.2000 172.1000 ;
	    RECT 12.6000 170.8000 13.0000 173.1000 ;
	    RECT 16.6000 172.4000 17.0000 173.2000 ;
	    RECT 23.0000 173.1000 23.4000 173.2000 ;
	    RECT 15.8000 170.8000 16.2000 172.1000 ;
	    RECT 16.6000 170.8000 17.0000 172.1000 ;
	    RECT 18.2000 170.8000 18.6000 173.1000 ;
	    RECT 21.2000 170.8000 21.6000 173.1000 ;
	    RECT 23.0000 172.8000 24.1000 173.1000 ;
	    RECT 23.0000 172.4000 23.4000 172.8000 ;
	    RECT 23.8000 172.1000 24.1000 172.8000 ;
	    RECT 23.0000 170.8000 23.4000 172.1000 ;
	    RECT 23.8000 170.8000 24.2000 172.1000 ;
	    RECT 25.4000 170.8000 25.8000 172.1000 ;
	    RECT 26.2000 170.8000 26.6000 172.1000 ;
	    RECT 29.4000 170.8000 29.8000 173.1000 ;
	    RECT 30.2000 170.8000 30.6000 172.1000 ;
	    RECT 31.8000 170.8000 32.2000 172.9000 ;
	    RECT 33.4000 172.4000 33.8000 173.2000 ;
	    RECT 33.4000 170.8000 33.8000 172.1000 ;
	    RECT 36.6000 170.8000 37.0000 173.1000 ;
	    RECT 37.4000 172.4000 37.8000 173.2000 ;
	    RECT 37.4000 170.8000 37.8000 172.1000 ;
	    RECT 40.6000 170.8000 41.0000 173.1000 ;
	    RECT 41.4000 172.4000 41.8000 173.2000 ;
	    RECT 41.4000 172.1000 41.7000 172.4000 ;
	    RECT 41.4000 170.8000 41.8000 172.1000 ;
	    RECT 44.6000 170.8000 45.0000 173.1000 ;
	    RECT 45.4000 170.8000 45.8000 173.1000 ;
	    RECT 48.6000 172.4000 49.0000 173.2000 ;
	    RECT 48.6000 170.8000 49.0000 172.1000 ;
	    RECT 50.2000 170.8000 50.6000 173.1000 ;
	    RECT 52.6000 170.8000 53.0000 173.0000 ;
	    RECT 55.4000 170.8000 55.8000 172.1000 ;
	    RECT 57.0000 170.8000 57.5000 172.1000 ;
	    RECT 59.8000 170.8000 60.2000 173.1000 ;
	    RECT 63.8000 170.8000 64.2000 173.1000 ;
	    RECT 66.5000 170.8000 67.0000 172.1000 ;
	    RECT 68.2000 170.8000 68.6000 172.1000 ;
	    RECT 71.0000 170.8000 71.4000 173.0000 ;
	    RECT 73.4000 170.8000 73.8000 173.1000 ;
	    RECT 75.8000 170.8000 76.2000 173.1000 ;
	    RECT 78.2000 170.8000 78.6000 173.1000 ;
	    RECT 80.6000 170.8000 81.0000 173.1000 ;
	    RECT 83.3000 170.8000 83.8000 172.1000 ;
	    RECT 85.0000 170.8000 85.4000 172.1000 ;
	    RECT 87.8000 170.8000 88.2000 173.0000 ;
	    RECT 89.4000 170.8000 89.8000 172.1000 ;
	    RECT 91.0000 170.8000 91.4000 172.1000 ;
	    RECT 92.6000 170.8000 93.0000 172.1000 ;
	    RECT 94.2000 170.8000 94.6000 173.1000 ;
	    RECT 96.6000 170.8000 97.0000 173.1000 ;
	    RECT 99.0000 170.8000 99.4000 173.1000 ;
	    RECT 101.7000 170.8000 102.2000 172.1000 ;
	    RECT 103.4000 170.8000 103.8000 172.1000 ;
	    RECT 106.2000 170.8000 106.6000 173.0000 ;
	    RECT 108.6000 170.8000 109.0000 173.1000 ;
	    RECT 112.6000 170.8000 113.0000 173.1000 ;
	    RECT 115.0000 170.8000 115.4000 173.0000 ;
	    RECT 117.8000 170.8000 118.2000 172.1000 ;
	    RECT 119.4000 170.8000 119.9000 172.1000 ;
	    RECT 122.2000 170.8000 122.6000 173.1000 ;
	    RECT 124.6000 170.8000 125.0000 173.1000 ;
	    RECT 126.2000 170.8000 126.6000 172.1000 ;
	    RECT 127.8000 170.8000 128.2000 172.1000 ;
	    RECT 129.4000 170.8000 129.8000 172.1000 ;
	    RECT 131.0000 170.8000 131.4000 173.1000 ;
	    RECT 133.4000 170.8000 133.8000 173.1000 ;
	    RECT 136.1000 170.8000 136.6000 172.1000 ;
	    RECT 137.8000 170.8000 138.2000 172.1000 ;
	    RECT 140.6000 170.8000 141.0000 173.0000 ;
	    RECT 143.0000 170.8000 143.4000 173.1000 ;
	    RECT 145.4000 170.8000 145.8000 173.1000 ;
	    RECT 147.8000 170.8000 148.2000 173.1000 ;
	    RECT 150.2000 170.8000 150.6000 173.1000 ;
	    RECT 152.6000 170.8000 153.0000 173.1000 ;
	    RECT 155.0000 170.8000 155.4000 173.0000 ;
	    RECT 157.8000 170.8000 158.2000 172.1000 ;
	    RECT 159.4000 170.8000 159.9000 172.1000 ;
	    RECT 162.2000 170.8000 162.6000 173.1000 ;
	    RECT 165.4000 170.8000 165.8000 172.1000 ;
	    RECT 167.8000 170.8000 168.2000 173.1000 ;
	    RECT 170.2000 170.8000 170.6000 173.1000 ;
	    RECT 172.6000 170.8000 173.0000 173.1000 ;
	    RECT 175.0000 170.8000 175.4000 173.1000 ;
	    RECT 177.7000 170.8000 178.2000 172.1000 ;
	    RECT 179.4000 170.8000 179.8000 172.1000 ;
	    RECT 182.2000 170.8000 182.6000 173.0000 ;
	    RECT 183.8000 170.8000 184.2000 172.1000 ;
	    RECT 185.4000 170.8000 185.8000 172.1000 ;
	    RECT 187.0000 170.8000 187.4000 172.1000 ;
	    RECT 188.6000 170.8000 189.0000 173.1000 ;
	    RECT 191.0000 170.8000 191.4000 173.1000 ;
	    RECT 193.7000 170.8000 194.2000 172.1000 ;
	    RECT 195.4000 170.8000 195.8000 172.1000 ;
	    RECT 198.2000 170.8000 198.6000 173.0000 ;
	    RECT 200.6000 170.8000 201.0000 172.7000 ;
	    RECT 203.3000 170.8000 203.7000 173.1000 ;
	    RECT 205.4000 170.8000 205.8000 172.1000 ;
	    RECT 207.0000 170.8000 207.4000 173.1000 ;
	    RECT 209.7000 170.8000 210.2000 172.1000 ;
	    RECT 211.4000 170.8000 211.8000 172.1000 ;
	    RECT 214.2000 170.8000 214.6000 173.0000 ;
	    RECT 217.4000 170.8000 217.8000 172.1000 ;
	    RECT 219.0000 170.8000 219.4000 172.1000 ;
	    RECT 220.6000 170.8000 221.0000 172.7000 ;
	    RECT 224.6000 170.8000 225.0000 173.1000 ;
	    RECT 225.7000 170.8000 226.1000 173.1000 ;
	    RECT 227.8000 170.8000 228.2000 172.1000 ;
	    RECT 229.4000 170.8000 229.8000 173.1000 ;
	    RECT 232.1000 170.8000 232.6000 172.1000 ;
	    RECT 233.8000 170.8000 234.2000 172.1000 ;
	    RECT 236.6000 170.8000 237.0000 173.0000 ;
	    RECT 238.2000 170.8000 238.6000 173.1000 ;
	    RECT 240.6000 170.8000 241.0000 172.1000 ;
	    RECT 242.2000 170.8000 242.6000 172.1000 ;
	    RECT 243.0000 170.8000 243.4000 172.1000 ;
	    RECT 244.6000 170.8000 245.0000 172.1000 ;
	    RECT 246.2000 170.8000 246.6000 172.1000 ;
	    RECT 247.0000 170.8000 247.4000 172.1000 ;
	    RECT 248.6000 170.8000 249.0000 172.1000 ;
	    RECT 250.7000 170.8000 251.1000 173.0000 ;
	    RECT 252.6000 170.8000 253.0000 172.1000 ;
	    RECT 254.2000 170.8000 254.6000 172.1000 ;
	    RECT 255.0000 170.8000 255.4000 172.1000 ;
	    RECT 257.4000 170.8000 257.8000 173.1000 ;
	    RECT 260.1000 170.8000 260.6000 172.1000 ;
	    RECT 261.8000 170.8000 262.2000 172.1000 ;
	    RECT 264.6000 170.8000 265.0000 173.0000 ;
	    RECT 267.0000 170.8000 267.4000 172.1000 ;
	    RECT 268.6000 170.8000 269.0000 173.1000 ;
	    RECT 0.2000 170.2000 271.0000 170.8000 ;
	    RECT 1.4000 167.9000 1.8000 170.2000 ;
	    RECT 4.6000 168.3000 5.0000 170.2000 ;
	    RECT 6.2000 168.9000 6.6000 170.2000 ;
	    RECT 6.2000 167.8000 6.6000 168.6000 ;
	    RECT 7.8000 166.9000 8.2000 170.2000 ;
	    RECT 11.2000 167.9000 11.6000 170.2000 ;
	    RECT 14.2000 167.9000 14.6000 170.2000 ;
	    RECT 15.8000 168.9000 16.2000 170.2000 ;
	    RECT 17.4000 168.9000 17.8000 170.2000 ;
	    RECT 18.2000 168.9000 18.6000 170.2000 ;
	    RECT 15.8000 167.8000 16.2000 168.6000 ;
	    RECT 18.2000 167.8000 18.6000 168.6000 ;
	    RECT 19.8000 167.9000 20.2000 170.2000 ;
	    RECT 22.8000 167.9000 23.2000 170.2000 ;
	    RECT 23.8000 168.9000 24.2000 170.2000 ;
	    RECT 25.4000 168.9000 25.8000 170.2000 ;
	    RECT 27.0000 168.9000 27.4000 170.2000 ;
	    RECT 27.0000 168.1000 27.4000 168.6000 ;
	    RECT 27.8000 168.1000 28.2000 170.2000 ;
	    RECT 31.0000 168.9000 31.4000 170.2000 ;
	    RECT 27.0000 167.8000 28.2000 168.1000 ;
	    RECT 34.2000 167.9000 34.6000 170.2000 ;
	    RECT 35.8000 168.3000 36.2000 170.2000 ;
	    RECT 38.2000 168.9000 38.6000 170.2000 ;
	    RECT 39.8000 167.9000 40.2000 170.2000 ;
	    RECT 27.8000 166.9000 28.2000 167.8000 ;
	    RECT 34.2000 166.8000 34.6000 167.6000 ;
	    RECT 43.8000 166.9000 44.2000 170.2000 ;
	    RECT 44.6000 168.9000 45.0000 170.2000 ;
	    RECT 46.2000 167.9000 46.6000 170.2000 ;
	    RECT 49.2000 169.2000 49.6000 170.2000 ;
	    RECT 49.2000 168.8000 49.8000 169.2000 ;
	    RECT 49.2000 167.9000 49.6000 168.8000 ;
	    RECT 50.2000 167.9000 50.6000 170.2000 ;
	    RECT 51.8000 168.9000 52.2000 170.2000 ;
	    RECT 53.9000 169.2000 54.3000 170.2000 ;
	    RECT 53.9000 168.8000 54.6000 169.2000 ;
	    RECT 55.0000 168.9000 55.4000 170.2000 ;
	    RECT 56.6000 168.9000 57.0000 170.2000 ;
	    RECT 53.9000 167.9000 54.3000 168.8000 ;
	    RECT 59.8000 168.3000 60.2000 170.2000 ;
	    RECT 62.2000 168.9000 62.6000 170.2000 ;
	    RECT 64.1000 167.9000 64.5000 170.2000 ;
	    RECT 66.2000 168.9000 66.6000 170.2000 ;
	    RECT 67.0000 168.9000 67.4000 170.2000 ;
	    RECT 69.1000 167.9000 69.5000 170.2000 ;
	    RECT 71.0000 168.9000 71.4000 170.2000 ;
	    RECT 71.8000 168.9000 72.2000 170.2000 ;
	    RECT 73.9000 167.9000 74.3000 170.2000 ;
	    RECT 75.8000 168.9000 76.2000 170.2000 ;
	    RECT 77.4000 168.0000 77.8000 170.2000 ;
	    RECT 80.2000 168.9000 80.6000 170.2000 ;
	    RECT 81.8000 168.9000 82.3000 170.2000 ;
	    RECT 84.6000 167.9000 85.0000 170.2000 ;
	    RECT 87.0000 167.9000 87.4000 170.2000 ;
	    RECT 89.7000 168.9000 90.2000 170.2000 ;
	    RECT 91.4000 168.9000 91.8000 170.2000 ;
	    RECT 94.2000 168.0000 94.6000 170.2000 ;
	    RECT 95.8000 168.9000 96.2000 170.2000 ;
	    RECT 97.4000 168.9000 97.8000 170.2000 ;
	    RECT 99.0000 168.9000 99.4000 170.2000 ;
	    RECT 99.8000 167.9000 100.2000 170.2000 ;
	    RECT 102.8000 167.9000 103.2000 170.2000 ;
	    RECT 104.6000 168.9000 105.0000 170.2000 ;
	    RECT 107.8000 167.9000 108.2000 170.2000 ;
	    RECT 110.5000 168.9000 111.0000 170.2000 ;
	    RECT 112.2000 168.9000 112.6000 170.2000 ;
	    RECT 115.0000 168.0000 115.4000 170.2000 ;
	    RECT 116.6000 168.9000 117.0000 170.2000 ;
	    RECT 118.5000 167.9000 118.9000 170.2000 ;
	    RECT 120.6000 168.9000 121.0000 170.2000 ;
	    RECT 122.2000 168.0000 122.6000 170.2000 ;
	    RECT 125.0000 168.9000 125.4000 170.2000 ;
	    RECT 126.6000 168.9000 127.1000 170.2000 ;
	    RECT 129.4000 167.9000 129.8000 170.2000 ;
	    RECT 131.0000 168.9000 131.4000 170.2000 ;
	    RECT 132.6000 168.9000 133.0000 170.2000 ;
	    RECT 134.2000 168.9000 134.6000 170.2000 ;
	    RECT 135.0000 168.9000 135.4000 170.2000 ;
	    RECT 137.1000 167.9000 137.5000 170.2000 ;
	    RECT 139.0000 168.9000 139.4000 170.2000 ;
	    RECT 139.8000 168.9000 140.2000 170.2000 ;
	    RECT 141.4000 168.9000 141.8000 170.2000 ;
	    RECT 143.0000 168.9000 143.4000 170.2000 ;
	    RECT 144.6000 168.0000 145.0000 170.2000 ;
	    RECT 147.4000 168.9000 147.8000 170.2000 ;
	    RECT 149.0000 168.9000 149.5000 170.2000 ;
	    RECT 151.8000 167.9000 152.2000 170.2000 ;
	    RECT 153.4000 168.9000 153.8000 170.2000 ;
	    RECT 155.8000 168.0000 156.2000 170.2000 ;
	    RECT 158.6000 168.9000 159.0000 170.2000 ;
	    RECT 160.2000 168.9000 160.7000 170.2000 ;
	    RECT 163.0000 167.9000 163.4000 170.2000 ;
	    RECT 166.2000 168.9000 166.6000 170.2000 ;
	    RECT 167.8000 168.9000 168.2000 170.2000 ;
	    RECT 168.6000 168.9000 169.0000 170.2000 ;
	    RECT 170.2000 168.9000 170.6000 170.2000 ;
	    RECT 171.8000 168.9000 172.2000 170.2000 ;
	    RECT 173.4000 167.9000 173.8000 170.2000 ;
	    RECT 176.1000 168.9000 176.6000 170.2000 ;
	    RECT 177.8000 168.9000 178.2000 170.2000 ;
	    RECT 180.6000 168.0000 181.0000 170.2000 ;
	    RECT 182.2000 168.9000 182.6000 170.2000 ;
	    RECT 183.8000 168.9000 184.2000 170.2000 ;
	    RECT 185.4000 168.9000 185.8000 170.2000 ;
	    RECT 187.0000 168.0000 187.4000 170.2000 ;
	    RECT 189.8000 168.9000 190.2000 170.2000 ;
	    RECT 191.4000 168.9000 191.9000 170.2000 ;
	    RECT 194.2000 167.9000 194.6000 170.2000 ;
	    RECT 196.6000 167.9000 197.0000 170.2000 ;
	    RECT 199.3000 168.9000 199.8000 170.2000 ;
	    RECT 201.0000 168.9000 201.4000 170.2000 ;
	    RECT 203.8000 168.0000 204.2000 170.2000 ;
	    RECT 205.4000 168.9000 205.8000 170.2000 ;
	    RECT 207.5000 167.9000 207.9000 170.2000 ;
	    RECT 208.6000 168.9000 209.0000 170.2000 ;
	    RECT 210.2000 168.9000 210.6000 170.2000 ;
	    RECT 214.2000 167.9000 214.6000 170.2000 ;
	    RECT 216.6000 168.3000 217.0000 170.2000 ;
	    RECT 218.2000 168.9000 218.6000 170.2000 ;
	    RECT 219.8000 168.9000 220.2000 170.2000 ;
	    RECT 222.2000 167.9000 222.6000 170.2000 ;
	    RECT 223.0000 167.9000 223.4000 170.2000 ;
	    RECT 225.4000 168.9000 225.8000 170.2000 ;
	    RECT 227.0000 168.9000 227.4000 170.2000 ;
	    RECT 228.6000 168.9000 229.0000 170.2000 ;
	    RECT 230.2000 168.3000 230.6000 170.2000 ;
	    RECT 233.4000 168.3000 233.8000 170.2000 ;
	    RECT 236.6000 168.3000 237.0000 170.2000 ;
	    RECT 241.4000 168.3000 241.8000 170.2000 ;
	    RECT 244.1000 168.0000 244.5000 170.2000 ;
	    RECT 247.0000 168.3000 247.4000 170.2000 ;
	    RECT 249.4000 167.9000 249.8000 170.2000 ;
	    RECT 251.0000 167.9000 251.4000 170.2000 ;
	    RECT 253.4000 168.3000 253.8000 170.2000 ;
	    RECT 255.8000 168.9000 256.2000 170.2000 ;
	    RECT 257.9000 167.9000 258.3000 170.2000 ;
	    RECT 259.0000 168.9000 259.4000 170.2000 ;
	    RECT 261.1000 167.9000 261.5000 170.2000 ;
	    RECT 263.0000 168.2000 263.5000 170.2000 ;
	    RECT 266.1000 169.9000 266.5000 170.2000 ;
	    RECT 266.1000 168.2000 266.6000 169.9000 ;
	    RECT 268.6000 167.9000 269.0000 170.2000 ;
	    RECT 270.2000 167.9000 270.6000 170.2000 ;
	    RECT 46.2000 167.1000 46.5000 167.9000 ;
	    RECT 47.0000 167.1000 47.4000 167.2000 ;
	    RECT 46.2000 166.8000 47.4000 167.1000 ;
	    RECT 47.1000 166.6000 47.4000 166.8000 ;
	    RECT 48.6000 167.1000 49.0000 167.2000 ;
	    RECT 49.4000 167.1000 49.8000 167.2000 ;
	    RECT 48.6000 166.8000 49.8000 167.1000 ;
	    RECT 53.4000 167.1000 53.8000 167.2000 ;
	    RECT 54.2000 167.1000 54.6000 167.2000 ;
	    RECT 53.4000 166.8000 54.6000 167.1000 ;
	    RECT 0.6000 165.8000 1.0000 166.6000 ;
	    RECT 47.1000 166.2000 47.5000 166.6000 ;
	    RECT 48.6000 166.4000 49.0000 166.8000 ;
	    RECT 53.4000 166.4000 53.8000 166.8000 ;
	    RECT 59.8000 165.8000 60.2000 166.6000 ;
	    RECT 11.0000 153.4000 11.4000 154.2000 ;
	    RECT 11.8000 153.4000 12.2000 154.2000 ;
	    RECT 32.6000 154.1000 33.0000 154.6000 ;
	    RECT 34.1000 154.4000 34.5000 154.8000 ;
	    RECT 0.6000 152.4000 1.0000 153.2000 ;
	    RECT 0.6000 150.8000 1.0000 152.1000 ;
	    RECT 2.2000 150.8000 2.6000 153.1000 ;
	    RECT 5.2000 150.8000 5.6000 153.1000 ;
	    RECT 7.0000 152.4000 7.4000 153.2000 ;
	    RECT 7.0000 150.8000 7.4000 152.1000 ;
	    RECT 7.8000 150.8000 8.2000 152.1000 ;
	    RECT 11.0000 150.8000 11.4000 153.1000 ;
	    RECT 11.8000 150.8000 12.2000 153.1000 ;
	    RECT 14.2000 150.8000 14.6000 154.1000 ;
	    RECT 31.0000 153.8000 33.0000 154.1000 ;
	    RECT 34.2000 154.2000 34.5000 154.4000 ;
	    RECT 34.2000 154.1000 34.6000 154.2000 ;
	    RECT 36.6000 154.1000 37.0000 154.6000 ;
	    RECT 42.2000 154.4000 42.6000 155.2000 ;
	    RECT 34.2000 153.8000 37.0000 154.1000 ;
	    RECT 17.4000 150.8000 17.8000 152.1000 ;
	    RECT 19.0000 150.8000 19.4000 152.1000 ;
	    RECT 19.8000 150.8000 20.2000 152.1000 ;
	    RECT 21.4000 150.8000 21.8000 152.9000 ;
	    RECT 23.8000 150.8000 24.2000 152.7000 ;
	    RECT 26.2000 150.8000 26.6000 152.1000 ;
	    RECT 27.8000 150.8000 28.2000 152.1000 ;
	    RECT 31.0000 150.8000 31.4000 153.8000 ;
	    RECT 35.0000 153.1000 35.3000 153.8000 ;
	    RECT 32.0000 150.8000 32.4000 153.1000 ;
	    RECT 35.0000 150.8000 35.4000 153.1000 ;
	    RECT 36.1000 150.8000 36.5000 153.1000 ;
	    RECT 38.2000 150.8000 38.6000 152.1000 ;
	    RECT 39.0000 150.8000 39.4000 152.1000 ;
	    RECT 40.6000 150.8000 41.0000 152.1000 ;
	    RECT 42.2000 150.8000 42.6000 152.7000 ;
	    RECT 45.4000 150.8000 45.8000 153.1000 ;
	    RECT 47.0000 150.8000 47.4000 152.1000 ;
	    RECT 48.6000 150.8000 49.0000 152.1000 ;
	    RECT 50.2000 150.8000 50.6000 152.1000 ;
	    RECT 51.8000 150.8000 52.2000 153.0000 ;
	    RECT 54.6000 150.8000 55.0000 152.1000 ;
	    RECT 56.2000 150.8000 56.7000 152.1000 ;
	    RECT 59.0000 150.8000 59.4000 153.1000 ;
	    RECT 63.0000 150.8000 63.4000 153.1000 ;
	    RECT 65.7000 150.8000 66.2000 152.1000 ;
	    RECT 67.4000 150.8000 67.8000 152.1000 ;
	    RECT 70.2000 150.8000 70.6000 153.0000 ;
	    RECT 71.8000 150.8000 72.2000 153.1000 ;
	    RECT 73.4000 150.8000 73.8000 153.1000 ;
	    RECT 75.8000 150.8000 76.2000 153.1000 ;
	    RECT 77.4000 150.8000 77.8000 152.1000 ;
	    RECT 79.0000 150.8000 79.4000 152.1000 ;
	    RECT 80.6000 150.8000 81.0000 152.1000 ;
	    RECT 81.4000 150.8000 81.8000 153.1000 ;
	    RECT 83.0000 150.8000 83.4000 153.1000 ;
	    RECT 86.2000 150.8000 86.6000 152.7000 ;
	    RECT 87.8000 150.8000 88.2000 152.1000 ;
	    RECT 89.4000 150.8000 89.8000 152.1000 ;
	    RECT 91.0000 150.8000 91.4000 152.7000 ;
	    RECT 93.4000 150.8000 93.8000 153.1000 ;
	    RECT 95.8000 150.8000 96.2000 152.1000 ;
	    RECT 97.4000 150.8000 97.8000 152.1000 ;
	    RECT 98.2000 150.8000 98.6000 152.1000 ;
	    RECT 99.8000 150.8000 100.2000 153.1000 ;
	    RECT 102.2000 150.8000 102.6000 152.1000 ;
	    RECT 103.8000 150.8000 104.2000 152.1000 ;
	    RECT 106.2000 150.8000 106.6000 152.7000 ;
	    RECT 109.4000 150.8000 109.8000 153.1000 ;
	    RECT 112.6000 150.8000 113.0000 153.0000 ;
	    RECT 115.4000 150.8000 115.8000 152.1000 ;
	    RECT 117.0000 150.8000 117.5000 152.1000 ;
	    RECT 119.8000 150.8000 120.2000 153.1000 ;
	    RECT 122.2000 150.8000 122.6000 153.1000 ;
	    RECT 124.6000 150.8000 125.0000 153.1000 ;
	    RECT 127.3000 150.8000 127.8000 152.1000 ;
	    RECT 129.0000 150.8000 129.4000 152.1000 ;
	    RECT 131.8000 150.8000 132.2000 153.0000 ;
	    RECT 133.4000 150.8000 133.8000 152.1000 ;
	    RECT 135.0000 150.8000 135.4000 152.9000 ;
	    RECT 136.6000 150.8000 137.0000 152.1000 ;
	    RECT 138.7000 150.8000 139.1000 153.1000 ;
	    RECT 140.6000 150.8000 141.0000 152.1000 ;
	    RECT 142.2000 150.8000 142.6000 153.1000 ;
	    RECT 144.9000 150.8000 145.4000 152.1000 ;
	    RECT 146.6000 150.8000 147.0000 152.1000 ;
	    RECT 149.4000 150.8000 149.8000 153.0000 ;
	    RECT 151.0000 150.8000 151.4000 153.1000 ;
	    RECT 154.0000 150.8000 154.4000 153.1000 ;
	    RECT 155.8000 150.8000 156.2000 153.1000 ;
	    RECT 159.8000 150.8000 160.2000 153.0000 ;
	    RECT 162.6000 150.8000 163.0000 152.1000 ;
	    RECT 164.2000 150.8000 164.7000 152.1000 ;
	    RECT 167.0000 150.8000 167.4000 153.1000 ;
	    RECT 168.6000 150.8000 169.0000 152.1000 ;
	    RECT 170.7000 150.8000 171.1000 153.1000 ;
	    RECT 173.4000 150.8000 173.8000 152.7000 ;
	    RECT 175.0000 150.8000 175.4000 152.1000 ;
	    RECT 176.6000 150.8000 177.0000 152.1000 ;
	    RECT 179.0000 150.8000 179.4000 153.1000 ;
	    RECT 179.8000 150.8000 180.2000 153.1000 ;
	    RECT 182.2000 150.8000 182.6000 152.1000 ;
	    RECT 183.8000 150.8000 184.2000 152.1000 ;
	    RECT 184.6000 150.8000 185.0000 152.1000 ;
	    RECT 186.7000 150.8000 187.1000 153.1000 ;
	    RECT 189.4000 150.8000 189.8000 152.7000 ;
	    RECT 191.0000 150.8000 191.4000 152.1000 ;
	    RECT 192.6000 150.8000 193.0000 152.1000 ;
	    RECT 194.2000 150.8000 194.6000 152.7000 ;
	    RECT 196.9000 150.8000 197.3000 153.1000 ;
	    RECT 199.0000 150.8000 199.4000 152.1000 ;
	    RECT 201.4000 150.8000 201.8000 153.1000 ;
	    RECT 203.0000 150.8000 203.4000 153.1000 ;
	    RECT 205.7000 150.8000 206.2000 152.1000 ;
	    RECT 207.4000 150.8000 207.8000 152.1000 ;
	    RECT 210.2000 150.8000 210.6000 153.0000 ;
	    RECT 214.5000 150.8000 214.9000 153.0000 ;
	    RECT 216.6000 150.8000 217.0000 152.1000 ;
	    RECT 218.2000 150.8000 218.6000 152.1000 ;
	    RECT 219.8000 150.8000 220.2000 152.7000 ;
	    RECT 223.0000 150.8000 223.4000 152.7000 ;
	    RECT 226.2000 150.8000 226.6000 152.1000 ;
	    RECT 227.0000 150.8000 227.4000 152.1000 ;
	    RECT 228.6000 150.8000 229.0000 152.1000 ;
	    RECT 230.2000 150.8000 230.6000 153.1000 ;
	    RECT 231.8000 150.8000 232.2000 153.1000 ;
	    RECT 232.6000 150.8000 233.0000 152.1000 ;
	    RECT 234.2000 150.8000 234.6000 152.1000 ;
	    RECT 235.8000 150.8000 236.3000 152.8000 ;
	    RECT 238.9000 151.1000 239.4000 152.8000 ;
	    RECT 238.9000 150.8000 239.3000 151.1000 ;
	    RECT 240.6000 150.8000 241.0000 152.1000 ;
	    RECT 242.2000 150.8000 242.6000 152.1000 ;
	    RECT 243.0000 150.8000 243.4000 152.1000 ;
	    RECT 244.6000 150.8000 245.0000 152.1000 ;
	    RECT 245.7000 150.8000 246.1000 153.1000 ;
	    RECT 247.8000 150.8000 248.2000 152.1000 ;
	    RECT 248.6000 150.8000 249.0000 152.1000 ;
	    RECT 250.2000 150.8000 250.6000 152.1000 ;
	    RECT 251.0000 150.8000 251.4000 152.1000 ;
	    RECT 253.1000 150.8000 253.5000 153.1000 ;
	    RECT 255.0000 150.8000 255.4000 152.7000 ;
	    RECT 257.4000 150.8000 257.8000 152.1000 ;
	    RECT 259.0000 150.8000 259.4000 152.1000 ;
	    RECT 259.8000 150.8000 260.2000 152.1000 ;
	    RECT 261.4000 150.8000 261.8000 152.1000 ;
	    RECT 263.0000 150.8000 263.4000 152.1000 ;
	    RECT 265.4000 150.8000 265.8000 153.1000 ;
	    RECT 267.0000 150.8000 267.4000 152.9000 ;
	    RECT 268.6000 150.8000 269.0000 152.1000 ;
	    RECT 0.2000 150.2000 271.0000 150.8000 ;
	    RECT 0.6000 148.9000 1.0000 150.2000 ;
	    RECT 2.2000 148.9000 2.6000 150.2000 ;
	    RECT 3.8000 148.3000 4.2000 150.2000 ;
	    RECT 7.0000 148.3000 7.4000 150.2000 ;
	    RECT 11.8000 148.3000 12.2000 150.2000 ;
	    RECT 13.4000 148.9000 13.8000 150.2000 ;
	    RECT 17.4000 146.9000 17.8000 150.2000 ;
	    RECT 19.8000 147.9000 20.2000 150.2000 ;
	    RECT 21.4000 148.3000 21.8000 150.2000 ;
	    RECT 24.1000 147.9000 24.5000 150.2000 ;
	    RECT 26.2000 148.9000 26.6000 150.2000 ;
	    RECT 27.3000 147.9000 27.7000 150.2000 ;
	    RECT 29.4000 148.9000 29.8000 150.2000 ;
	    RECT 31.0000 147.9000 31.4000 150.2000 ;
	    RECT 33.7000 148.9000 34.2000 150.2000 ;
	    RECT 35.4000 148.9000 35.8000 150.2000 ;
	    RECT 38.2000 148.0000 38.6000 150.2000 ;
	    RECT 39.8000 148.9000 40.2000 150.2000 ;
	    RECT 42.2000 148.3000 42.6000 150.2000 ;
	    RECT 46.2000 148.9000 46.6000 150.2000 ;
	    RECT 50.2000 149.1000 50.6000 150.2000 ;
	    RECT 51.8000 148.9000 52.2000 150.2000 ;
	    RECT 55.0000 148.3000 55.4000 150.2000 ;
	    RECT 57.4000 148.9000 57.8000 150.2000 ;
	    RECT 60.6000 148.9000 61.0000 150.2000 ;
	    RECT 61.7000 147.9000 62.1000 150.2000 ;
	    RECT 63.8000 148.9000 64.2000 150.2000 ;
	    RECT 65.4000 147.9000 65.8000 150.2000 ;
	    RECT 68.1000 148.9000 68.6000 150.2000 ;
	    RECT 69.8000 148.9000 70.2000 150.2000 ;
	    RECT 72.6000 148.0000 73.0000 150.2000 ;
	    RECT 75.0000 148.0000 75.4000 150.2000 ;
	    RECT 77.8000 148.9000 78.2000 150.2000 ;
	    RECT 79.4000 148.9000 79.9000 150.2000 ;
	    RECT 82.2000 147.9000 82.6000 150.2000 ;
	    RECT 85.4000 147.9000 85.8000 150.2000 ;
	    RECT 87.0000 147.9000 87.4000 150.2000 ;
	    RECT 89.7000 148.9000 90.2000 150.2000 ;
	    RECT 91.4000 148.9000 91.8000 150.2000 ;
	    RECT 94.2000 148.0000 94.6000 150.2000 ;
	    RECT 95.8000 148.9000 96.2000 150.2000 ;
	    RECT 97.4000 148.9000 97.8000 150.2000 ;
	    RECT 99.8000 148.3000 100.2000 150.2000 ;
	    RECT 102.2000 148.9000 102.6000 150.2000 ;
	    RECT 19.8000 146.8000 20.2000 147.6000 ;
	    RECT 103.0000 146.9000 103.4000 150.2000 ;
	    RECT 107.8000 147.9000 108.2000 150.2000 ;
	    RECT 110.2000 148.9000 110.6000 150.2000 ;
	    RECT 111.8000 148.9000 112.2000 150.2000 ;
	    RECT 112.6000 148.9000 113.0000 150.2000 ;
	    RECT 114.2000 148.9000 114.6000 150.2000 ;
	    RECT 115.0000 147.9000 115.4000 150.2000 ;
	    RECT 117.4000 146.9000 117.8000 150.2000 ;
	    RECT 121.4000 148.9000 121.8000 150.2000 ;
	    RECT 123.0000 148.0000 123.4000 150.2000 ;
	    RECT 125.8000 148.9000 126.2000 150.2000 ;
	    RECT 127.4000 148.9000 127.9000 150.2000 ;
	    RECT 130.2000 147.9000 130.6000 150.2000 ;
	    RECT 131.8000 147.9000 132.2000 150.2000 ;
	    RECT 133.7000 147.9000 134.1000 150.2000 ;
	    RECT 135.8000 148.9000 136.2000 150.2000 ;
	    RECT 136.6000 148.9000 137.0000 150.2000 ;
	    RECT 138.4000 147.9000 138.8000 150.2000 ;
	    RECT 141.4000 147.9000 141.8000 150.2000 ;
	    RECT 142.2000 147.9000 142.6000 150.2000 ;
	    RECT 145.2000 147.9000 145.6000 150.2000 ;
	    RECT 147.0000 148.9000 147.4000 150.2000 ;
	    RECT 148.6000 148.0000 149.0000 150.2000 ;
	    RECT 151.4000 148.9000 151.8000 150.2000 ;
	    RECT 153.0000 148.9000 153.5000 150.2000 ;
	    RECT 155.8000 147.9000 156.2000 150.2000 ;
	    RECT 157.4000 147.9000 157.8000 150.2000 ;
	    RECT 159.0000 147.9000 159.4000 150.2000 ;
	    RECT 163.0000 147.9000 163.4000 150.2000 ;
	    RECT 165.7000 148.9000 166.2000 150.2000 ;
	    RECT 167.4000 148.9000 167.8000 150.2000 ;
	    RECT 170.2000 148.0000 170.6000 150.2000 ;
	    RECT 171.8000 148.9000 172.2000 150.2000 ;
	    RECT 173.4000 148.9000 173.8000 150.2000 ;
	    RECT 175.0000 148.9000 175.4000 150.2000 ;
	    RECT 177.4000 148.3000 177.8000 150.2000 ;
	    RECT 180.1000 148.0000 180.5000 150.2000 ;
	    RECT 182.2000 148.9000 182.6000 150.2000 ;
	    RECT 183.8000 148.9000 184.2000 150.2000 ;
	    RECT 185.4000 148.9000 185.8000 150.2000 ;
	    RECT 186.2000 148.9000 186.6000 150.2000 ;
	    RECT 187.8000 148.9000 188.2000 150.2000 ;
	    RECT 189.4000 148.3000 189.8000 150.2000 ;
	    RECT 191.8000 148.9000 192.2000 150.2000 ;
	    RECT 193.4000 148.9000 193.8000 150.2000 ;
	    RECT 195.0000 148.3000 195.4000 150.2000 ;
	    RECT 198.2000 148.0000 198.6000 150.2000 ;
	    RECT 201.0000 148.9000 201.4000 150.2000 ;
	    RECT 202.6000 148.9000 203.1000 150.2000 ;
	    RECT 205.4000 147.9000 205.8000 150.2000 ;
	    RECT 207.0000 148.9000 207.4000 150.2000 ;
	    RECT 209.1000 147.9000 209.5000 150.2000 ;
	    RECT 211.8000 147.9000 212.2000 150.2000 ;
	    RECT 214.5000 147.9000 214.9000 150.2000 ;
	    RECT 216.6000 148.9000 217.0000 150.2000 ;
	    RECT 217.7000 147.9000 218.1000 150.2000 ;
	    RECT 219.8000 148.9000 220.2000 150.2000 ;
	    RECT 222.2000 148.3000 222.6000 150.2000 ;
	    RECT 223.8000 148.9000 224.2000 150.2000 ;
	    RECT 225.4000 148.9000 225.8000 150.2000 ;
	    RECT 226.2000 148.9000 226.6000 150.2000 ;
	    RECT 227.8000 148.9000 228.2000 150.2000 ;
	    RECT 228.6000 148.9000 229.0000 150.2000 ;
	    RECT 230.2000 148.9000 230.6000 150.2000 ;
	    RECT 231.8000 147.9000 232.2000 150.2000 ;
	    RECT 233.4000 147.9000 233.8000 150.2000 ;
	    RECT 235.0000 147.9000 235.4000 150.2000 ;
	    RECT 236.6000 147.9000 237.0000 150.2000 ;
	    RECT 237.4000 148.9000 237.8000 150.2000 ;
	    RECT 239.0000 148.9000 239.4000 150.2000 ;
	    RECT 239.8000 148.9000 240.2000 150.2000 ;
	    RECT 241.4000 148.9000 241.8000 150.2000 ;
	    RECT 243.0000 148.9000 243.4000 150.2000 ;
	    RECT 243.8000 146.9000 244.2000 150.2000 ;
	    RECT 247.0000 148.9000 247.4000 150.2000 ;
	    RECT 248.6000 148.9000 249.0000 150.2000 ;
	    RECT 251.0000 148.3000 251.4000 150.2000 ;
	    RECT 254.2000 148.3000 254.6000 150.2000 ;
	    RECT 256.9000 148.0000 257.3000 150.2000 ;
	    RECT 259.0000 148.9000 259.4000 150.2000 ;
	    RECT 260.6000 148.9000 261.0000 150.2000 ;
	    RECT 263.0000 148.3000 263.4000 150.2000 ;
	    RECT 264.6000 148.9000 265.0000 150.2000 ;
	    RECT 266.2000 148.9000 266.6000 150.2000 ;
	    RECT 267.0000 147.9000 267.4000 150.2000 ;
	    RECT 270.2000 148.9000 270.6000 150.2000 ;
	    RECT 10.2000 145.8000 10.6000 146.6000 ;
	    RECT 11.8000 145.8000 12.2000 146.6000 ;
	    RECT 5.2000 134.2000 5.6000 134.6000 ;
	    RECT 18.4000 134.2000 18.8000 134.6000 ;
	    RECT 89.4000 134.4000 89.8000 135.2000 ;
	    RECT 147.8000 134.4000 148.2000 135.2000 ;
	    RECT 3.0000 130.8000 3.4000 134.1000 ;
	    RECT 5.3000 133.8000 5.8000 134.2000 ;
	    RECT 8.6000 133.4000 9.0000 134.2000 ;
	    RECT 15.0000 133.4000 15.4000 134.2000 ;
	    RECT 18.2000 133.8000 18.7000 134.2000 ;
	    RECT 4.6000 130.8000 5.0000 132.9000 ;
	    RECT 6.2000 130.8000 6.6000 132.1000 ;
	    RECT 8.6000 130.8000 9.0000 133.1000 ;
	    RECT 11.0000 132.4000 11.4000 133.2000 ;
	    RECT 9.4000 130.8000 9.8000 132.1000 ;
	    RECT 11.0000 130.8000 11.4000 132.1000 ;
	    RECT 12.6000 130.8000 13.0000 133.1000 ;
	    RECT 13.4000 130.8000 13.8000 133.1000 ;
	    RECT 15.0000 130.8000 15.4000 133.1000 ;
	    RECT 17.4000 130.8000 17.8000 132.1000 ;
	    RECT 19.0000 130.8000 19.4000 132.9000 ;
	    RECT 20.6000 130.8000 21.0000 134.1000 ;
	    RECT 23.8000 130.8000 24.2000 132.1000 ;
	    RECT 25.4000 130.8000 25.8000 132.1000 ;
	    RECT 27.3000 130.8000 27.7000 133.0000 ;
	    RECT 29.4000 130.8000 29.8000 133.1000 ;
	    RECT 32.6000 130.8000 33.0000 132.7000 ;
	    RECT 36.6000 130.8000 37.0000 132.7000 ;
	    RECT 39.0000 130.8000 39.4000 132.1000 ;
	    RECT 40.6000 130.8000 41.0000 133.1000 ;
	    RECT 43.3000 130.8000 43.8000 132.1000 ;
	    RECT 45.0000 130.8000 45.4000 132.1000 ;
	    RECT 47.8000 130.8000 48.2000 133.0000 ;
	    RECT 49.4000 130.8000 49.8000 132.1000 ;
	    RECT 51.0000 130.8000 51.4000 132.1000 ;
	    RECT 53.1000 130.8000 53.5000 133.0000 ;
	    RECT 57.4000 130.8000 57.8000 132.7000 ;
	    RECT 60.6000 130.8000 61.0000 132.1000 ;
	    RECT 63.0000 130.8000 63.4000 133.0000 ;
	    RECT 65.8000 130.8000 66.2000 132.1000 ;
	    RECT 67.4000 130.8000 67.9000 132.1000 ;
	    RECT 70.2000 130.8000 70.6000 133.1000 ;
	    RECT 71.8000 130.8000 72.2000 133.1000 ;
	    RECT 73.4000 130.8000 73.8000 133.1000 ;
	    RECT 75.8000 130.8000 76.2000 133.0000 ;
	    RECT 78.6000 130.8000 79.0000 132.1000 ;
	    RECT 80.2000 130.8000 80.7000 132.1000 ;
	    RECT 83.0000 130.8000 83.4000 133.1000 ;
	    RECT 84.6000 130.8000 85.0000 133.1000 ;
	    RECT 86.2000 130.8000 86.6000 133.1000 ;
	    RECT 87.8000 130.8000 88.2000 132.1000 ;
	    RECT 90.2000 130.8000 90.6000 133.1000 ;
	    RECT 91.8000 130.8000 92.2000 133.1000 ;
	    RECT 93.4000 130.8000 93.8000 133.1000 ;
	    RECT 95.0000 130.8000 95.4000 133.1000 ;
	    RECT 96.6000 130.8000 97.0000 133.1000 ;
	    RECT 98.2000 130.8000 98.6000 133.1000 ;
	    RECT 99.0000 130.8000 99.4000 132.1000 ;
	    RECT 100.6000 130.8000 101.0000 133.1000 ;
	    RECT 106.2000 130.8000 106.6000 131.9000 ;
	    RECT 107.8000 130.8000 108.2000 132.1000 ;
	    RECT 111.0000 130.8000 111.4000 132.1000 ;
	    RECT 112.6000 130.8000 113.0000 132.1000 ;
	    RECT 114.7000 130.8000 115.1000 133.0000 ;
	    RECT 116.6000 130.8000 117.0000 132.1000 ;
	    RECT 118.2000 130.8000 118.6000 132.1000 ;
	    RECT 119.8000 130.8000 120.2000 133.0000 ;
	    RECT 122.6000 130.8000 123.0000 132.1000 ;
	    RECT 124.2000 130.8000 124.7000 132.1000 ;
	    RECT 127.0000 130.8000 127.4000 133.1000 ;
	    RECT 129.4000 130.8000 129.8000 133.0000 ;
	    RECT 132.2000 130.8000 132.6000 132.1000 ;
	    RECT 133.8000 130.8000 134.3000 132.1000 ;
	    RECT 136.6000 130.8000 137.0000 133.1000 ;
	    RECT 139.0000 130.8000 139.4000 133.0000 ;
	    RECT 141.8000 130.8000 142.2000 132.1000 ;
	    RECT 143.4000 130.8000 143.9000 132.1000 ;
	    RECT 146.2000 130.8000 146.6000 133.1000 ;
	    RECT 148.6000 130.8000 149.0000 133.1000 ;
	    RECT 151.0000 130.8000 151.4000 133.0000 ;
	    RECT 153.8000 130.8000 154.2000 132.1000 ;
	    RECT 155.4000 130.8000 155.9000 132.1000 ;
	    RECT 158.2000 130.8000 158.6000 133.1000 ;
	    RECT 161.4000 130.8000 161.8000 133.1000 ;
	    RECT 163.0000 130.8000 163.4000 133.1000 ;
	    RECT 164.6000 130.8000 165.0000 133.1000 ;
	    RECT 166.2000 130.8000 166.6000 133.1000 ;
	    RECT 167.8000 130.8000 168.2000 133.1000 ;
	    RECT 168.6000 130.8000 169.0000 133.1000 ;
	    RECT 170.2000 130.8000 170.6000 133.1000 ;
	    RECT 171.8000 130.8000 172.2000 133.1000 ;
	    RECT 173.4000 130.8000 173.8000 133.1000 ;
	    RECT 175.0000 130.8000 175.4000 133.1000 ;
	    RECT 175.8000 130.8000 176.2000 134.1000 ;
	    RECT 179.8000 130.8000 180.2000 133.1000 ;
	    RECT 181.4000 130.8000 181.8000 133.1000 ;
	    RECT 183.0000 130.8000 183.4000 133.1000 ;
	    RECT 184.6000 130.8000 185.0000 133.1000 ;
	    RECT 186.2000 130.8000 186.6000 133.1000 ;
	    RECT 187.8000 130.8000 188.2000 133.1000 ;
	    RECT 189.4000 130.8000 189.8000 133.1000 ;
	    RECT 191.0000 130.8000 191.4000 133.1000 ;
	    RECT 191.8000 130.8000 192.2000 133.1000 ;
	    RECT 193.4000 130.8000 193.8000 133.1000 ;
	    RECT 194.2000 130.8000 194.6000 132.1000 ;
	    RECT 195.8000 130.8000 196.2000 132.1000 ;
	    RECT 196.6000 130.8000 197.0000 134.1000 ;
	    RECT 200.6000 130.8000 201.0000 132.1000 ;
	    RECT 203.0000 130.8000 203.4000 133.1000 ;
	    RECT 203.8000 130.8000 204.2000 132.1000 ;
	    RECT 205.4000 130.8000 205.8000 132.1000 ;
	    RECT 207.0000 130.8000 207.4000 132.1000 ;
	    RECT 209.4000 130.8000 209.8000 132.7000 ;
	    RECT 212.6000 130.8000 213.0000 132.1000 ;
	    RECT 214.7000 130.8000 215.1000 133.1000 ;
	    RECT 215.8000 130.8000 216.2000 133.1000 ;
	    RECT 218.2000 130.8000 218.6000 133.1000 ;
	    RECT 220.6000 130.8000 221.0000 133.1000 ;
	    RECT 223.8000 130.8000 224.2000 132.1000 ;
	    RECT 224.6000 130.8000 225.0000 133.1000 ;
	    RECT 227.0000 130.8000 227.4000 133.1000 ;
	    RECT 229.4000 130.8000 229.8000 133.1000 ;
	    RECT 231.8000 130.8000 232.2000 133.1000 ;
	    RECT 234.2000 130.8000 234.6000 133.1000 ;
	    RECT 236.6000 130.8000 237.0000 132.1000 ;
	    RECT 238.2000 130.8000 238.6000 132.1000 ;
	    RECT 239.0000 130.8000 239.4000 132.1000 ;
	    RECT 240.6000 130.8000 241.0000 132.1000 ;
	    RECT 241.4000 130.8000 241.8000 132.1000 ;
	    RECT 243.0000 130.8000 243.4000 132.1000 ;
	    RECT 245.4000 130.8000 245.8000 132.7000 ;
	    RECT 247.8000 130.8000 248.2000 132.7000 ;
	    RECT 251.0000 130.8000 251.4000 132.7000 ;
	    RECT 255.0000 130.8000 255.4000 132.7000 ;
	    RECT 259.0000 130.8000 259.4000 132.7000 ;
	    RECT 260.6000 130.8000 261.0000 132.1000 ;
	    RECT 262.2000 130.8000 262.6000 132.1000 ;
	    RECT 264.1000 130.8000 264.5000 133.0000 ;
	    RECT 267.0000 130.8000 267.4000 133.1000 ;
	    RECT 268.6000 130.8000 269.0000 133.1000 ;
	    RECT 0.2000 130.2000 271.0000 130.8000 ;
	    RECT 1.5000 129.9000 1.9000 130.2000 ;
	    RECT 1.4000 128.2000 1.9000 129.9000 ;
	    RECT 4.5000 128.2000 5.0000 130.2000 ;
	    RECT 6.5000 127.9000 6.9000 130.2000 ;
	    RECT 8.6000 128.9000 9.0000 130.2000 ;
	    RECT 9.4000 128.9000 9.8000 130.2000 ;
	    RECT 11.0000 128.9000 11.4000 130.2000 ;
	    RECT 12.6000 128.9000 13.0000 130.2000 ;
	    RECT 14.3000 129.9000 14.7000 130.2000 ;
	    RECT 9.4000 127.8000 9.8000 128.6000 ;
	    RECT 14.2000 128.2000 14.7000 129.9000 ;
	    RECT 17.3000 128.2000 17.8000 130.2000 ;
	    RECT 19.0000 128.9000 19.4000 130.2000 ;
	    RECT 20.6000 128.9000 21.0000 130.2000 ;
	    RECT 20.6000 127.8000 21.0000 128.6000 ;
	    RECT 21.7000 127.9000 22.1000 130.2000 ;
	    RECT 23.8000 128.9000 24.2000 130.2000 ;
	    RECT 24.6000 128.9000 25.0000 130.2000 ;
	    RECT 26.2000 128.9000 26.6000 130.2000 ;
	    RECT 27.8000 128.9000 28.2000 130.2000 ;
	    RECT 27.8000 127.8000 28.2000 128.6000 ;
	    RECT 29.4000 128.3000 29.8000 130.2000 ;
	    RECT 31.8000 127.9000 32.2000 130.2000 ;
	    RECT 34.8000 127.9000 35.2000 130.2000 ;
	    RECT 35.8000 128.9000 36.2000 130.2000 ;
	    RECT 39.0000 127.9000 39.4000 130.2000 ;
	    RECT 41.4000 128.3000 41.8000 130.2000 ;
	    RECT 43.8000 128.9000 44.2000 130.2000 ;
	    RECT 45.4000 127.9000 45.8000 130.2000 ;
	    RECT 48.1000 128.9000 48.6000 130.2000 ;
	    RECT 49.8000 128.9000 50.2000 130.2000 ;
	    RECT 52.6000 128.0000 53.0000 130.2000 ;
	    RECT 55.5000 128.0000 55.9000 130.2000 ;
	    RECT 59.8000 128.1000 60.2000 130.2000 ;
	    RECT 61.4000 128.9000 61.8000 130.2000 ;
	    RECT 62.2000 128.9000 62.6000 130.2000 ;
	    RECT 63.8000 128.1000 64.2000 130.2000 ;
	    RECT 66.7000 128.0000 67.1000 130.2000 ;
	    RECT 69.4000 128.0000 69.8000 130.2000 ;
	    RECT 72.2000 128.9000 72.6000 130.2000 ;
	    RECT 73.8000 128.9000 74.3000 130.2000 ;
	    RECT 76.6000 127.9000 77.0000 130.2000 ;
	    RECT 78.2000 128.9000 78.6000 130.2000 ;
	    RECT 80.3000 127.9000 80.7000 130.2000 ;
	    RECT 83.0000 128.3000 83.4000 130.2000 ;
	    RECT 84.6000 127.9000 85.0000 130.2000 ;
	    RECT 86.2000 127.9000 86.6000 130.2000 ;
	    RECT 87.8000 127.9000 88.2000 130.2000 ;
	    RECT 89.4000 127.9000 89.8000 130.2000 ;
	    RECT 91.0000 127.9000 91.4000 130.2000 ;
	    RECT 91.8000 128.9000 92.2000 130.2000 ;
	    RECT 93.4000 128.9000 93.8000 130.2000 ;
	    RECT 94.2000 127.9000 94.6000 130.2000 ;
	    RECT 95.8000 127.9000 96.2000 130.2000 ;
	    RECT 98.7000 128.0000 99.1000 130.2000 ;
	    RECT 100.6000 127.9000 101.0000 130.2000 ;
	    RECT 103.8000 128.3000 104.2000 130.2000 ;
	    RECT 106.2000 128.9000 106.6000 130.2000 ;
	    RECT 107.8000 128.1000 108.2000 130.2000 ;
	    RECT 112.6000 127.9000 113.0000 130.2000 ;
	    RECT 2.2000 127.7000 3.0000 127.8000 ;
	    RECT 2.0000 127.4000 3.0000 127.7000 ;
	    RECT 3.9000 127.4000 4.3000 127.8000 ;
	    RECT 15.0000 127.7000 15.8000 127.8000 ;
	    RECT 2.0000 127.2000 2.3000 127.4000 ;
	    RECT 0.6000 126.9000 2.3000 127.2000 ;
	    RECT 4.0000 127.2000 4.3000 127.4000 ;
	    RECT 14.8000 127.4000 15.8000 127.7000 ;
	    RECT 16.7000 127.4000 17.1000 127.8000 ;
	    RECT 14.8000 127.2000 15.1000 127.4000 ;
	    RECT 0.6000 126.8000 1.4000 126.9000 ;
	    RECT 4.0000 126.8000 4.4000 127.2000 ;
	    RECT 13.4000 126.9000 15.1000 127.2000 ;
	    RECT 16.8000 127.2000 17.1000 127.4000 ;
	    RECT 13.4000 126.8000 14.2000 126.9000 ;
	    RECT 16.8000 126.8000 17.2000 127.2000 ;
	    RECT 113.4000 126.9000 113.8000 130.2000 ;
	    RECT 117.7000 128.0000 118.1000 130.2000 ;
	    RECT 120.6000 128.9000 121.0000 130.2000 ;
	    RECT 121.4000 128.9000 121.8000 130.2000 ;
	    RECT 123.0000 128.9000 123.4000 130.2000 ;
	    RECT 124.6000 128.3000 125.0000 130.2000 ;
	    RECT 127.0000 128.9000 127.4000 130.2000 ;
	    RECT 128.6000 128.9000 129.0000 130.2000 ;
	    RECT 130.2000 127.9000 130.6000 130.2000 ;
	    RECT 132.9000 128.9000 133.4000 130.2000 ;
	    RECT 134.6000 128.9000 135.0000 130.2000 ;
	    RECT 137.4000 128.0000 137.8000 130.2000 ;
	    RECT 139.3000 127.9000 139.7000 130.2000 ;
	    RECT 141.4000 128.9000 141.8000 130.2000 ;
	    RECT 143.8000 128.3000 144.2000 130.2000 ;
	    RECT 145.4000 128.9000 145.8000 130.2000 ;
	    RECT 147.0000 128.9000 147.4000 130.2000 ;
	    RECT 148.1000 129.2000 148.5000 130.2000 ;
	    RECT 147.8000 128.8000 148.5000 129.2000 ;
	    RECT 150.2000 128.9000 150.6000 130.2000 ;
	    RECT 148.1000 127.9000 148.5000 128.8000 ;
	    RECT 151.0000 127.9000 151.4000 130.2000 ;
	    RECT 154.2000 128.9000 154.6000 130.2000 ;
	    RECT 155.8000 128.3000 156.2000 130.2000 ;
	    RECT 158.2000 128.9000 158.6000 130.2000 ;
	    RECT 159.8000 128.9000 160.2000 130.2000 ;
	    RECT 163.0000 127.9000 163.4000 130.2000 ;
	    RECT 164.6000 127.9000 165.0000 130.2000 ;
	    RECT 166.2000 127.9000 166.6000 130.2000 ;
	    RECT 168.9000 128.9000 169.4000 130.2000 ;
	    RECT 170.6000 128.9000 171.0000 130.2000 ;
	    RECT 173.4000 128.0000 173.8000 130.2000 ;
	    RECT 176.6000 127.9000 177.0000 130.2000 ;
	    RECT 177.4000 127.9000 177.8000 130.2000 ;
	    RECT 179.0000 127.9000 179.4000 130.2000 ;
	    RECT 182.2000 127.9000 182.6000 130.2000 ;
	    RECT 183.0000 127.9000 183.4000 130.2000 ;
	    RECT 184.6000 127.9000 185.0000 130.2000 ;
	    RECT 187.8000 127.9000 188.2000 130.2000 ;
	    RECT 188.6000 127.9000 189.0000 130.2000 ;
	    RECT 191.8000 127.9000 192.2000 130.2000 ;
	    RECT 195.0000 126.9000 195.4000 130.2000 ;
	    RECT 196.6000 128.0000 197.0000 130.2000 ;
	    RECT 199.4000 128.9000 199.8000 130.2000 ;
	    RECT 201.0000 128.9000 201.5000 130.2000 ;
	    RECT 203.8000 127.9000 204.2000 130.2000 ;
	    RECT 205.4000 128.9000 205.8000 130.2000 ;
	    RECT 207.0000 128.9000 207.4000 130.2000 ;
	    RECT 207.8000 127.9000 208.2000 130.2000 ;
	    RECT 209.4000 127.9000 209.8000 130.2000 ;
	    RECT 212.6000 128.9000 213.0000 130.2000 ;
	    RECT 214.2000 128.9000 214.6000 130.2000 ;
	    RECT 215.0000 128.9000 215.4000 130.2000 ;
	    RECT 216.6000 128.9000 217.0000 130.2000 ;
	    RECT 217.4000 128.9000 217.8000 130.2000 ;
	    RECT 219.5000 127.9000 219.9000 130.2000 ;
	    RECT 220.6000 128.9000 221.0000 130.2000 ;
	    RECT 222.2000 128.9000 222.6000 130.2000 ;
	    RECT 223.0000 128.9000 223.4000 130.2000 ;
	    RECT 224.6000 128.9000 225.0000 130.2000 ;
	    RECT 225.4000 127.9000 225.8000 130.2000 ;
	    RECT 227.8000 127.9000 228.2000 130.2000 ;
	    RECT 229.4000 127.9000 229.8000 130.2000 ;
	    RECT 231.0000 127.9000 231.4000 130.2000 ;
	    RECT 232.6000 127.9000 233.0000 130.2000 ;
	    RECT 233.4000 128.9000 233.8000 130.2000 ;
	    RECT 235.0000 128.9000 235.4000 130.2000 ;
	    RECT 235.8000 128.9000 236.2000 130.2000 ;
	    RECT 237.4000 128.9000 237.8000 130.2000 ;
	    RECT 238.2000 128.9000 238.6000 130.2000 ;
	    RECT 240.6000 128.3000 241.0000 130.2000 ;
	    RECT 243.0000 128.9000 243.4000 130.2000 ;
	    RECT 244.6000 128.9000 245.0000 130.2000 ;
	    RECT 246.2000 128.9000 246.6000 130.2000 ;
	    RECT 247.8000 128.9000 248.2000 130.2000 ;
	    RECT 248.6000 128.9000 249.0000 130.2000 ;
	    RECT 250.2000 128.9000 250.6000 130.2000 ;
	    RECT 251.8000 128.3000 252.2000 130.2000 ;
	    RECT 255.0000 128.9000 255.4000 130.2000 ;
	    RECT 255.8000 128.9000 256.2000 130.2000 ;
	    RECT 257.9000 127.9000 258.3000 130.2000 ;
	    RECT 259.0000 128.9000 259.4000 130.2000 ;
	    RECT 260.9000 127.9000 261.3000 130.2000 ;
	    RECT 263.0000 128.9000 263.4000 130.2000 ;
	    RECT 263.8000 128.9000 264.2000 130.2000 ;
	    RECT 265.9000 127.9000 266.3000 130.2000 ;
	    RECT 268.6000 127.9000 269.0000 130.2000 ;
	    RECT 123.0000 114.4000 123.4000 115.2000 ;
	    RECT 13.2000 113.8000 13.6000 114.2000 ;
	    RECT 16.2000 114.1000 17.0000 114.2000 ;
	    RECT 13.3000 113.6000 13.6000 113.8000 ;
	    RECT 15.3000 113.8000 17.0000 114.1000 ;
	    RECT 15.3000 113.6000 15.6000 113.8000 ;
	    RECT 13.3000 113.2000 13.7000 113.6000 ;
	    RECT 14.6000 113.3000 15.6000 113.6000 ;
	    RECT 14.6000 113.2000 15.4000 113.3000 ;
	    RECT 3.8000 112.4000 4.2000 113.2000 ;
	    RECT 0.6000 110.8000 1.0000 112.1000 ;
	    RECT 2.2000 110.8000 2.6000 112.1000 ;
	    RECT 3.8000 110.8000 4.2000 112.1000 ;
	    RECT 4.9000 111.2000 5.3000 113.1000 ;
	    RECT 7.8000 112.4000 8.2000 113.2000 ;
	    RECT 4.6000 110.8000 5.3000 111.2000 ;
	    RECT 7.0000 110.8000 7.4000 112.1000 ;
	    RECT 7.8000 110.8000 8.2000 112.1000 ;
	    RECT 9.4000 110.8000 9.8000 112.1000 ;
	    RECT 11.0000 110.8000 11.4000 112.1000 ;
	    RECT 12.6000 110.8000 13.1000 112.8000 ;
	    RECT 15.7000 111.1000 16.2000 112.8000 ;
	    RECT 15.7000 110.8000 16.1000 111.1000 ;
	    RECT 18.2000 110.8000 18.6000 112.7000 ;
	    RECT 20.6000 110.8000 21.0000 113.1000 ;
	    RECT 24.3000 110.8000 24.7000 113.0000 ;
	    RECT 27.0000 110.8000 27.4000 112.7000 ;
	    RECT 30.2000 110.8000 30.6000 112.7000 ;
	    RECT 32.6000 110.8000 33.0000 113.1000 ;
	    RECT 35.6000 110.8000 36.0000 113.1000 ;
	    RECT 37.4000 110.8000 37.8000 113.1000 ;
	    RECT 40.1000 110.8000 40.6000 112.1000 ;
	    RECT 41.8000 110.8000 42.2000 112.1000 ;
	    RECT 44.6000 110.8000 45.0000 113.0000 ;
	    RECT 46.2000 110.8000 46.6000 113.1000 ;
	    RECT 49.4000 110.8000 49.8000 112.1000 ;
	    RECT 51.0000 110.8000 51.4000 113.1000 ;
	    RECT 53.7000 110.8000 54.2000 112.1000 ;
	    RECT 55.4000 110.8000 55.8000 112.1000 ;
	    RECT 58.2000 110.8000 58.6000 113.0000 ;
	    RECT 62.2000 110.8000 62.6000 112.9000 ;
	    RECT 63.8000 110.8000 64.2000 112.1000 ;
	    RECT 65.4000 110.8000 65.8000 113.1000 ;
	    RECT 68.1000 110.8000 68.6000 112.1000 ;
	    RECT 69.8000 110.8000 70.2000 112.1000 ;
	    RECT 72.6000 110.8000 73.0000 113.0000 ;
	    RECT 74.2000 110.8000 74.6000 114.1000 ;
	    RECT 78.2000 110.8000 78.6000 113.0000 ;
	    RECT 81.0000 110.8000 81.4000 112.1000 ;
	    RECT 82.6000 110.8000 83.1000 112.1000 ;
	    RECT 85.4000 110.8000 85.8000 113.1000 ;
	    RECT 87.0000 110.8000 87.4000 112.1000 ;
	    RECT 88.6000 110.8000 89.0000 112.1000 ;
	    RECT 90.2000 110.8000 90.6000 113.1000 ;
	    RECT 92.9000 110.8000 93.4000 112.1000 ;
	    RECT 94.6000 110.8000 95.0000 112.1000 ;
	    RECT 97.4000 110.8000 97.8000 113.0000 ;
	    RECT 99.8000 110.8000 100.2000 112.1000 ;
	    RECT 100.6000 110.8000 101.0000 112.1000 ;
	    RECT 102.2000 110.8000 102.6000 113.1000 ;
	    RECT 105.2000 110.8000 105.6000 113.1000 ;
	    RECT 106.2000 110.8000 106.6000 112.1000 ;
	    RECT 107.8000 110.8000 108.2000 112.1000 ;
	    RECT 111.0000 110.8000 111.4000 112.1000 ;
	    RECT 112.6000 110.8000 113.0000 112.1000 ;
	    RECT 113.4000 110.8000 113.8000 113.1000 ;
	    RECT 116.6000 110.8000 117.0000 112.1000 ;
	    RECT 117.4000 110.8000 117.8000 113.1000 ;
	    RECT 120.6000 110.8000 121.0000 112.1000 ;
	    RECT 122.2000 110.8000 122.6000 113.1000 ;
	    RECT 123.8000 110.8000 124.2000 112.1000 ;
	    RECT 125.4000 110.8000 125.8000 112.1000 ;
	    RECT 126.2000 110.8000 126.6000 112.1000 ;
	    RECT 127.8000 110.8000 128.2000 114.1000 ;
	    RECT 131.8000 110.8000 132.2000 112.1000 ;
	    RECT 134.2000 110.8000 134.6000 112.7000 ;
	    RECT 136.1000 110.8000 136.5000 113.1000 ;
	    RECT 138.2000 110.8000 138.6000 112.1000 ;
	    RECT 140.6000 110.8000 141.0000 112.7000 ;
	    RECT 142.2000 110.8000 142.6000 112.1000 ;
	    RECT 144.3000 110.8000 144.7000 113.1000 ;
	    RECT 146.2000 110.8000 146.6000 112.1000 ;
	    RECT 147.0000 110.8000 147.4000 112.1000 ;
	    RECT 149.1000 110.8000 149.5000 113.1000 ;
	    RECT 150.2000 110.8000 150.6000 113.1000 ;
	    RECT 153.4000 110.8000 153.8000 112.7000 ;
	    RECT 155.8000 110.8000 156.2000 113.1000 ;
	    RECT 157.4000 110.8000 157.8000 113.1000 ;
	    RECT 161.4000 110.8000 161.8000 113.1000 ;
	    RECT 164.1000 110.8000 164.6000 112.1000 ;
	    RECT 165.8000 110.8000 166.2000 112.1000 ;
	    RECT 168.6000 110.8000 169.0000 113.0000 ;
	    RECT 170.2000 110.8000 170.6000 113.1000 ;
	    RECT 172.6000 110.8000 173.0000 112.1000 ;
	    RECT 174.2000 110.8000 174.6000 111.9000 ;
	    RECT 179.3000 110.8000 179.7000 113.0000 ;
	    RECT 182.2000 110.8000 182.6000 113.1000 ;
	    RECT 184.9000 110.8000 185.4000 112.1000 ;
	    RECT 186.6000 110.8000 187.0000 112.1000 ;
	    RECT 189.4000 110.8000 189.8000 113.0000 ;
	    RECT 191.8000 110.8000 192.2000 113.1000 ;
	    RECT 194.5000 110.8000 195.0000 112.1000 ;
	    RECT 196.2000 110.8000 196.6000 112.1000 ;
	    RECT 199.0000 110.8000 199.4000 113.0000 ;
	    RECT 200.6000 110.8000 201.0000 113.1000 ;
	    RECT 202.2000 110.8000 202.6000 113.1000 ;
	    RECT 203.8000 110.8000 204.2000 113.1000 ;
	    RECT 204.6000 110.8000 205.0000 112.1000 ;
	    RECT 206.2000 110.8000 206.6000 112.1000 ;
	    RECT 208.6000 110.8000 209.0000 113.1000 ;
	    RECT 209.4000 110.8000 209.8000 112.1000 ;
	    RECT 213.4000 110.8000 213.8000 112.7000 ;
	    RECT 215.8000 110.8000 216.2000 112.1000 ;
	    RECT 217.4000 110.8000 217.8000 112.1000 ;
	    RECT 219.0000 110.8000 219.4000 112.1000 ;
	    RECT 219.8000 110.8000 220.2000 112.1000 ;
	    RECT 221.4000 110.8000 221.8000 112.1000 ;
	    RECT 223.8000 110.8000 224.2000 112.7000 ;
	    RECT 226.7000 110.8000 227.1000 113.0000 ;
	    RECT 228.6000 110.8000 229.0000 113.1000 ;
	    RECT 231.0000 110.8000 231.4000 112.1000 ;
	    RECT 232.6000 110.8000 233.0000 112.1000 ;
	    RECT 233.4000 110.8000 233.8000 112.1000 ;
	    RECT 235.0000 110.8000 235.4000 112.1000 ;
	    RECT 235.8000 110.8000 236.2000 113.1000 ;
	    RECT 239.5000 110.8000 239.9000 113.0000 ;
	    RECT 241.4000 110.8000 241.8000 113.1000 ;
	    RECT 245.4000 110.8000 245.8000 113.1000 ;
	    RECT 246.2000 110.8000 246.6000 113.1000 ;
	    RECT 250.2000 110.8000 250.6000 113.1000 ;
	    RECT 251.0000 110.8000 251.4000 112.1000 ;
	    RECT 252.6000 110.8000 253.0000 112.1000 ;
	    RECT 253.4000 110.8000 253.8000 112.1000 ;
	    RECT 255.0000 110.8000 255.4000 112.1000 ;
	    RECT 255.8000 110.8000 256.2000 112.1000 ;
	    RECT 257.4000 110.8000 257.8000 112.1000 ;
	    RECT 258.2000 110.8000 258.6000 112.1000 ;
	    RECT 259.8000 110.8000 260.2000 112.1000 ;
	    RECT 261.4000 110.8000 261.8000 112.7000 ;
	    RECT 264.6000 110.8000 265.0000 112.7000 ;
	    RECT 268.6000 110.8000 269.0000 113.1000 ;
	    RECT 0.2000 110.2000 271.0000 110.8000 ;
	    RECT 1.4000 108.3000 1.8000 110.2000 ;
	    RECT 3.8000 107.9000 4.2000 110.2000 ;
	    RECT 6.2000 108.9000 6.6000 110.2000 ;
	    RECT 7.8000 108.9000 8.2000 110.2000 ;
	    RECT 8.9000 107.9000 9.3000 110.2000 ;
	    RECT 11.0000 108.9000 11.4000 110.2000 ;
	    RECT 11.8000 107.9000 12.2000 110.2000 ;
	    RECT 15.0000 108.2000 15.5000 110.2000 ;
	    RECT 18.1000 109.9000 18.5000 110.2000 ;
	    RECT 18.1000 108.2000 18.6000 109.9000 ;
	    RECT 19.8000 108.9000 20.2000 110.2000 ;
	    RECT 21.4000 108.9000 21.8000 110.2000 ;
	    RECT 23.0000 108.9000 23.4000 110.2000 ;
	    RECT 21.4000 107.8000 21.8000 108.6000 ;
	    RECT 24.6000 108.0000 25.0000 110.2000 ;
	    RECT 27.4000 108.9000 27.8000 110.2000 ;
	    RECT 29.0000 108.9000 29.5000 110.2000 ;
	    RECT 31.8000 107.9000 32.2000 110.2000 ;
	    RECT 33.4000 108.9000 33.8000 110.2000 ;
	    RECT 35.0000 108.9000 35.4000 110.2000 ;
	    RECT 36.6000 108.9000 37.0000 110.2000 ;
	    RECT 40.6000 109.1000 41.0000 110.2000 ;
	    RECT 42.2000 108.9000 42.6000 110.2000 ;
	    RECT 44.6000 108.9000 45.0000 110.2000 ;
	    RECT 45.4000 108.9000 45.8000 110.2000 ;
	    RECT 47.0000 108.9000 47.4000 110.2000 ;
	    RECT 48.6000 108.3000 49.0000 110.2000 ;
	    RECT 51.0000 108.9000 51.4000 110.2000 ;
	    RECT 52.6000 108.9000 53.0000 110.2000 ;
	    RECT 55.0000 108.3000 55.4000 110.2000 ;
	    RECT 58.2000 108.9000 58.6000 110.2000 ;
	    RECT 60.3000 107.9000 60.7000 110.2000 ;
	    RECT 61.7000 107.9000 62.1000 110.2000 ;
	    RECT 63.8000 108.9000 64.2000 110.2000 ;
	    RECT 13.4000 107.1000 13.8000 107.2000 ;
	    RECT 14.2000 107.1000 15.0000 107.2000 ;
	    RECT 13.4000 106.8000 15.0000 107.1000 ;
	    RECT 67.0000 106.9000 67.4000 110.2000 ;
	    RECT 68.6000 108.0000 69.0000 110.2000 ;
	    RECT 71.4000 108.9000 71.8000 110.2000 ;
	    RECT 73.0000 108.9000 73.5000 110.2000 ;
	    RECT 75.8000 107.9000 76.2000 110.2000 ;
	    RECT 77.4000 108.9000 77.8000 110.2000 ;
	    RECT 79.5000 107.9000 79.9000 110.2000 ;
	    RECT 82.2000 108.3000 82.6000 110.2000 ;
	    RECT 83.8000 108.9000 84.2000 110.2000 ;
	    RECT 85.9000 107.9000 86.3000 110.2000 ;
	    RECT 88.6000 108.3000 89.0000 110.2000 ;
	    RECT 90.2000 107.9000 90.6000 110.2000 ;
	    RECT 93.4000 108.9000 93.8000 110.2000 ;
	    RECT 96.6000 106.9000 97.0000 110.2000 ;
	    RECT 97.4000 108.9000 97.8000 110.2000 ;
	    RECT 99.0000 108.9000 99.4000 110.2000 ;
	    RECT 99.8000 108.9000 100.2000 110.2000 ;
	    RECT 101.4000 108.1000 101.8000 110.2000 ;
	    RECT 103.8000 108.3000 104.2000 110.2000 ;
	    RECT 108.6000 106.9000 109.0000 110.2000 ;
	    RECT 111.0000 107.9000 111.4000 110.2000 ;
	    RECT 114.0000 107.9000 114.4000 110.2000 ;
	    RECT 115.3000 107.9000 115.7000 110.2000 ;
	    RECT 117.4000 108.9000 117.8000 110.2000 ;
	    RECT 118.2000 108.9000 118.6000 110.2000 ;
	    RECT 119.8000 108.9000 120.2000 110.2000 ;
	    RECT 122.2000 108.3000 122.6000 110.2000 ;
	    RECT 124.6000 108.0000 125.0000 110.2000 ;
	    RECT 127.4000 108.9000 127.8000 110.2000 ;
	    RECT 129.0000 108.9000 129.5000 110.2000 ;
	    RECT 131.8000 107.9000 132.2000 110.2000 ;
	    RECT 134.2000 108.0000 134.6000 110.2000 ;
	    RECT 137.0000 108.9000 137.4000 110.2000 ;
	    RECT 138.6000 108.9000 139.1000 110.2000 ;
	    RECT 141.4000 107.9000 141.8000 110.2000 ;
	    RECT 143.0000 108.9000 143.4000 110.2000 ;
	    RECT 144.6000 108.9000 145.0000 110.2000 ;
	    RECT 148.6000 109.1000 149.0000 110.2000 ;
	    RECT 150.2000 108.9000 150.6000 110.2000 ;
	    RECT 152.9000 108.0000 153.3000 110.2000 ;
	    RECT 155.0000 108.9000 155.4000 110.2000 ;
	    RECT 156.6000 108.1000 157.0000 110.2000 ;
	    RECT 158.5000 107.9000 158.9000 110.2000 ;
	    RECT 160.6000 108.9000 161.0000 110.2000 ;
	    RECT 163.8000 108.9000 164.2000 110.2000 ;
	    RECT 167.0000 106.9000 167.4000 110.2000 ;
	    RECT 169.1000 108.0000 169.5000 110.2000 ;
	    RECT 171.0000 106.9000 171.4000 110.2000 ;
	    RECT 174.2000 107.9000 174.6000 110.2000 ;
	    RECT 178.2000 106.9000 178.6000 110.2000 ;
	    RECT 179.0000 108.9000 179.4000 110.2000 ;
	    RECT 181.1000 107.9000 181.5000 110.2000 ;
	    RECT 183.0000 108.3000 183.4000 110.2000 ;
	    RECT 186.2000 108.2000 186.7000 110.2000 ;
	    RECT 189.3000 109.9000 189.7000 110.2000 ;
	    RECT 189.3000 108.2000 189.8000 109.9000 ;
	    RECT 191.0000 108.9000 191.4000 110.2000 ;
	    RECT 193.1000 107.9000 193.5000 110.2000 ;
	    RECT 195.0000 108.3000 195.4000 110.2000 ;
	    RECT 198.2000 108.2000 198.7000 110.2000 ;
	    RECT 201.3000 109.9000 201.7000 110.2000 ;
	    RECT 201.3000 108.2000 201.8000 109.9000 ;
	    RECT 203.0000 107.9000 203.4000 110.2000 ;
	    RECT 206.2000 108.3000 206.6000 110.2000 ;
	    RECT 208.6000 108.9000 209.0000 110.2000 ;
	    RECT 210.7000 107.9000 211.1000 110.2000 ;
	    RECT 215.0000 108.3000 215.4000 110.2000 ;
	    RECT 217.4000 107.7000 217.8000 110.2000 ;
	    RECT 220.0000 107.5000 220.4000 110.2000 ;
	    RECT 222.2000 108.9000 222.6000 110.2000 ;
	    RECT 224.6000 108.3000 225.0000 110.2000 ;
	    RECT 227.5000 108.0000 227.9000 110.2000 ;
	    RECT 229.4000 107.9000 229.8000 110.2000 ;
	    RECT 231.0000 107.9000 231.4000 110.2000 ;
	    RECT 232.6000 108.9000 233.0000 110.2000 ;
	    RECT 234.2000 108.9000 234.6000 110.2000 ;
	    RECT 235.0000 108.9000 235.4000 110.2000 ;
	    RECT 236.6000 108.9000 237.0000 110.2000 ;
	    RECT 237.4000 108.9000 237.8000 110.2000 ;
	    RECT 239.0000 108.9000 239.4000 110.2000 ;
	    RECT 239.8000 108.9000 240.2000 110.2000 ;
	    RECT 242.3000 109.9000 242.7000 110.2000 ;
	    RECT 242.2000 108.2000 242.7000 109.9000 ;
	    RECT 245.3000 108.2000 245.8000 110.2000 ;
	    RECT 247.0000 108.9000 247.4000 110.2000 ;
	    RECT 248.6000 108.9000 249.0000 110.2000 ;
	    RECT 249.4000 108.9000 249.8000 110.2000 ;
	    RECT 251.5000 107.9000 251.9000 110.2000 ;
	    RECT 253.4000 108.3000 253.8000 110.2000 ;
	    RECT 256.7000 109.9000 257.1000 110.2000 ;
	    RECT 256.6000 108.2000 257.1000 109.9000 ;
	    RECT 259.7000 108.2000 260.2000 110.2000 ;
	    RECT 263.0000 108.3000 263.4000 110.2000 ;
	    RECT 266.2000 108.3000 266.6000 110.2000 ;
	    RECT 268.6000 108.9000 269.0000 110.2000 ;
	    RECT 3.0000 94.4000 3.4000 95.2000 ;
	    RECT 4.6000 94.4000 5.0000 95.2000 ;
	    RECT 8.7000 94.4000 9.1000 94.8000 ;
	    RECT 8.7000 94.2000 9.0000 94.4000 ;
	    RECT 8.6000 94.1000 9.0000 94.2000 ;
	    RECT 7.8000 93.8000 9.0000 94.1000 ;
	    RECT 10.2000 93.8000 10.6000 94.6000 ;
	    RECT 17.4000 93.8000 18.2000 94.2000 ;
	    RECT 7.8000 93.1000 8.1000 93.8000 ;
	    RECT 0.6000 90.8000 1.0000 92.1000 ;
	    RECT 3.0000 90.8000 3.4000 92.7000 ;
	    RECT 6.2000 90.8000 6.6000 92.1000 ;
	    RECT 7.8000 90.8000 8.2000 93.1000 ;
	    RECT 10.8000 90.8000 11.2000 93.1000 ;
	    RECT 13.4000 90.8000 13.8000 93.1000 ;
	    RECT 15.5000 90.8000 15.9000 93.0000 ;
	    RECT 18.2000 90.8000 18.7000 92.8000 ;
	    RECT 21.3000 91.1000 21.8000 92.8000 ;
	    RECT 21.3000 90.8000 21.7000 91.1000 ;
	    RECT 23.8000 90.8000 24.2000 92.7000 ;
	    RECT 27.8000 90.8000 28.2000 93.1000 ;
	    RECT 28.9000 91.2000 29.3000 93.1000 ;
	    RECT 31.8000 92.4000 32.2000 93.2000 ;
	    RECT 28.6000 90.8000 29.3000 91.2000 ;
	    RECT 31.0000 90.8000 31.4000 92.1000 ;
	    RECT 31.8000 90.8000 32.2000 92.1000 ;
	    RECT 33.4000 90.8000 33.8000 92.1000 ;
	    RECT 35.0000 90.8000 35.4000 92.1000 ;
	    RECT 35.8000 90.8000 36.2000 92.1000 ;
	    RECT 38.2000 90.8000 38.7000 92.8000 ;
	    RECT 41.3000 91.1000 41.8000 92.8000 ;
	    RECT 41.3000 90.8000 41.7000 91.1000 ;
	    RECT 43.0000 90.8000 43.4000 92.1000 ;
	    RECT 44.6000 90.8000 45.0000 92.1000 ;
	    RECT 46.2000 90.8000 46.6000 92.1000 ;
	    RECT 47.0000 90.8000 47.4000 92.1000 ;
	    RECT 49.1000 90.8000 49.5000 93.1000 ;
	    RECT 50.2000 90.8000 50.6000 92.1000 ;
	    RECT 51.8000 90.8000 52.2000 92.1000 ;
	    RECT 54.2000 90.8000 54.6000 92.7000 ;
	    RECT 55.8000 90.8000 56.2000 92.1000 ;
	    RECT 59.0000 90.8000 59.4000 92.1000 ;
	    RECT 61.1000 90.8000 61.5000 93.1000 ;
	    RECT 63.0000 90.8000 63.4000 93.1000 ;
	    RECT 65.7000 90.8000 66.2000 92.1000 ;
	    RECT 67.4000 90.8000 67.8000 92.1000 ;
	    RECT 70.2000 90.8000 70.6000 93.0000 ;
	    RECT 71.8000 90.8000 72.2000 94.1000 ;
	    RECT 75.0000 90.8000 75.4000 92.1000 ;
	    RECT 76.6000 90.8000 77.0000 92.1000 ;
	    RECT 79.0000 90.8000 79.4000 93.1000 ;
	    RECT 82.2000 90.8000 82.6000 94.1000 ;
	    RECT 85.4000 90.8000 85.8000 94.1000 ;
	    RECT 86.2000 90.8000 86.6000 93.1000 ;
	    RECT 87.8000 90.8000 88.2000 93.1000 ;
	    RECT 89.4000 90.8000 89.8000 93.1000 ;
	    RECT 91.0000 90.8000 91.4000 93.1000 ;
	    RECT 92.6000 90.8000 93.0000 93.1000 ;
	    RECT 94.2000 90.8000 94.6000 93.1000 ;
	    RECT 97.4000 90.8000 97.8000 92.7000 ;
	    RECT 99.0000 90.8000 99.4000 92.1000 ;
	    RECT 101.1000 90.8000 101.5000 93.1000 ;
	    RECT 103.0000 90.8000 103.4000 92.1000 ;
	    RECT 104.6000 90.8000 105.0000 93.1000 ;
	    RECT 107.3000 90.8000 107.8000 92.1000 ;
	    RECT 109.0000 90.8000 109.4000 92.1000 ;
	    RECT 111.8000 90.8000 112.2000 93.0000 ;
	    RECT 115.8000 90.8000 116.2000 93.1000 ;
	    RECT 118.5000 90.8000 119.0000 92.1000 ;
	    RECT 120.2000 90.8000 120.6000 92.1000 ;
	    RECT 123.0000 90.8000 123.4000 93.0000 ;
	    RECT 125.4000 90.8000 125.8000 93.1000 ;
	    RECT 126.2000 90.8000 126.6000 92.1000 ;
	    RECT 128.6000 90.8000 129.0000 93.0000 ;
	    RECT 131.4000 90.8000 131.8000 92.1000 ;
	    RECT 133.0000 90.8000 133.5000 92.1000 ;
	    RECT 135.8000 90.8000 136.2000 93.1000 ;
	    RECT 137.7000 90.8000 138.1000 93.1000 ;
	    RECT 139.8000 90.8000 140.2000 92.1000 ;
	    RECT 142.2000 90.8000 142.6000 92.7000 ;
	    RECT 144.6000 90.8000 145.0000 92.7000 ;
	    RECT 147.0000 90.8000 147.4000 93.1000 ;
	    RECT 148.6000 90.8000 149.0000 93.1000 ;
	    RECT 150.2000 90.8000 150.6000 93.1000 ;
	    RECT 151.8000 90.8000 152.2000 93.1000 ;
	    RECT 153.4000 90.8000 153.8000 93.1000 ;
	    RECT 155.0000 90.8000 155.4000 93.1000 ;
	    RECT 157.7000 90.8000 158.2000 92.1000 ;
	    RECT 159.4000 90.8000 159.8000 92.1000 ;
	    RECT 162.2000 90.8000 162.6000 93.0000 ;
	    RECT 165.4000 90.8000 165.8000 92.1000 ;
	    RECT 167.5000 90.8000 167.9000 93.1000 ;
	    RECT 170.2000 90.8000 170.6000 93.1000 ;
	    RECT 171.3000 90.8000 171.7000 93.1000 ;
	    RECT 173.4000 90.8000 173.8000 92.1000 ;
	    RECT 175.0000 90.8000 175.4000 93.1000 ;
	    RECT 177.7000 90.8000 178.2000 92.1000 ;
	    RECT 179.4000 90.8000 179.8000 92.1000 ;
	    RECT 182.2000 90.8000 182.6000 93.0000 ;
	    RECT 183.8000 90.8000 184.2000 93.1000 ;
	    RECT 187.0000 90.8000 187.4000 92.7000 ;
	    RECT 190.2000 90.8000 190.6000 92.1000 ;
	    RECT 191.8000 90.8000 192.2000 93.1000 ;
	    RECT 194.5000 90.8000 195.0000 92.1000 ;
	    RECT 196.2000 90.8000 196.6000 92.1000 ;
	    RECT 199.0000 90.8000 199.4000 93.0000 ;
	    RECT 200.6000 90.8000 201.0000 92.1000 ;
	    RECT 202.7000 90.8000 203.1000 93.1000 ;
	    RECT 205.4000 90.8000 205.8000 92.7000 ;
	    RECT 207.0000 90.8000 207.4000 93.1000 ;
	    RECT 209.4000 90.8000 209.8000 92.1000 ;
	    RECT 211.0000 90.8000 211.4000 92.1000 ;
	    RECT 215.0000 90.8000 215.4000 93.1000 ;
	    RECT 216.6000 91.1000 217.1000 92.8000 ;
	    RECT 216.7000 90.8000 217.1000 91.1000 ;
	    RECT 219.7000 90.8000 220.2000 92.8000 ;
	    RECT 221.4000 90.8000 221.8000 92.1000 ;
	    RECT 223.0000 90.8000 223.4000 92.1000 ;
	    RECT 224.6000 90.8000 225.0000 93.1000 ;
	    RECT 226.2000 90.8000 226.6000 93.1000 ;
	    RECT 227.8000 90.8000 228.2000 92.1000 ;
	    RECT 230.2000 90.8000 230.6000 93.1000 ;
	    RECT 232.6000 90.8000 233.0000 93.1000 ;
	    RECT 234.2000 90.8000 234.6000 93.1000 ;
	    RECT 235.8000 90.8000 236.2000 93.1000 ;
	    RECT 237.4000 90.8000 237.8000 92.9000 ;
	    RECT 239.0000 90.8000 239.4000 92.1000 ;
	    RECT 241.4000 90.8000 241.8000 93.1000 ;
	    RECT 242.2000 90.8000 242.6000 92.1000 ;
	    RECT 243.8000 90.8000 244.2000 92.1000 ;
	    RECT 244.6000 90.8000 245.0000 92.1000 ;
	    RECT 246.2000 90.8000 246.6000 92.1000 ;
	    RECT 247.0000 90.8000 247.4000 92.1000 ;
	    RECT 248.6000 90.8000 249.0000 92.1000 ;
	    RECT 250.2000 90.8000 250.6000 93.3000 ;
	    RECT 252.8000 90.8000 253.2000 93.5000 ;
	    RECT 254.2000 90.8000 254.6000 92.1000 ;
	    RECT 255.8000 90.8000 256.2000 92.1000 ;
	    RECT 257.4000 91.1000 257.9000 92.8000 ;
	    RECT 257.5000 90.8000 257.9000 91.1000 ;
	    RECT 260.5000 90.8000 261.0000 92.8000 ;
	    RECT 263.0000 90.8000 263.5000 92.8000 ;
	    RECT 266.1000 91.1000 266.6000 92.8000 ;
	    RECT 266.1000 90.8000 266.5000 91.1000 ;
	    RECT 267.8000 90.8000 268.2000 92.1000 ;
	    RECT 269.4000 90.8000 269.8000 92.1000 ;
	    RECT 0.2000 90.2000 271.0000 90.8000 ;
	    RECT 2.2000 88.3000 2.6000 90.2000 ;
	    RECT 4.6000 88.9000 5.0000 90.2000 ;
	    RECT 4.6000 88.1000 5.0000 88.6000 ;
	    RECT 5.6000 88.2000 6.0000 90.2000 ;
	    RECT 5.4000 88.1000 6.0000 88.2000 ;
	    RECT 4.6000 87.9000 6.0000 88.1000 ;
	    RECT 8.6000 87.9000 9.0000 90.2000 ;
	    RECT 10.2000 88.9000 10.6000 90.2000 ;
	    RECT 11.9000 89.9000 12.3000 90.2000 ;
	    RECT 4.6000 87.8000 5.8000 87.9000 ;
	    RECT 10.2000 87.8000 10.6000 88.6000 ;
	    RECT 11.8000 88.2000 12.3000 89.9000 ;
	    RECT 14.9000 88.2000 15.4000 90.2000 ;
	    RECT 18.2000 87.9000 18.6000 90.2000 ;
	    RECT 19.0000 88.9000 19.4000 90.2000 ;
	    RECT 20.6000 88.9000 21.0000 90.2000 ;
	    RECT 22.3000 89.9000 22.7000 90.2000 ;
	    RECT 22.2000 88.2000 22.7000 89.9000 ;
	    RECT 25.3000 88.2000 25.8000 90.2000 ;
	    RECT 27.8000 88.2000 28.3000 90.2000 ;
	    RECT 30.9000 89.9000 31.3000 90.2000 ;
	    RECT 33.5000 89.9000 33.9000 90.2000 ;
	    RECT 30.9000 88.2000 31.4000 89.9000 ;
	    RECT 33.4000 88.2000 33.9000 89.9000 ;
	    RECT 36.5000 88.2000 37.0000 90.2000 ;
	    RECT 39.0000 88.0000 39.4000 90.2000 ;
	    RECT 41.8000 88.9000 42.2000 90.2000 ;
	    RECT 43.4000 88.9000 43.9000 90.2000 ;
	    RECT 46.2000 87.9000 46.6000 90.2000 ;
	    RECT 47.8000 88.9000 48.2000 90.2000 ;
	    RECT 49.4000 88.9000 49.8000 90.2000 ;
	    RECT 28.5000 87.4000 28.9000 87.8000 ;
	    RECT 29.8000 87.7000 30.6000 87.8000 ;
	    RECT 29.8000 87.4000 30.8000 87.7000 ;
	    RECT 28.5000 87.2000 28.8000 87.4000 ;
	    RECT 10.2000 87.1000 10.6000 87.2000 ;
	    RECT 11.0000 87.1000 11.8000 87.2000 ;
	    RECT 10.2000 87.0000 12.1000 87.1000 ;
	    RECT 10.2000 86.8000 13.2000 87.0000 ;
	    RECT 25.8000 86.8000 26.6000 87.2000 ;
	    RECT 28.4000 86.8000 28.8000 87.2000 ;
	    RECT 30.5000 87.2000 30.8000 87.4000 ;
	    RECT 30.5000 86.9000 32.2000 87.2000 ;
	    RECT 31.4000 86.8000 32.2000 86.9000 ;
	    RECT 37.0000 86.8000 37.8000 87.2000 ;
	    RECT 52.6000 86.9000 53.0000 90.2000 ;
	    RECT 54.2000 88.1000 54.6000 90.2000 ;
	    RECT 55.8000 88.9000 56.2000 90.2000 ;
	    RECT 58.2000 87.9000 58.6000 90.2000 ;
	    RECT 62.2000 88.3000 62.6000 90.2000 ;
	    RECT 66.2000 86.9000 66.6000 90.2000 ;
	    RECT 67.8000 88.0000 68.2000 90.2000 ;
	    RECT 70.6000 88.9000 71.0000 90.2000 ;
	    RECT 72.2000 88.9000 72.7000 90.2000 ;
	    RECT 75.0000 87.9000 75.4000 90.2000 ;
	    RECT 76.6000 88.9000 77.0000 90.2000 ;
	    RECT 78.2000 88.9000 78.6000 90.2000 ;
	    RECT 79.8000 87.9000 80.2000 90.2000 ;
	    RECT 82.5000 88.9000 83.0000 90.2000 ;
	    RECT 84.2000 88.9000 84.6000 90.2000 ;
	    RECT 87.0000 88.0000 87.4000 90.2000 ;
	    RECT 89.4000 88.0000 89.8000 90.2000 ;
	    RECT 92.2000 88.9000 92.6000 90.2000 ;
	    RECT 93.8000 88.9000 94.3000 90.2000 ;
	    RECT 96.6000 87.9000 97.0000 90.2000 ;
	    RECT 99.0000 88.3000 99.4000 90.2000 ;
	    RECT 101.4000 87.9000 101.8000 90.2000 ;
	    RECT 103.0000 87.9000 103.4000 90.2000 ;
	    RECT 104.6000 87.9000 105.0000 90.2000 ;
	    RECT 106.2000 87.9000 106.6000 90.2000 ;
	    RECT 107.8000 87.9000 108.2000 90.2000 ;
	    RECT 110.2000 88.9000 110.6000 90.2000 ;
	    RECT 112.3000 87.9000 112.7000 90.2000 ;
	    RECT 113.4000 86.9000 113.8000 90.2000 ;
	    RECT 116.6000 88.9000 117.0000 90.2000 ;
	    RECT 119.8000 87.9000 120.2000 90.2000 ;
	    RECT 121.4000 88.0000 121.8000 90.2000 ;
	    RECT 124.2000 88.9000 124.6000 90.2000 ;
	    RECT 125.8000 88.9000 126.3000 90.2000 ;
	    RECT 128.6000 87.9000 129.0000 90.2000 ;
	    RECT 130.2000 88.9000 130.6000 90.2000 ;
	    RECT 131.8000 88.9000 132.2000 90.2000 ;
	    RECT 132.6000 88.9000 133.0000 90.2000 ;
	    RECT 134.2000 88.9000 134.6000 90.2000 ;
	    RECT 135.8000 88.9000 136.2000 90.2000 ;
	    RECT 137.4000 87.9000 137.8000 90.2000 ;
	    RECT 140.1000 88.9000 140.6000 90.2000 ;
	    RECT 141.8000 88.9000 142.2000 90.2000 ;
	    RECT 144.6000 88.0000 145.0000 90.2000 ;
	    RECT 147.0000 88.0000 147.4000 90.2000 ;
	    RECT 149.8000 88.9000 150.2000 90.2000 ;
	    RECT 151.4000 88.9000 151.9000 90.2000 ;
	    RECT 154.2000 87.9000 154.6000 90.2000 ;
	    RECT 155.8000 87.9000 156.2000 90.2000 ;
	    RECT 159.8000 88.3000 160.2000 90.2000 ;
	    RECT 163.0000 88.9000 163.4000 90.2000 ;
	    RECT 165.1000 87.9000 165.5000 90.2000 ;
	    RECT 166.2000 88.9000 166.6000 90.2000 ;
	    RECT 167.8000 87.9000 168.2000 90.2000 ;
	    RECT 171.8000 87.9000 172.2000 90.2000 ;
	    RECT 173.4000 87.9000 173.8000 90.2000 ;
	    RECT 176.1000 88.9000 176.6000 90.2000 ;
	    RECT 177.8000 88.9000 178.2000 90.2000 ;
	    RECT 180.6000 88.0000 181.0000 90.2000 ;
	    RECT 183.0000 88.9000 183.4000 90.2000 ;
	    RECT 183.8000 88.9000 184.2000 90.2000 ;
	    RECT 185.4000 88.9000 185.8000 90.2000 ;
	    RECT 187.8000 87.9000 188.2000 90.2000 ;
	    RECT 188.6000 88.9000 189.0000 90.2000 ;
	    RECT 190.7000 87.9000 191.1000 90.2000 ;
	    RECT 191.8000 88.9000 192.2000 90.2000 ;
	    RECT 193.4000 88.9000 193.8000 90.2000 ;
	    RECT 196.6000 86.9000 197.0000 90.2000 ;
	    RECT 197.4000 88.9000 197.8000 90.2000 ;
	    RECT 199.0000 88.9000 199.4000 90.2000 ;
	    RECT 200.6000 88.9000 201.0000 90.2000 ;
	    RECT 202.2000 88.3000 202.6000 90.2000 ;
	    RECT 206.2000 87.9000 206.6000 90.2000 ;
	    RECT 207.0000 88.9000 207.4000 90.2000 ;
	    RECT 208.6000 88.9000 209.0000 90.2000 ;
	    RECT 209.4000 88.9000 209.8000 90.2000 ;
	    RECT 213.4000 88.3000 213.8000 90.2000 ;
	    RECT 217.4000 88.3000 217.8000 90.2000 ;
	    RECT 219.0000 88.9000 219.4000 90.2000 ;
	    RECT 221.1000 87.9000 221.5000 90.2000 ;
	    RECT 223.0000 88.3000 223.4000 90.2000 ;
	    RECT 226.2000 88.3000 226.6000 90.2000 ;
	    RECT 229.4000 88.9000 229.8000 90.2000 ;
	    RECT 231.0000 88.9000 231.4000 90.2000 ;
	    RECT 232.7000 89.9000 233.1000 90.2000 ;
	    RECT 232.6000 88.2000 233.1000 89.9000 ;
	    RECT 235.7000 88.2000 236.2000 90.2000 ;
	    RECT 237.4000 88.9000 237.8000 90.2000 ;
	    RECT 239.0000 87.9000 239.4000 90.2000 ;
	    RECT 240.6000 87.9000 241.0000 90.2000 ;
	    RECT 241.4000 88.9000 241.8000 90.2000 ;
	    RECT 243.8000 88.3000 244.2000 90.2000 ;
	    RECT 247.0000 88.3000 247.4000 90.2000 ;
	    RECT 249.4000 88.9000 249.8000 90.2000 ;
	    RECT 251.0000 88.9000 251.4000 90.2000 ;
	    RECT 252.6000 88.3000 253.0000 90.2000 ;
	    RECT 255.8000 88.3000 256.2000 90.2000 ;
	    RECT 259.1000 89.9000 259.5000 90.2000 ;
	    RECT 259.0000 88.2000 259.5000 89.9000 ;
	    RECT 262.1000 88.2000 262.6000 90.2000 ;
	    RECT 264.6000 88.2000 265.1000 90.2000 ;
	    RECT 267.7000 89.9000 268.1000 90.2000 ;
	    RECT 267.7000 88.2000 268.2000 89.9000 ;
	    RECT 11.8000 86.7000 13.2000 86.8000 ;
	    RECT 12.8000 86.6000 13.2000 86.7000 ;
	    RECT 3.1000 74.4000 3.5000 74.8000 ;
	    RECT 3.1000 74.2000 3.4000 74.4000 ;
	    RECT 3.0000 74.1000 3.4000 74.2000 ;
	    RECT 2.2000 73.8000 3.4000 74.1000 ;
	    RECT 4.6000 74.1000 5.0000 74.6000 ;
	    RECT 7.0000 74.4000 7.4000 75.2000 ;
	    RECT 8.6000 74.4000 9.0000 75.2000 ;
	    RECT 38.8000 74.3000 39.2000 74.4000 ;
	    RECT 38.8000 74.2000 40.2000 74.3000 ;
	    RECT 5.4000 74.1000 5.8000 74.2000 ;
	    RECT 4.6000 73.8000 5.8000 74.1000 ;
	    RECT 38.8000 74.0000 41.0000 74.2000 ;
	    RECT 39.9000 73.9000 41.0000 74.0000 ;
	    RECT 40.2000 73.8000 41.0000 73.9000 ;
	    RECT 2.2000 73.1000 2.5000 73.8000 ;
	    RECT 0.6000 70.8000 1.0000 72.1000 ;
	    RECT 2.2000 70.8000 2.6000 73.1000 ;
	    RECT 5.2000 72.2000 5.6000 73.1000 ;
	    RECT 5.2000 71.8000 5.8000 72.2000 ;
	    RECT 5.2000 70.8000 5.6000 71.8000 ;
	    RECT 8.6000 70.8000 9.0000 72.7000 ;
	    RECT 11.8000 72.4000 12.2000 73.2000 ;
	    RECT 11.0000 70.8000 11.4000 72.1000 ;
	    RECT 11.8000 70.8000 12.2000 72.1000 ;
	    RECT 13.4000 70.8000 13.8000 73.1000 ;
	    RECT 16.4000 70.8000 16.8000 73.1000 ;
	    RECT 19.0000 70.8000 19.4000 72.7000 ;
	    RECT 21.4000 72.4000 21.8000 73.2000 ;
	    RECT 21.4000 70.8000 21.8000 72.1000 ;
	    RECT 22.2000 70.8000 22.6000 73.1000 ;
	    RECT 25.9000 70.8000 26.3000 73.0000 ;
	    RECT 28.6000 70.8000 29.0000 72.7000 ;
	    RECT 32.6000 70.8000 33.0000 73.1000 ;
	    RECT 33.4000 70.8000 33.8000 72.1000 ;
	    RECT 35.0000 70.8000 35.4000 72.1000 ;
	    RECT 36.6000 70.8000 37.1000 72.8000 ;
	    RECT 39.7000 71.1000 40.2000 72.8000 ;
	    RECT 39.7000 70.8000 40.1000 71.1000 ;
	    RECT 41.4000 70.8000 41.8000 72.1000 ;
	    RECT 44.6000 70.8000 45.0000 72.7000 ;
	    RECT 46.4000 70.8000 46.8000 73.1000 ;
	    RECT 49.4000 70.8000 49.8000 73.1000 ;
	    RECT 51.0000 70.8000 51.4000 72.1000 ;
	    RECT 52.6000 70.8000 53.0000 72.7000 ;
	    RECT 55.0000 70.8000 55.4000 74.1000 ;
	    RECT 60.6000 70.8000 61.0000 73.0000 ;
	    RECT 63.4000 70.8000 63.8000 72.1000 ;
	    RECT 65.0000 70.8000 65.5000 72.1000 ;
	    RECT 67.8000 70.8000 68.2000 73.1000 ;
	    RECT 69.4000 70.8000 69.8000 72.1000 ;
	    RECT 71.5000 70.8000 71.9000 73.1000 ;
	    RECT 74.2000 70.8000 74.6000 72.7000 ;
	    RECT 77.4000 70.8000 77.8000 72.7000 ;
	    RECT 79.8000 70.8000 80.2000 73.0000 ;
	    RECT 82.6000 70.8000 83.0000 72.1000 ;
	    RECT 84.2000 70.8000 84.7000 72.1000 ;
	    RECT 87.0000 70.8000 87.4000 73.1000 ;
	    RECT 89.4000 70.8000 89.8000 72.1000 ;
	    RECT 91.8000 70.8000 92.2000 73.1000 ;
	    RECT 93.4000 70.8000 93.8000 72.7000 ;
	    RECT 95.8000 70.8000 96.2000 72.1000 ;
	    RECT 97.4000 70.8000 97.8000 72.1000 ;
	    RECT 98.2000 70.8000 98.6000 73.1000 ;
	    RECT 99.8000 70.8000 100.2000 73.1000 ;
	    RECT 101.7000 70.8000 102.1000 73.1000 ;
	    RECT 103.8000 70.8000 104.2000 72.1000 ;
	    RECT 107.0000 70.8000 107.4000 73.1000 ;
	    RECT 109.7000 70.8000 110.2000 72.1000 ;
	    RECT 111.4000 70.8000 111.8000 72.1000 ;
	    RECT 114.2000 70.8000 114.6000 73.0000 ;
	    RECT 116.6000 70.8000 117.0000 73.1000 ;
	    RECT 118.2000 70.8000 118.6000 73.1000 ;
	    RECT 119.8000 70.8000 120.2000 73.1000 ;
	    RECT 122.5000 70.8000 123.0000 72.1000 ;
	    RECT 124.2000 70.8000 124.6000 72.1000 ;
	    RECT 127.0000 70.8000 127.4000 73.0000 ;
	    RECT 129.4000 70.8000 129.8000 73.0000 ;
	    RECT 132.2000 70.8000 132.6000 72.1000 ;
	    RECT 133.8000 70.8000 134.3000 72.1000 ;
	    RECT 136.6000 70.8000 137.0000 73.1000 ;
	    RECT 139.0000 70.8000 139.4000 73.1000 ;
	    RECT 140.6000 70.8000 141.0000 73.1000 ;
	    RECT 142.2000 70.8000 142.6000 72.7000 ;
	    RECT 144.6000 70.8000 145.0000 73.1000 ;
	    RECT 146.2000 70.8000 146.6000 73.1000 ;
	    RECT 147.8000 70.8000 148.2000 73.1000 ;
	    RECT 149.4000 70.8000 149.8000 73.1000 ;
	    RECT 151.0000 70.8000 151.4000 73.1000 ;
	    RECT 151.8000 70.8000 152.2000 73.1000 ;
	    RECT 153.4000 70.8000 153.8000 73.1000 ;
	    RECT 155.0000 70.8000 155.4000 73.1000 ;
	    RECT 156.6000 70.8000 157.0000 73.1000 ;
	    RECT 158.2000 70.8000 158.6000 73.1000 ;
	    RECT 161.9000 70.8000 162.3000 73.0000 ;
	    RECT 163.8000 70.8000 164.2000 73.1000 ;
	    RECT 167.0000 70.8000 167.4000 72.1000 ;
	    RECT 168.6000 70.8000 169.0000 73.1000 ;
	    RECT 171.3000 70.8000 171.8000 72.1000 ;
	    RECT 173.0000 70.8000 173.4000 72.1000 ;
	    RECT 175.8000 70.8000 176.2000 73.0000 ;
	    RECT 179.0000 70.8000 179.4000 73.1000 ;
	    RECT 179.8000 70.8000 180.2000 72.1000 ;
	    RECT 181.9000 70.8000 182.3000 73.1000 ;
	    RECT 185.4000 70.8000 185.8000 74.1000 ;
	    RECT 186.2000 70.8000 186.6000 72.1000 ;
	    RECT 187.8000 70.8000 188.2000 72.1000 ;
	    RECT 190.2000 70.8000 190.6000 73.1000 ;
	    RECT 191.0000 70.8000 191.4000 72.1000 ;
	    RECT 192.6000 70.8000 193.0000 72.9000 ;
	    RECT 195.8000 70.8000 196.2000 72.7000 ;
	    RECT 198.2000 70.8000 198.6000 72.9000 ;
	    RECT 199.8000 70.8000 200.2000 72.1000 ;
	    RECT 200.6000 70.8000 201.0000 72.1000 ;
	    RECT 202.2000 70.8000 202.6000 72.1000 ;
	    RECT 204.6000 70.8000 205.0000 73.1000 ;
	    RECT 205.4000 70.8000 205.8000 72.1000 ;
	    RECT 207.5000 70.8000 207.9000 73.1000 ;
	    RECT 211.0000 70.8000 211.4000 73.1000 ;
	    RECT 213.7000 70.8000 214.2000 72.1000 ;
	    RECT 215.4000 70.8000 215.8000 72.1000 ;
	    RECT 218.2000 70.8000 218.6000 73.0000 ;
	    RECT 220.6000 70.8000 221.0000 72.1000 ;
	    RECT 221.4000 70.8000 221.8000 72.1000 ;
	    RECT 223.8000 70.8000 224.2000 72.1000 ;
	    RECT 225.4000 70.8000 225.8000 72.7000 ;
	    RECT 227.8000 70.8000 228.2000 74.1000 ;
	    RECT 231.8000 70.8000 232.2000 72.7000 ;
	    RECT 235.8000 70.8000 236.2000 72.7000 ;
	    RECT 237.4000 70.8000 237.8000 72.1000 ;
	    RECT 239.0000 70.8000 239.4000 72.1000 ;
	    RECT 240.6000 70.8000 241.0000 72.1000 ;
	    RECT 241.4000 70.8000 241.8000 73.1000 ;
	    RECT 243.8000 70.8000 244.2000 72.1000 ;
	    RECT 245.4000 70.8000 245.8000 72.1000 ;
	    RECT 247.0000 71.1000 247.5000 72.8000 ;
	    RECT 247.1000 70.8000 247.5000 71.1000 ;
	    RECT 250.1000 70.8000 250.6000 72.8000 ;
	    RECT 254.2000 70.8000 254.6000 74.1000 ;
	    RECT 256.6000 70.8000 257.0000 73.1000 ;
	    RECT 259.0000 70.8000 259.4000 72.7000 ;
	    RECT 262.2000 70.8000 262.6000 72.7000 ;
	    RECT 263.8000 70.8000 264.2000 72.1000 ;
	    RECT 265.4000 70.8000 265.8000 72.1000 ;
	    RECT 266.2000 70.8000 266.6000 73.1000 ;
	    RECT 269.4000 70.8000 269.8000 72.1000 ;
	    RECT 0.2000 70.2000 271.0000 70.8000 ;
	    RECT 0.6000 68.9000 1.0000 70.2000 ;
	    RECT 2.2000 67.9000 2.6000 70.2000 ;
	    RECT 4.6000 68.9000 5.0000 70.2000 ;
	    RECT 6.2000 68.9000 6.6000 70.2000 ;
	    RECT 7.0000 68.9000 7.4000 70.2000 ;
	    RECT 6.2000 67.8000 6.6000 68.6000 ;
	    RECT 9.1000 67.9000 9.5000 70.2000 ;
	    RECT 11.8000 68.3000 12.2000 70.2000 ;
	    RECT 13.4000 68.9000 13.8000 70.2000 ;
	    RECT 15.0000 68.9000 15.4000 70.2000 ;
	    RECT 16.1000 67.9000 16.5000 70.2000 ;
	    RECT 18.2000 68.9000 18.6000 70.2000 ;
	    RECT 20.6000 67.9000 21.0000 70.2000 ;
	    RECT 21.7000 67.9000 22.1000 70.2000 ;
	    RECT 23.8000 68.9000 24.2000 70.2000 ;
	    RECT 24.6000 68.9000 25.0000 70.2000 ;
	    RECT 26.2000 68.9000 26.6000 70.2000 ;
	    RECT 27.0000 68.9000 27.4000 70.2000 ;
	    RECT 29.1000 67.9000 29.5000 70.2000 ;
	    RECT 30.2000 67.9000 30.6000 70.2000 ;
	    RECT 33.4000 68.9000 33.8000 70.2000 ;
	    RECT 35.8000 67.9000 36.2000 70.2000 ;
	    RECT 39.0000 68.3000 39.4000 70.2000 ;
	    RECT 2.2000 66.8000 2.6000 67.6000 ;
	    RECT 43.0000 66.9000 43.4000 70.2000 ;
	    RECT 45.4000 67.9000 45.8000 70.2000 ;
	    RECT 47.0000 68.9000 47.4000 70.2000 ;
	    RECT 47.8000 68.9000 48.2000 70.2000 ;
	    RECT 49.4000 68.9000 49.8000 70.2000 ;
	    RECT 51.0000 67.9000 51.4000 70.2000 ;
	    RECT 53.7000 68.9000 54.2000 70.2000 ;
	    RECT 55.4000 68.9000 55.8000 70.2000 ;
	    RECT 58.2000 68.0000 58.6000 70.2000 ;
	    RECT 61.4000 68.9000 61.8000 70.2000 ;
	    RECT 63.0000 68.9000 63.4000 70.2000 ;
	    RECT 63.8000 66.9000 64.2000 70.2000 ;
	    RECT 67.8000 68.3000 68.2000 70.2000 ;
	    RECT 70.2000 68.9000 70.6000 70.2000 ;
	    RECT 71.8000 68.9000 72.2000 70.2000 ;
	    RECT 73.4000 67.9000 73.8000 70.2000 ;
	    RECT 76.1000 68.9000 76.6000 70.2000 ;
	    RECT 77.8000 68.9000 78.2000 70.2000 ;
	    RECT 80.6000 68.0000 81.0000 70.2000 ;
	    RECT 83.8000 68.3000 84.2000 70.2000 ;
	    RECT 85.4000 68.9000 85.8000 70.2000 ;
	    RECT 87.5000 67.9000 87.9000 70.2000 ;
	    RECT 88.6000 66.9000 89.0000 70.2000 ;
	    RECT 91.8000 67.9000 92.2000 70.2000 ;
	    RECT 93.4000 67.9000 93.8000 70.2000 ;
	    RECT 95.0000 67.9000 95.4000 70.2000 ;
	    RECT 96.6000 67.9000 97.0000 70.2000 ;
	    RECT 98.2000 67.9000 98.6000 70.2000 ;
	    RECT 99.8000 67.9000 100.2000 70.2000 ;
	    RECT 101.4000 67.9000 101.8000 70.2000 ;
	    RECT 103.0000 67.9000 103.4000 70.2000 ;
	    RECT 104.6000 67.9000 105.0000 70.2000 ;
	    RECT 106.2000 67.9000 106.6000 70.2000 ;
	    RECT 110.2000 67.9000 110.6000 70.2000 ;
	    RECT 111.8000 67.9000 112.2000 70.2000 ;
	    RECT 113.4000 67.9000 113.8000 70.2000 ;
	    RECT 115.0000 67.9000 115.4000 70.2000 ;
	    RECT 115.8000 66.9000 116.2000 70.2000 ;
	    RECT 119.0000 68.9000 119.4000 70.2000 ;
	    RECT 121.1000 67.9000 121.5000 70.2000 ;
	    RECT 123.8000 68.3000 124.2000 70.2000 ;
	    RECT 127.0000 68.3000 127.4000 70.2000 ;
	    RECT 129.4000 67.9000 129.8000 70.2000 ;
	    RECT 131.0000 67.9000 131.4000 70.2000 ;
	    RECT 132.6000 67.9000 133.0000 70.2000 ;
	    RECT 134.2000 67.9000 134.6000 70.2000 ;
	    RECT 135.0000 67.9000 135.4000 70.2000 ;
	    RECT 136.6000 67.9000 137.0000 70.2000 ;
	    RECT 138.2000 67.9000 138.6000 70.2000 ;
	    RECT 140.6000 68.3000 141.0000 70.2000 ;
	    RECT 142.5000 67.9000 142.9000 70.2000 ;
	    RECT 144.6000 68.9000 145.0000 70.2000 ;
	    RECT 146.2000 68.3000 146.6000 70.2000 ;
	    RECT 148.9000 67.9000 149.3000 70.2000 ;
	    RECT 151.0000 68.9000 151.4000 70.2000 ;
	    RECT 152.6000 68.0000 153.0000 70.2000 ;
	    RECT 155.4000 68.9000 155.8000 70.2000 ;
	    RECT 157.0000 68.9000 157.5000 70.2000 ;
	    RECT 159.8000 67.9000 160.2000 70.2000 ;
	    RECT 163.0000 67.9000 163.4000 70.2000 ;
	    RECT 166.2000 68.9000 166.6000 70.2000 ;
	    RECT 167.0000 67.9000 167.4000 70.2000 ;
	    RECT 168.6000 67.9000 169.0000 70.2000 ;
	    RECT 171.0000 67.9000 171.4000 70.2000 ;
	    RECT 172.6000 67.9000 173.0000 70.2000 ;
	    RECT 174.2000 68.9000 174.6000 70.2000 ;
	    RECT 175.0000 68.9000 175.4000 70.2000 ;
	    RECT 178.2000 67.9000 178.6000 70.2000 ;
	    RECT 179.8000 67.7000 180.2000 70.2000 ;
	    RECT 182.4000 67.5000 182.8000 70.2000 ;
	    RECT 183.8000 68.9000 184.2000 70.2000 ;
	    RECT 185.4000 68.9000 185.8000 70.2000 ;
	    RECT 186.2000 68.9000 186.6000 70.2000 ;
	    RECT 187.8000 68.1000 188.2000 70.2000 ;
	    RECT 190.0000 67.5000 190.4000 70.2000 ;
	    RECT 192.6000 67.7000 193.0000 70.2000 ;
	    RECT 195.0000 68.2000 195.5000 70.2000 ;
	    RECT 198.1000 69.9000 198.5000 70.2000 ;
	    RECT 198.1000 68.2000 198.6000 69.9000 ;
	    RECT 200.6000 67.9000 201.0000 70.2000 ;
	    RECT 202.2000 67.9000 202.6000 70.2000 ;
	    RECT 205.4000 68.9000 205.8000 70.2000 ;
	    RECT 206.2000 67.9000 206.6000 70.2000 ;
	    RECT 207.8000 67.9000 208.2000 70.2000 ;
	    RECT 208.6000 68.9000 209.0000 70.2000 ;
	    RECT 210.2000 68.9000 210.6000 70.2000 ;
	    RECT 212.6000 68.9000 213.0000 70.2000 ;
	    RECT 214.2000 68.9000 214.6000 70.2000 ;
	    RECT 217.4000 66.9000 217.8000 70.2000 ;
	    RECT 218.2000 67.9000 218.6000 70.2000 ;
	    RECT 220.6000 68.9000 221.0000 70.2000 ;
	    RECT 222.7000 67.9000 223.1000 70.2000 ;
	    RECT 224.6000 68.3000 225.0000 70.2000 ;
	    RECT 227.0000 67.9000 227.4000 70.2000 ;
	    RECT 231.0000 68.3000 231.4000 70.2000 ;
	    RECT 232.6000 68.9000 233.0000 70.2000 ;
	    RECT 235.8000 68.3000 236.2000 70.2000 ;
	    RECT 238.2000 68.3000 238.6000 70.2000 ;
	    RECT 240.9000 67.9000 241.3000 70.2000 ;
	    RECT 243.0000 68.9000 243.4000 70.2000 ;
	    RECT 243.8000 68.9000 244.2000 70.2000 ;
	    RECT 245.4000 68.9000 245.8000 70.2000 ;
	    RECT 247.0000 66.9000 247.4000 70.2000 ;
	    RECT 250.2000 68.9000 250.6000 70.2000 ;
	    RECT 251.8000 68.9000 252.2000 70.2000 ;
	    RECT 253.4000 68.3000 253.8000 70.2000 ;
	    RECT 256.6000 68.9000 257.0000 70.2000 ;
	    RECT 258.3000 69.9000 258.7000 70.2000 ;
	    RECT 258.2000 68.2000 258.7000 69.9000 ;
	    RECT 261.3000 68.2000 261.8000 70.2000 ;
	    RECT 263.0000 67.9000 263.4000 70.2000 ;
	    RECT 264.6000 67.9000 265.0000 70.2000 ;
	    RECT 267.0000 67.9000 267.4000 70.2000 ;
	    RECT 268.6000 67.9000 269.0000 70.2000 ;
	    RECT 201.4000 65.8000 201.8000 66.6000 ;
	    RECT 152.6000 54.4000 153.0000 55.2000 ;
	    RECT 200.6000 55.1000 201.0000 55.2000 ;
	    RECT 200.6000 54.8000 203.1000 55.1000 ;
	    RECT 202.7000 54.7000 203.1000 54.8000 ;
	    RECT 5.0000 53.8000 5.8000 54.2000 ;
	    RECT 23.8000 53.4000 24.2000 54.2000 ;
	    RECT 1.4000 51.1000 1.9000 52.8000 ;
	    RECT 1.5000 50.8000 1.9000 51.1000 ;
	    RECT 4.5000 50.8000 5.0000 52.8000 ;
	    RECT 9.4000 52.4000 9.8000 53.2000 ;
	    RECT 6.2000 50.8000 6.6000 52.1000 ;
	    RECT 7.8000 50.8000 8.2000 52.1000 ;
	    RECT 9.4000 50.8000 9.8000 52.1000 ;
	    RECT 10.2000 50.8000 10.6000 52.1000 ;
	    RECT 13.4000 50.8000 13.8000 52.7000 ;
	    RECT 16.6000 52.4000 17.0000 53.2000 ;
	    RECT 15.0000 50.8000 15.4000 52.1000 ;
	    RECT 16.6000 50.8000 17.0000 52.1000 ;
	    RECT 18.2000 50.8000 18.6000 52.1000 ;
	    RECT 19.0000 50.8000 19.4000 52.1000 ;
	    RECT 21.1000 50.8000 21.5000 53.1000 ;
	    RECT 23.8000 50.8000 24.2000 53.1000 ;
	    RECT 25.4000 51.1000 25.9000 52.8000 ;
	    RECT 25.5000 50.8000 25.9000 51.1000 ;
	    RECT 28.5000 50.8000 29.0000 52.8000 ;
	    RECT 31.8000 50.8000 32.2000 52.7000 ;
	    RECT 33.4000 50.8000 33.8000 52.1000 ;
	    RECT 36.6000 50.8000 37.0000 53.1000 ;
	    RECT 37.7000 50.8000 38.1000 53.1000 ;
	    RECT 42.2000 52.4000 42.6000 53.2000 ;
	    RECT 39.8000 50.8000 40.2000 52.1000 ;
	    RECT 40.6000 50.8000 41.0000 52.1000 ;
	    RECT 42.2000 50.8000 42.6000 52.1000 ;
	    RECT 43.8000 50.8000 44.2000 53.0000 ;
	    RECT 46.6000 50.8000 47.0000 52.1000 ;
	    RECT 48.2000 50.8000 48.7000 52.1000 ;
	    RECT 51.0000 50.8000 51.4000 53.1000 ;
	    RECT 53.4000 50.8000 53.8000 52.9000 ;
	    RECT 55.0000 50.8000 55.4000 52.1000 ;
	    RECT 58.2000 50.8000 58.6000 53.0000 ;
	    RECT 61.0000 50.8000 61.4000 52.1000 ;
	    RECT 62.6000 50.8000 63.1000 52.1000 ;
	    RECT 65.4000 50.8000 65.8000 53.1000 ;
	    RECT 67.0000 50.8000 67.4000 52.1000 ;
	    RECT 69.1000 50.8000 69.5000 53.1000 ;
	    RECT 71.8000 50.8000 72.2000 52.7000 ;
	    RECT 75.0000 50.8000 75.4000 52.7000 ;
	    RECT 76.9000 50.8000 77.3000 53.1000 ;
	    RECT 79.0000 50.8000 79.4000 52.1000 ;
	    RECT 82.2000 50.8000 82.6000 54.1000 ;
	    RECT 83.8000 50.8000 84.2000 53.0000 ;
	    RECT 86.6000 50.8000 87.0000 52.1000 ;
	    RECT 88.2000 50.8000 88.7000 52.1000 ;
	    RECT 91.0000 50.8000 91.4000 53.1000 ;
	    RECT 92.6000 50.8000 93.0000 53.1000 ;
	    RECT 94.2000 50.8000 94.6000 53.1000 ;
	    RECT 95.8000 50.8000 96.2000 53.1000 ;
	    RECT 97.4000 50.8000 97.8000 53.1000 ;
	    RECT 100.3000 50.8000 100.7000 53.0000 ;
	    RECT 102.2000 50.8000 102.6000 53.1000 ;
	    RECT 104.6000 50.8000 105.0000 53.1000 ;
	    RECT 106.2000 50.8000 106.6000 53.1000 ;
	    RECT 110.2000 50.8000 110.6000 53.0000 ;
	    RECT 113.0000 50.8000 113.4000 52.1000 ;
	    RECT 114.6000 50.8000 115.1000 52.1000 ;
	    RECT 117.4000 50.8000 117.8000 53.1000 ;
	    RECT 119.0000 50.8000 119.4000 52.1000 ;
	    RECT 121.1000 50.8000 121.5000 53.1000 ;
	    RECT 122.2000 50.8000 122.6000 54.1000 ;
	    RECT 125.4000 50.8000 125.8000 53.1000 ;
	    RECT 127.0000 50.8000 127.4000 52.1000 ;
	    RECT 129.4000 50.8000 129.8000 52.7000 ;
	    RECT 132.1000 50.8000 132.5000 53.1000 ;
	    RECT 134.2000 50.8000 134.6000 52.1000 ;
	    RECT 135.8000 50.8000 136.2000 53.1000 ;
	    RECT 138.5000 50.8000 139.0000 52.1000 ;
	    RECT 140.2000 50.8000 140.6000 52.1000 ;
	    RECT 143.0000 50.8000 143.4000 53.0000 ;
	    RECT 147.0000 50.8000 147.4000 54.1000 ;
	    RECT 147.8000 50.8000 148.2000 54.1000 ;
	    RECT 151.8000 50.8000 152.2000 53.1000 ;
	    RECT 153.7000 50.8000 154.1000 53.1000 ;
	    RECT 155.8000 50.8000 156.2000 52.1000 ;
	    RECT 157.4000 50.8000 157.8000 52.7000 ;
	    RECT 162.2000 50.8000 162.6000 53.1000 ;
	    RECT 164.9000 50.8000 165.4000 52.1000 ;
	    RECT 166.6000 50.8000 167.0000 52.1000 ;
	    RECT 169.4000 50.8000 169.8000 53.0000 ;
	    RECT 171.0000 50.8000 171.4000 53.1000 ;
	    RECT 173.4000 50.8000 173.8000 52.1000 ;
	    RECT 175.5000 50.8000 175.9000 53.1000 ;
	    RECT 176.6000 50.8000 177.0000 52.1000 ;
	    RECT 178.2000 50.8000 178.6000 53.1000 ;
	    RECT 180.6000 50.8000 181.0000 52.1000 ;
	    RECT 182.7000 50.8000 183.1000 53.1000 ;
	    RECT 184.6000 50.8000 185.0000 53.1000 ;
	    RECT 187.3000 50.8000 187.8000 52.1000 ;
	    RECT 189.0000 50.8000 189.4000 52.1000 ;
	    RECT 191.8000 50.8000 192.2000 53.0000 ;
	    RECT 194.2000 50.8000 194.6000 52.1000 ;
	    RECT 195.8000 50.8000 196.2000 53.0000 ;
	    RECT 198.6000 50.8000 199.0000 52.1000 ;
	    RECT 200.2000 50.8000 200.7000 52.1000 ;
	    RECT 203.0000 50.8000 203.4000 53.1000 ;
	    RECT 204.6000 50.8000 205.0000 52.1000 ;
	    RECT 206.7000 50.8000 207.1000 53.1000 ;
	    RECT 210.2000 50.8000 210.6000 53.1000 ;
	    RECT 212.9000 50.8000 213.4000 52.1000 ;
	    RECT 214.6000 50.8000 215.0000 52.1000 ;
	    RECT 217.4000 50.8000 217.8000 53.0000 ;
	    RECT 219.8000 50.8000 220.2000 53.1000 ;
	    RECT 222.5000 50.8000 223.0000 52.1000 ;
	    RECT 224.2000 50.8000 224.6000 52.1000 ;
	    RECT 227.0000 50.8000 227.4000 53.0000 ;
	    RECT 228.6000 50.8000 229.0000 52.1000 ;
	    RECT 230.2000 50.8000 230.6000 52.1000 ;
	    RECT 232.3000 50.8000 232.7000 53.0000 ;
	    RECT 235.0000 50.8000 235.4000 53.0000 ;
	    RECT 237.8000 50.8000 238.2000 52.1000 ;
	    RECT 239.4000 50.8000 239.9000 52.1000 ;
	    RECT 242.2000 50.8000 242.6000 53.1000 ;
	    RECT 243.8000 50.8000 244.2000 52.1000 ;
	    RECT 246.7000 50.8000 247.1000 53.0000 ;
	    RECT 249.4000 50.8000 249.8000 52.1000 ;
	    RECT 251.0000 50.8000 251.4000 51.9000 ;
	    RECT 255.0000 50.8000 255.4000 52.1000 ;
	    RECT 256.6000 50.8000 257.0000 52.1000 ;
	    RECT 257.4000 50.8000 257.8000 52.1000 ;
	    RECT 259.5000 50.8000 259.9000 53.1000 ;
	    RECT 261.4000 50.8000 261.8000 52.7000 ;
	    RECT 263.8000 50.8000 264.2000 52.1000 ;
	    RECT 265.4000 50.8000 265.8000 53.1000 ;
	    RECT 267.8000 50.8000 268.2000 52.1000 ;
	    RECT 269.4000 50.8000 269.8000 52.1000 ;
	    RECT 0.2000 50.2000 271.0000 50.8000 ;
	    RECT 1.4000 48.2000 1.9000 50.2000 ;
	    RECT 4.5000 49.9000 4.9000 50.2000 ;
	    RECT 4.5000 48.2000 5.0000 49.9000 ;
	    RECT 6.2000 47.9000 6.6000 50.2000 ;
	    RECT 8.6000 48.9000 9.0000 50.2000 ;
	    RECT 10.7000 47.9000 11.1000 50.2000 ;
	    RECT 12.6000 48.9000 13.0000 50.2000 ;
	    RECT 13.4000 48.8000 13.8000 50.2000 ;
	    RECT 15.0000 48.9000 15.4000 50.2000 ;
	    RECT 17.4000 47.9000 17.8000 50.2000 ;
	    RECT 19.1000 49.9000 19.5000 50.2000 ;
	    RECT 19.0000 48.2000 19.5000 49.9000 ;
	    RECT 22.1000 48.2000 22.6000 50.2000 ;
	    RECT 23.8000 48.9000 24.2000 50.2000 ;
	    RECT 27.0000 47.9000 27.4000 50.2000 ;
	    RECT 27.8000 48.9000 28.2000 50.2000 ;
	    RECT 29.4000 48.9000 29.8000 50.2000 ;
	    RECT 31.0000 48.9000 31.4000 50.2000 ;
	    RECT 32.7000 49.9000 33.1000 50.2000 ;
	    RECT 32.6000 48.2000 33.1000 49.9000 ;
	    RECT 35.7000 48.2000 36.2000 50.2000 ;
	    RECT 38.2000 48.9000 38.6000 50.2000 ;
	    RECT 39.0000 47.9000 39.4000 50.2000 ;
	    RECT 41.4000 48.9000 41.8000 50.2000 ;
	    RECT 43.8000 48.0000 44.2000 50.2000 ;
	    RECT 46.6000 48.9000 47.0000 50.2000 ;
	    RECT 48.2000 48.9000 48.7000 50.2000 ;
	    RECT 51.0000 47.9000 51.4000 50.2000 ;
	    RECT 53.4000 48.1000 53.8000 50.2000 ;
	    RECT 55.0000 48.9000 55.4000 50.2000 ;
	    RECT 56.6000 47.9000 57.0000 50.2000 ;
	    RECT 58.2000 47.9000 58.6000 50.2000 ;
	    RECT 60.6000 48.9000 61.0000 50.2000 ;
	    RECT 65.4000 49.1000 65.8000 50.2000 ;
	    RECT 67.0000 48.9000 67.4000 50.2000 ;
	    RECT 68.6000 48.9000 69.0000 50.2000 ;
	    RECT 70.2000 48.9000 70.6000 50.2000 ;
	    RECT 71.8000 48.9000 72.2000 50.2000 ;
	    RECT 72.6000 48.9000 73.0000 50.2000 ;
	    RECT 74.2000 48.9000 74.6000 50.2000 ;
	    RECT 75.8000 48.9000 76.2000 50.2000 ;
	    RECT 78.2000 48.3000 78.6000 50.2000 ;
	    RECT 80.6000 47.9000 81.0000 50.2000 ;
	    RECT 83.3000 48.9000 83.8000 50.2000 ;
	    RECT 85.0000 48.9000 85.4000 50.2000 ;
	    RECT 87.8000 48.0000 88.2000 50.2000 ;
	    RECT 91.0000 48.3000 91.4000 50.2000 ;
	    RECT 92.9000 47.9000 93.3000 50.2000 ;
	    RECT 95.0000 48.9000 95.4000 50.2000 ;
	    RECT 96.1000 47.9000 96.5000 50.2000 ;
	    RECT 98.2000 48.9000 98.6000 50.2000 ;
	    RECT 100.6000 48.3000 101.0000 50.2000 ;
	    RECT 103.0000 48.3000 103.4000 50.2000 ;
	    RECT 105.7000 47.9000 106.1000 50.2000 ;
	    RECT 107.8000 48.9000 108.2000 50.2000 ;
	    RECT 0.6000 46.8000 1.4000 47.2000 ;
	    RECT 22.6000 46.8000 23.4000 47.2000 ;
	    RECT 39.0000 46.8000 39.4000 47.6000 ;
	    RECT 112.6000 46.9000 113.0000 50.2000 ;
	    RECT 114.2000 48.0000 114.6000 50.2000 ;
	    RECT 117.0000 48.9000 117.4000 50.2000 ;
	    RECT 118.6000 48.9000 119.1000 50.2000 ;
	    RECT 121.4000 47.9000 121.8000 50.2000 ;
	    RECT 123.0000 47.9000 123.4000 50.2000 ;
	    RECT 125.4000 48.9000 125.8000 50.2000 ;
	    RECT 127.0000 48.9000 127.4000 50.2000 ;
	    RECT 127.8000 48.9000 128.2000 50.2000 ;
	    RECT 129.9000 47.9000 130.3000 50.2000 ;
	    RECT 132.3000 48.0000 132.7000 50.2000 ;
	    RECT 134.2000 47.9000 134.6000 50.2000 ;
	    RECT 135.8000 47.9000 136.2000 50.2000 ;
	    RECT 137.4000 47.9000 137.8000 50.2000 ;
	    RECT 139.0000 47.9000 139.4000 50.2000 ;
	    RECT 140.6000 47.9000 141.0000 50.2000 ;
	    RECT 142.2000 47.9000 142.6000 50.2000 ;
	    RECT 144.9000 48.9000 145.4000 50.2000 ;
	    RECT 146.6000 48.9000 147.0000 50.2000 ;
	    RECT 149.4000 48.0000 149.8000 50.2000 ;
	    RECT 151.8000 47.9000 152.2000 50.2000 ;
	    RECT 154.5000 48.9000 155.0000 50.2000 ;
	    RECT 156.2000 48.9000 156.6000 50.2000 ;
	    RECT 159.0000 48.0000 159.4000 50.2000 ;
	    RECT 162.2000 48.9000 162.6000 50.2000 ;
	    RECT 163.8000 48.9000 164.2000 50.2000 ;
	    RECT 165.4000 48.9000 165.8000 50.2000 ;
	    RECT 167.0000 48.0000 167.4000 50.2000 ;
	    RECT 169.8000 48.9000 170.2000 50.2000 ;
	    RECT 171.4000 48.9000 171.9000 50.2000 ;
	    RECT 174.2000 47.9000 174.6000 50.2000 ;
	    RECT 175.8000 48.9000 176.2000 50.2000 ;
	    RECT 178.2000 48.0000 178.6000 50.2000 ;
	    RECT 181.0000 48.9000 181.4000 50.2000 ;
	    RECT 182.6000 48.9000 183.1000 50.2000 ;
	    RECT 185.4000 47.9000 185.8000 50.2000 ;
	    RECT 188.3000 48.0000 188.7000 50.2000 ;
	    RECT 191.0000 47.9000 191.4000 50.2000 ;
	    RECT 193.7000 48.9000 194.2000 50.2000 ;
	    RECT 195.4000 48.9000 195.8000 50.2000 ;
	    RECT 198.2000 48.0000 198.6000 50.2000 ;
	    RECT 200.9000 48.0000 201.3000 50.2000 ;
	    RECT 203.8000 48.3000 204.2000 50.2000 ;
	    RECT 207.0000 47.9000 207.4000 50.2000 ;
	    RECT 211.0000 47.9000 211.4000 50.2000 ;
	    RECT 213.7000 48.9000 214.2000 50.2000 ;
	    RECT 215.4000 48.9000 215.8000 50.2000 ;
	    RECT 218.2000 48.0000 218.6000 50.2000 ;
	    RECT 220.6000 47.9000 221.0000 50.2000 ;
	    RECT 223.3000 48.9000 223.8000 50.2000 ;
	    RECT 225.0000 48.9000 225.4000 50.2000 ;
	    RECT 227.8000 48.0000 228.2000 50.2000 ;
	    RECT 230.2000 48.0000 230.6000 50.2000 ;
	    RECT 233.0000 48.9000 233.4000 50.2000 ;
	    RECT 234.6000 48.9000 235.1000 50.2000 ;
	    RECT 237.4000 47.9000 237.8000 50.2000 ;
	    RECT 239.8000 48.0000 240.2000 50.2000 ;
	    RECT 242.6000 48.9000 243.0000 50.2000 ;
	    RECT 244.2000 48.9000 244.7000 50.2000 ;
	    RECT 247.0000 47.9000 247.4000 50.2000 ;
	    RECT 249.4000 48.3000 249.8000 50.2000 ;
	    RECT 253.4000 48.3000 253.8000 50.2000 ;
	    RECT 255.3000 47.9000 255.7000 50.2000 ;
	    RECT 257.4000 48.9000 257.8000 50.2000 ;
	    RECT 259.0000 48.0000 259.4000 50.2000 ;
	    RECT 261.8000 48.9000 262.2000 50.2000 ;
	    RECT 263.4000 48.9000 263.9000 50.2000 ;
	    RECT 266.2000 47.9000 266.6000 50.2000 ;
	    RECT 269.4000 47.9000 269.8000 50.2000 ;
	    RECT 13.4000 45.4000 13.8000 46.2000 ;
	    RECT 249.4000 45.8000 249.8000 46.6000 ;
	    RECT 7.8000 44.4000 8.2000 45.2000 ;
	    RECT 251.0000 45.1000 251.4000 45.2000 ;
	    RECT 250.7000 44.8000 251.4000 45.1000 ;
	    RECT 250.7000 44.2000 251.0000 44.8000 ;
	    RECT 250.6000 43.8000 251.0000 44.2000 ;
	    RECT 23.0000 34.8000 23.4000 35.6000 ;
	    RECT 235.4000 35.2000 235.8000 35.4000 ;
	    RECT 235.0000 34.9000 235.8000 35.2000 ;
	    RECT 235.0000 34.8000 235.4000 34.9000 ;
	    RECT 251.0000 34.8000 251.4000 35.6000 ;
	    RECT 5.0000 33.8000 5.8000 34.2000 ;
	    RECT 10.6000 34.1000 11.4000 34.2000 ;
	    RECT 11.8000 34.1000 12.2000 34.2000 ;
	    RECT 10.6000 33.8000 12.2000 34.1000 ;
	    RECT 35.8000 33.8000 36.6000 34.2000 ;
	    RECT 1.4000 31.1000 1.9000 32.8000 ;
	    RECT 1.5000 30.8000 1.9000 31.1000 ;
	    RECT 4.5000 30.8000 5.0000 32.8000 ;
	    RECT 7.0000 31.1000 7.5000 32.8000 ;
	    RECT 7.1000 30.8000 7.5000 31.1000 ;
	    RECT 10.1000 30.8000 10.6000 32.8000 ;
	    RECT 11.8000 32.4000 12.2000 33.2000 ;
	    RECT 11.8000 30.8000 12.2000 32.1000 ;
	    RECT 13.4000 30.8000 13.8000 33.1000 ;
	    RECT 15.8000 30.8000 16.2000 32.1000 ;
	    RECT 17.4000 30.8000 17.8000 32.1000 ;
	    RECT 19.8000 30.8000 20.2000 32.7000 ;
	    RECT 21.4000 30.8000 21.8000 32.1000 ;
	    RECT 23.0000 30.8000 23.4000 32.2000 ;
	    RECT 23.8000 30.8000 24.2000 32.1000 ;
	    RECT 26.2000 30.8000 26.6000 32.7000 ;
	    RECT 28.6000 30.8000 29.0000 32.1000 ;
	    RECT 30.2000 30.8000 30.6000 32.1000 ;
	    RECT 31.0000 30.8000 31.4000 32.1000 ;
	    RECT 32.6000 30.8000 33.0000 32.1000 ;
	    RECT 35.0000 30.8000 35.4000 33.1000 ;
	    RECT 36.6000 30.8000 37.1000 32.8000 ;
	    RECT 39.7000 31.1000 40.2000 32.8000 ;
	    RECT 39.7000 30.8000 40.1000 31.1000 ;
	    RECT 41.4000 30.8000 41.8000 32.1000 ;
	    RECT 43.0000 30.8000 43.4000 32.1000 ;
	    RECT 44.6000 30.8000 45.0000 32.1000 ;
	    RECT 45.4000 30.8000 45.8000 33.1000 ;
	    RECT 47.0000 30.8000 47.4000 33.1000 ;
	    RECT 48.6000 30.8000 49.0000 33.1000 ;
	    RECT 51.0000 30.8000 51.4000 33.0000 ;
	    RECT 53.8000 30.8000 54.2000 32.1000 ;
	    RECT 55.4000 30.8000 55.9000 32.1000 ;
	    RECT 58.2000 30.8000 58.6000 33.1000 ;
	    RECT 63.8000 30.8000 64.2000 34.1000 ;
	    RECT 64.6000 30.8000 65.0000 33.1000 ;
	    RECT 67.0000 30.8000 67.4000 32.1000 ;
	    RECT 69.4000 30.8000 69.8000 32.7000 ;
	    RECT 72.6000 30.8000 73.0000 33.0000 ;
	    RECT 75.4000 30.8000 75.8000 32.1000 ;
	    RECT 77.0000 30.8000 77.5000 32.1000 ;
	    RECT 79.8000 30.8000 80.2000 33.1000 ;
	    RECT 81.4000 30.8000 81.8000 34.1000 ;
	    RECT 84.6000 30.8000 85.0000 34.1000 ;
	    RECT 91.0000 30.8000 91.4000 31.9000 ;
	    RECT 92.6000 30.8000 93.0000 32.1000 ;
	    RECT 95.0000 30.8000 95.4000 32.1000 ;
	    RECT 97.4000 30.8000 97.8000 32.7000 ;
	    RECT 99.8000 30.8000 100.2000 32.7000 ;
	    RECT 103.0000 30.8000 103.4000 32.7000 ;
	    RECT 107.8000 30.8000 108.2000 33.1000 ;
	    RECT 110.5000 30.8000 111.0000 32.1000 ;
	    RECT 112.2000 30.8000 112.6000 32.1000 ;
	    RECT 115.0000 30.8000 115.4000 33.0000 ;
	    RECT 117.4000 30.8000 117.8000 32.7000 ;
	    RECT 119.8000 30.8000 120.2000 33.1000 ;
	    RECT 122.8000 30.8000 123.2000 33.1000 ;
	    RECT 123.8000 30.8000 124.2000 34.1000 ;
	    RECT 248.6000 33.4000 249.0000 34.2000 ;
	    RECT 127.8000 30.8000 128.2000 33.1000 ;
	    RECT 130.5000 30.8000 131.0000 32.1000 ;
	    RECT 132.2000 30.8000 132.6000 32.1000 ;
	    RECT 135.0000 30.8000 135.4000 33.0000 ;
	    RECT 137.9000 30.8000 138.3000 33.0000 ;
	    RECT 140.6000 30.8000 141.0000 32.9000 ;
	    RECT 142.2000 30.8000 142.6000 32.1000 ;
	    RECT 143.8000 30.8000 144.2000 33.1000 ;
	    RECT 146.5000 30.8000 147.0000 32.1000 ;
	    RECT 148.2000 30.8000 148.6000 32.1000 ;
	    RECT 151.0000 30.8000 151.4000 33.0000 ;
	    RECT 152.6000 30.8000 153.0000 33.1000 ;
	    RECT 155.0000 30.8000 155.4000 33.1000 ;
	    RECT 158.2000 30.8000 158.6000 32.1000 ;
	    RECT 161.4000 30.8000 161.8000 33.0000 ;
	    RECT 164.2000 30.8000 164.6000 32.1000 ;
	    RECT 165.8000 30.8000 166.3000 32.1000 ;
	    RECT 168.6000 30.8000 169.0000 33.1000 ;
	    RECT 170.2000 30.8000 170.6000 32.1000 ;
	    RECT 171.8000 30.8000 172.2000 32.1000 ;
	    RECT 173.4000 30.8000 173.8000 32.1000 ;
	    RECT 175.0000 30.8000 175.4000 32.1000 ;
	    RECT 176.6000 30.8000 177.0000 33.1000 ;
	    RECT 178.2000 30.8000 178.6000 33.1000 ;
	    RECT 179.8000 30.8000 180.2000 33.1000 ;
	    RECT 182.5000 30.8000 183.0000 32.1000 ;
	    RECT 184.2000 30.8000 184.6000 32.1000 ;
	    RECT 187.0000 30.8000 187.4000 33.0000 ;
	    RECT 188.9000 30.8000 189.3000 33.1000 ;
	    RECT 191.0000 30.8000 191.4000 32.1000 ;
	    RECT 192.6000 30.8000 193.0000 32.7000 ;
	    RECT 195.8000 30.8000 196.2000 33.1000 ;
	    RECT 198.5000 30.8000 199.0000 32.1000 ;
	    RECT 200.2000 30.8000 200.6000 32.1000 ;
	    RECT 203.0000 30.8000 203.4000 33.0000 ;
	    RECT 205.9000 30.8000 206.3000 33.0000 ;
	    RECT 210.2000 30.8000 210.6000 33.1000 ;
	    RECT 212.9000 30.8000 213.4000 32.1000 ;
	    RECT 214.6000 30.8000 215.0000 32.1000 ;
	    RECT 217.4000 30.8000 217.8000 33.0000 ;
	    RECT 220.3000 30.8000 220.7000 33.0000 ;
	    RECT 223.0000 30.8000 223.4000 33.1000 ;
	    RECT 225.7000 30.8000 226.2000 32.1000 ;
	    RECT 227.4000 30.8000 227.8000 32.1000 ;
	    RECT 230.2000 30.8000 230.6000 33.0000 ;
	    RECT 233.4000 30.8000 233.8000 32.7000 ;
	    RECT 235.3000 32.2000 235.7000 33.1000 ;
	    RECT 235.0000 31.8000 235.7000 32.2000 ;
	    RECT 235.3000 30.8000 235.7000 31.8000 ;
	    RECT 237.4000 30.8000 237.8000 32.1000 ;
	    RECT 239.8000 30.8000 240.2000 32.7000 ;
	    RECT 241.4000 32.4000 241.8000 33.2000 ;
	    RECT 241.4000 30.8000 241.8000 32.1000 ;
	    RECT 243.0000 30.8000 243.4000 32.1000 ;
	    RECT 243.8000 30.8000 244.2000 32.1000 ;
	    RECT 245.9000 30.8000 246.3000 33.1000 ;
	    RECT 247.0000 30.8000 247.4000 33.1000 ;
	    RECT 248.6000 30.8000 249.0000 33.1000 ;
	    RECT 249.4000 32.4000 249.8000 33.2000 ;
	    RECT 249.4000 30.8000 249.8000 32.1000 ;
	    RECT 251.0000 30.8000 251.4000 32.2000 ;
	    RECT 251.8000 30.8000 252.2000 32.1000 ;
	    RECT 254.2000 30.8000 254.6000 32.7000 ;
	    RECT 257.7000 30.8000 258.1000 33.0000 ;
	    RECT 260.6000 30.8000 261.0000 32.7000 ;
	    RECT 263.8000 30.8000 264.2000 32.1000 ;
	    RECT 264.6000 30.8000 265.0000 32.1000 ;
	    RECT 266.7000 30.8000 267.1000 33.1000 ;
	    RECT 267.8000 30.8000 268.2000 32.1000 ;
	    RECT 0.2000 30.2000 271.0000 30.8000 ;
	    RECT 0.6000 28.9000 1.0000 30.2000 ;
	    RECT 2.2000 28.9000 2.6000 30.2000 ;
	    RECT 3.8000 28.9000 4.2000 30.2000 ;
	    RECT 3.8000 27.8000 4.2000 28.6000 ;
	    RECT 4.6000 27.9000 5.0000 30.2000 ;
	    RECT 7.3000 27.9000 7.7000 30.2000 ;
	    RECT 9.4000 28.9000 9.8000 30.2000 ;
	    RECT 10.2000 28.9000 10.6000 30.2000 ;
	    RECT 11.8000 28.9000 12.2000 30.2000 ;
	    RECT 13.4000 28.9000 13.8000 30.2000 ;
	    RECT 11.8000 27.8000 12.2000 28.6000 ;
	    RECT 14.2000 27.9000 14.6000 30.2000 ;
	    RECT 16.6000 28.9000 17.0000 30.2000 ;
	    RECT 18.7000 27.9000 19.1000 30.2000 ;
	    RECT 20.6000 28.9000 21.0000 30.2000 ;
	    RECT 23.0000 27.9000 23.4000 30.2000 ;
	    RECT 25.4000 28.3000 25.8000 30.2000 ;
	    RECT 27.0000 28.9000 27.4000 30.2000 ;
	    RECT 28.6000 28.9000 29.0000 30.2000 ;
	    RECT 29.4000 27.9000 29.8000 30.2000 ;
	    RECT 32.6000 28.9000 33.0000 30.2000 ;
	    RECT 32.6000 27.8000 33.0000 28.6000 ;
	    RECT 34.2000 27.9000 34.6000 30.2000 ;
	    RECT 36.9000 28.9000 37.4000 30.2000 ;
	    RECT 38.6000 28.9000 39.0000 30.2000 ;
	    RECT 41.4000 28.0000 41.8000 30.2000 ;
	    RECT 43.8000 27.9000 44.2000 30.2000 ;
	    RECT 46.5000 28.9000 47.0000 30.2000 ;
	    RECT 48.2000 28.9000 48.6000 30.2000 ;
	    RECT 51.0000 28.0000 51.4000 30.2000 ;
	    RECT 52.6000 28.9000 53.0000 30.2000 ;
	    RECT 54.2000 28.9000 54.6000 30.2000 ;
	    RECT 55.8000 28.9000 56.2000 30.2000 ;
	    RECT 59.0000 27.9000 59.4000 30.2000 ;
	    RECT 61.7000 28.9000 62.2000 30.2000 ;
	    RECT 63.4000 28.9000 63.8000 30.2000 ;
	    RECT 66.2000 28.0000 66.6000 30.2000 ;
	    RECT 68.6000 28.3000 69.0000 30.2000 ;
	    RECT 71.0000 28.9000 71.4000 30.2000 ;
	    RECT 72.6000 28.9000 73.0000 30.2000 ;
	    RECT 74.2000 27.9000 74.6000 30.2000 ;
	    RECT 76.9000 28.9000 77.4000 30.2000 ;
	    RECT 78.6000 28.9000 79.0000 30.2000 ;
	    RECT 81.4000 28.0000 81.8000 30.2000 ;
	    RECT 83.8000 28.0000 84.2000 30.2000 ;
	    RECT 86.6000 28.9000 87.0000 30.2000 ;
	    RECT 88.2000 28.9000 88.7000 30.2000 ;
	    RECT 91.0000 27.9000 91.4000 30.2000 ;
	    RECT 92.6000 28.9000 93.0000 30.2000 ;
	    RECT 94.2000 28.9000 94.6000 30.2000 ;
	    RECT 96.6000 27.9000 97.0000 30.2000 ;
	    RECT 97.7000 27.9000 98.1000 30.2000 ;
	    RECT 99.8000 28.9000 100.2000 30.2000 ;
	    RECT 100.6000 27.9000 101.0000 30.2000 ;
	    RECT 103.8000 27.9000 104.2000 30.2000 ;
	    RECT 105.4000 28.3000 105.8000 30.2000 ;
	    RECT 109.7000 27.9000 110.1000 30.2000 ;
	    RECT 111.8000 28.9000 112.2000 30.2000 ;
	    RECT 113.4000 27.9000 113.8000 30.2000 ;
	    RECT 116.1000 28.9000 116.6000 30.2000 ;
	    RECT 117.8000 28.9000 118.2000 30.2000 ;
	    RECT 120.6000 28.0000 121.0000 30.2000 ;
	    RECT 122.2000 28.9000 122.6000 30.2000 ;
	    RECT 125.4000 27.9000 125.8000 30.2000 ;
	    RECT 126.2000 28.9000 126.6000 30.2000 ;
	    RECT 127.8000 28.9000 128.2000 30.2000 ;
	    RECT 129.4000 28.1000 129.8000 30.2000 ;
	    RECT 131.0000 28.9000 131.4000 30.2000 ;
	    RECT 131.8000 28.9000 132.2000 30.2000 ;
	    RECT 133.4000 28.9000 133.8000 30.2000 ;
	    RECT 135.8000 27.9000 136.2000 30.2000 ;
	    RECT 138.2000 28.3000 138.6000 30.2000 ;
	    RECT 140.6000 28.9000 141.0000 30.2000 ;
	    RECT 142.2000 28.0000 142.6000 30.2000 ;
	    RECT 145.0000 28.9000 145.4000 30.2000 ;
	    RECT 146.6000 28.9000 147.1000 30.2000 ;
	    RECT 149.4000 27.9000 149.8000 30.2000 ;
	    RECT 151.3000 27.9000 151.7000 30.2000 ;
	    RECT 153.4000 28.9000 153.8000 30.2000 ;
	    RECT 155.0000 27.9000 155.4000 30.2000 ;
	    RECT 157.7000 28.9000 158.2000 30.2000 ;
	    RECT 159.4000 28.9000 159.8000 30.2000 ;
	    RECT 162.2000 28.0000 162.6000 30.2000 ;
	    RECT 166.2000 28.3000 166.6000 30.2000 ;
	    RECT 169.4000 27.9000 169.8000 30.2000 ;
	    RECT 172.1000 28.9000 172.6000 30.2000 ;
	    RECT 173.8000 28.9000 174.2000 30.2000 ;
	    RECT 176.6000 28.0000 177.0000 30.2000 ;
	    RECT 178.2000 28.9000 178.6000 30.2000 ;
	    RECT 179.8000 28.9000 180.2000 30.2000 ;
	    RECT 181.4000 28.9000 181.8000 30.2000 ;
	    RECT 182.2000 27.9000 182.6000 30.2000 ;
	    RECT 183.8000 27.9000 184.2000 30.2000 ;
	    RECT 185.4000 27.9000 185.8000 30.2000 ;
	    RECT 187.0000 27.9000 187.4000 30.2000 ;
	    RECT 188.6000 27.9000 189.0000 30.2000 ;
	    RECT 190.2000 27.9000 190.6000 30.2000 ;
	    RECT 192.9000 28.9000 193.4000 30.2000 ;
	    RECT 194.6000 28.9000 195.0000 30.2000 ;
	    RECT 197.4000 28.0000 197.8000 30.2000 ;
	    RECT 199.0000 27.9000 199.4000 30.2000 ;
	    RECT 4.6000 26.8000 5.0000 27.6000 ;
	    RECT 201.2000 27.5000 201.6000 30.2000 ;
	    RECT 203.8000 27.7000 204.2000 30.2000 ;
	    RECT 206.5000 28.0000 206.9000 30.2000 ;
	    RECT 209.4000 28.3000 209.8000 30.2000 ;
	    RECT 214.2000 28.9000 214.6000 30.2000 ;
	    RECT 216.6000 27.9000 217.0000 30.2000 ;
	    RECT 217.4000 27.9000 217.8000 30.2000 ;
	    RECT 220.6000 27.9000 221.0000 30.2000 ;
	    RECT 221.4000 27.9000 221.8000 30.2000 ;
	    RECT 223.8000 28.9000 224.2000 30.2000 ;
	    RECT 225.4000 28.9000 225.8000 30.2000 ;
	    RECT 223.8000 27.8000 224.2000 28.6000 ;
	    RECT 227.0000 28.3000 227.4000 30.2000 ;
	    RECT 229.7000 27.9000 230.1000 30.2000 ;
	    RECT 231.8000 28.9000 232.2000 30.2000 ;
	    RECT 234.2000 27.9000 234.6000 30.2000 ;
	    RECT 236.6000 28.3000 237.0000 30.2000 ;
	    RECT 238.5000 27.9000 238.9000 30.2000 ;
	    RECT 240.6000 28.9000 241.0000 30.2000 ;
	    RECT 241.4000 27.9000 241.8000 30.2000 ;
	    RECT 243.0000 27.9000 243.4000 30.2000 ;
	    RECT 244.7000 29.9000 245.1000 30.2000 ;
	    RECT 244.6000 28.2000 245.1000 29.9000 ;
	    RECT 247.7000 28.2000 248.2000 30.2000 ;
	    RECT 250.2000 27.9000 250.6000 30.2000 ;
	    RECT 252.9000 28.9000 253.4000 30.2000 ;
	    RECT 254.6000 28.9000 255.0000 30.2000 ;
	    RECT 257.4000 28.0000 257.8000 30.2000 ;
	    RECT 259.0000 28.9000 259.4000 30.2000 ;
	    RECT 261.4000 27.9000 261.8000 30.2000 ;
	    RECT 264.1000 28.9000 264.6000 30.2000 ;
	    RECT 265.8000 28.9000 266.2000 30.2000 ;
	    RECT 268.6000 28.0000 269.0000 30.2000 ;
	    RECT 220.6000 26.8000 221.0000 27.6000 ;
	    RECT 15.8000 24.4000 16.2000 25.2000 ;
	    RECT 194.6000 16.8000 195.0000 17.2000 ;
	    RECT 194.7000 16.2000 195.0000 16.8000 ;
	    RECT 194.7000 15.9000 195.4000 16.2000 ;
	    RECT 195.0000 15.8000 195.4000 15.9000 ;
	    RECT 218.2000 15.8000 218.6000 17.2000 ;
	    RECT 27.8000 14.4000 28.2000 15.2000 ;
	    RECT 187.0000 14.8000 187.4000 15.6000 ;
	    RECT 259.4000 15.2000 259.8000 15.4000 ;
	    RECT 190.2000 14.8000 190.6000 15.2000 ;
	    RECT 190.3000 14.4000 190.6000 14.8000 ;
	    RECT 215.0000 14.4000 215.4000 15.2000 ;
	    RECT 259.4000 14.9000 260.2000 15.2000 ;
	    RECT 259.8000 14.8000 260.2000 14.9000 ;
	    RECT 190.2000 14.0000 190.8000 14.4000 ;
	    RECT 1.4000 10.8000 1.8000 12.1000 ;
	    RECT 2.2000 10.8000 2.6000 12.1000 ;
	    RECT 3.8000 10.8000 4.2000 12.1000 ;
	    RECT 5.4000 10.8000 5.8000 13.0000 ;
	    RECT 8.2000 10.8000 8.6000 12.1000 ;
	    RECT 9.8000 10.8000 10.3000 12.1000 ;
	    RECT 12.6000 10.8000 13.0000 13.1000 ;
	    RECT 14.2000 10.8000 14.6000 12.1000 ;
	    RECT 15.8000 10.8000 16.2000 12.1000 ;
	    RECT 17.4000 10.8000 17.8000 12.1000 ;
	    RECT 19.0000 10.8000 19.4000 13.0000 ;
	    RECT 21.8000 10.8000 22.2000 12.1000 ;
	    RECT 23.4000 10.8000 23.9000 12.1000 ;
	    RECT 26.2000 10.8000 26.6000 13.1000 ;
	    RECT 28.6000 10.8000 29.0000 13.1000 ;
	    RECT 31.0000 10.8000 31.4000 13.1000 ;
	    RECT 33.7000 10.8000 34.2000 12.1000 ;
	    RECT 35.4000 10.8000 35.8000 12.1000 ;
	    RECT 38.2000 10.8000 38.6000 13.0000 ;
	    RECT 40.6000 10.8000 41.0000 12.9000 ;
	    RECT 42.2000 10.8000 42.6000 12.1000 ;
	    RECT 43.0000 10.8000 43.4000 12.1000 ;
	    RECT 44.6000 10.8000 45.0000 12.1000 ;
	    RECT 46.2000 10.8000 46.6000 12.1000 ;
	    RECT 47.0000 10.8000 47.4000 12.1000 ;
	    RECT 48.6000 10.8000 49.0000 12.1000 ;
	    RECT 50.2000 10.8000 50.6000 12.1000 ;
	    RECT 51.8000 10.8000 52.3000 12.8000 ;
	    RECT 54.9000 11.1000 55.4000 12.8000 ;
	    RECT 54.9000 10.8000 55.3000 11.1000 ;
	    RECT 58.2000 10.8000 58.6000 12.1000 ;
	    RECT 60.3000 10.8000 60.7000 13.1000 ;
	    RECT 61.4000 10.8000 61.8000 13.1000 ;
	    RECT 65.4000 10.8000 65.8000 12.7000 ;
	    RECT 67.0000 10.8000 67.4000 12.1000 ;
	    RECT 69.4000 10.8000 69.8000 12.7000 ;
	    RECT 72.0000 10.8000 72.4000 13.1000 ;
	    RECT 75.0000 10.8000 75.4000 13.1000 ;
	    RECT 76.6000 10.8000 77.0000 12.1000 ;
	    RECT 77.4000 10.8000 77.8000 13.1000 ;
	    RECT 79.0000 10.8000 79.4000 13.1000 ;
	    RECT 80.6000 10.8000 81.0000 13.1000 ;
	    RECT 82.2000 10.8000 82.6000 13.1000 ;
	    RECT 83.8000 10.8000 84.2000 13.1000 ;
	    RECT 84.6000 10.8000 85.0000 12.1000 ;
	    RECT 86.2000 10.8000 86.6000 12.1000 ;
	    RECT 87.3000 10.8000 87.7000 13.1000 ;
	    RECT 89.4000 10.8000 89.8000 12.1000 ;
	    RECT 91.8000 10.8000 92.2000 12.7000 ;
	    RECT 93.4000 10.8000 93.8000 12.1000 ;
	    RECT 95.0000 10.8000 95.4000 12.1000 ;
	    RECT 97.4000 10.8000 97.8000 12.7000 ;
	    RECT 99.8000 10.8000 100.2000 12.1000 ;
	    RECT 100.6000 10.8000 101.0000 12.1000 ;
	    RECT 102.5000 10.8000 102.9000 13.1000 ;
	    RECT 104.6000 10.8000 105.0000 12.1000 ;
	    RECT 107.0000 10.8000 107.4000 13.1000 ;
	    RECT 111.0000 10.8000 111.4000 12.7000 ;
	    RECT 112.6000 10.8000 113.0000 12.1000 ;
	    RECT 114.2000 10.8000 114.6000 12.1000 ;
	    RECT 115.8000 10.8000 116.2000 12.1000 ;
	    RECT 116.6000 10.8000 117.0000 12.1000 ;
	    RECT 118.2000 10.8000 118.6000 12.1000 ;
	    RECT 119.0000 10.8000 119.4000 12.1000 ;
	    RECT 122.2000 10.8000 122.6000 13.1000 ;
	    RECT 123.8000 10.8000 124.2000 12.1000 ;
	    RECT 125.4000 10.8000 125.8000 13.0000 ;
	    RECT 128.2000 10.8000 128.6000 12.1000 ;
	    RECT 129.8000 10.8000 130.3000 12.1000 ;
	    RECT 132.6000 10.8000 133.0000 13.1000 ;
	    RECT 134.2000 10.8000 134.6000 12.1000 ;
	    RECT 135.8000 10.8000 136.2000 12.1000 ;
	    RECT 137.4000 10.8000 137.8000 12.1000 ;
	    RECT 139.0000 10.8000 139.5000 12.8000 ;
	    RECT 142.1000 11.1000 142.6000 12.8000 ;
	    RECT 142.1000 10.8000 142.5000 11.1000 ;
	    RECT 143.8000 10.8000 144.2000 12.1000 ;
	    RECT 145.4000 10.8000 145.8000 12.1000 ;
	    RECT 147.0000 10.8000 147.4000 12.1000 ;
	    RECT 147.8000 10.8000 148.2000 13.1000 ;
	    RECT 149.4000 10.8000 149.8000 13.1000 ;
	    RECT 151.0000 10.8000 151.4000 13.1000 ;
	    RECT 152.6000 10.8000 153.0000 13.1000 ;
	    RECT 154.2000 10.8000 154.6000 13.1000 ;
	    RECT 155.0000 10.8000 155.4000 13.1000 ;
	    RECT 156.6000 10.8000 157.0000 13.1000 ;
	    RECT 158.2000 10.8000 158.6000 12.1000 ;
	    RECT 161.4000 10.8000 161.8000 12.1000 ;
	    RECT 163.0000 10.8000 163.4000 12.1000 ;
	    RECT 163.8000 10.8000 164.2000 13.1000 ;
	    RECT 165.4000 10.8000 165.8000 13.1000 ;
	    RECT 167.0000 10.8000 167.4000 13.1000 ;
	    RECT 168.6000 10.8000 169.0000 13.1000 ;
	    RECT 170.2000 10.8000 170.6000 13.1000 ;
	    RECT 171.8000 10.8000 172.2000 13.1000 ;
	    RECT 174.2000 10.8000 174.6000 13.0000 ;
	    RECT 177.0000 10.8000 177.4000 12.1000 ;
	    RECT 178.6000 10.8000 179.1000 12.1000 ;
	    RECT 181.4000 10.8000 181.8000 13.1000 ;
	    RECT 183.0000 10.8000 183.4000 12.1000 ;
	    RECT 184.6000 10.8000 185.0000 12.1000 ;
	    RECT 186.2000 10.8000 186.6000 12.1000 ;
	    RECT 187.0000 10.8000 187.4000 12.2000 ;
	    RECT 188.6000 10.8000 189.0000 12.1000 ;
	    RECT 190.7000 10.8000 191.1000 13.0000 ;
	    RECT 193.4000 10.8000 193.8000 12.7000 ;
	    RECT 196.6000 10.8000 197.0000 13.2000 ;
	    RECT 199.3000 10.8000 199.8000 12.1000 ;
	    RECT 201.0000 10.8000 201.4000 12.1000 ;
	    RECT 203.8000 10.8000 204.2000 13.0000 ;
	    RECT 206.0000 10.8000 206.4000 13.5000 ;
	    RECT 249.4000 13.4000 249.8000 14.2000 ;
	    RECT 208.6000 10.8000 209.0000 13.3000 ;
	    RECT 210.2000 10.8000 210.6000 13.1000 ;
	    RECT 215.0000 10.8000 215.4000 12.7000 ;
	    RECT 216.6000 10.8000 217.0000 13.1000 ;
	    RECT 220.3000 10.8000 220.7000 13.0000 ;
	    RECT 222.2000 10.8000 222.6000 12.1000 ;
	    RECT 223.8000 10.8000 224.2000 12.1000 ;
	    RECT 226.2000 10.8000 226.6000 13.1000 ;
	    RECT 227.0000 12.4000 227.4000 13.2000 ;
	    RECT 227.0000 10.8000 227.4000 12.1000 ;
	    RECT 228.6000 10.8000 229.0000 12.1000 ;
	    RECT 229.4000 10.8000 229.8000 13.1000 ;
	    RECT 231.8000 10.8000 232.2000 12.1000 ;
	    RECT 233.4000 10.8000 233.8000 13.1000 ;
	    RECT 236.4000 10.8000 236.8000 13.1000 ;
	    RECT 239.0000 10.8000 239.4000 12.7000 ;
	    RECT 240.6000 10.8000 241.0000 12.1000 ;
	    RECT 242.2000 10.8000 242.6000 12.1000 ;
	    RECT 244.6000 10.8000 245.0000 13.1000 ;
	    RECT 246.2000 10.8000 246.6000 12.7000 ;
	    RECT 249.4000 10.8000 249.8000 13.1000 ;
	    RECT 250.2000 10.8000 250.6000 13.1000 ;
	    RECT 259.5000 12.2000 259.9000 13.1000 ;
	    RECT 251.8000 10.8000 252.2000 12.1000 ;
	    RECT 253.4000 10.8000 253.8000 12.1000 ;
	    RECT 255.0000 10.8000 255.4000 12.1000 ;
	    RECT 256.6000 10.8000 257.0000 12.1000 ;
	    RECT 257.4000 10.8000 257.8000 12.1000 ;
	    RECT 259.5000 11.8000 260.2000 12.2000 ;
	    RECT 259.5000 10.8000 259.9000 11.8000 ;
	    RECT 261.4000 10.8000 261.8000 13.1000 ;
	    RECT 264.1000 10.8000 264.6000 12.1000 ;
	    RECT 265.8000 10.8000 266.2000 12.1000 ;
	    RECT 268.6000 10.8000 269.0000 13.0000 ;
	    RECT 0.2000 10.2000 271.0000 10.8000 ;
	    RECT 1.4000 7.9000 1.8000 10.2000 ;
	    RECT 3.8000 7.9000 4.2000 10.2000 ;
	    RECT 5.4000 8.9000 5.8000 10.2000 ;
	    RECT 7.0000 8.9000 7.4000 10.2000 ;
	    RECT 8.6000 8.9000 9.0000 10.2000 ;
	    RECT 10.2000 8.0000 10.6000 10.2000 ;
	    RECT 13.0000 8.9000 13.4000 10.2000 ;
	    RECT 14.6000 8.9000 15.1000 10.2000 ;
	    RECT 17.4000 7.9000 17.8000 10.2000 ;
	    RECT 19.8000 7.9000 20.2000 10.2000 ;
	    RECT 21.4000 8.9000 21.8000 10.2000 ;
	    RECT 23.0000 8.9000 23.4000 10.2000 ;
	    RECT 24.6000 8.9000 25.0000 10.2000 ;
	    RECT 26.2000 7.9000 26.6000 10.2000 ;
	    RECT 28.9000 8.9000 29.4000 10.2000 ;
	    RECT 30.6000 8.9000 31.0000 10.2000 ;
	    RECT 33.4000 8.0000 33.8000 10.2000 ;
	    RECT 35.8000 7.9000 36.2000 10.2000 ;
	    RECT 37.4000 8.9000 37.8000 10.2000 ;
	    RECT 39.0000 8.9000 39.4000 10.2000 ;
	    RECT 40.6000 8.9000 41.0000 10.2000 ;
	    RECT 42.2000 7.9000 42.6000 10.2000 ;
	    RECT 44.9000 8.9000 45.4000 10.2000 ;
	    RECT 46.6000 8.9000 47.0000 10.2000 ;
	    RECT 49.4000 8.0000 49.8000 10.2000 ;
	    RECT 51.8000 7.9000 52.2000 10.2000 ;
	    RECT 54.3000 9.9000 54.7000 10.2000 ;
	    RECT 54.2000 8.2000 54.7000 9.9000 ;
	    RECT 57.3000 8.2000 57.8000 10.2000 ;
	    RECT 60.6000 8.9000 61.0000 10.2000 ;
	    RECT 62.2000 8.9000 62.6000 10.2000 ;
	    RECT 63.8000 8.9000 64.2000 10.2000 ;
	    RECT 65.4000 8.2000 65.9000 10.2000 ;
	    RECT 68.5000 9.9000 68.9000 10.2000 ;
	    RECT 71.1000 9.9000 71.5000 10.2000 ;
	    RECT 68.5000 8.2000 69.0000 9.9000 ;
	    RECT 71.0000 8.2000 71.5000 9.9000 ;
	    RECT 74.1000 8.2000 74.6000 10.2000 ;
	    RECT 75.8000 8.9000 76.2000 10.2000 ;
	    RECT 77.4000 8.9000 77.8000 10.2000 ;
	    RECT 78.2000 8.9000 78.6000 10.2000 ;
	    RECT 80.6000 8.3000 81.0000 10.2000 ;
	    RECT 84.0000 7.9000 84.4000 10.2000 ;
	    RECT 87.0000 7.9000 87.4000 10.2000 ;
	    RECT 88.6000 8.9000 89.0000 10.2000 ;
	    RECT 91.0000 7.9000 91.4000 10.2000 ;
	    RECT 91.8000 7.9000 92.2000 10.2000 ;
	    RECT 95.5000 8.0000 95.9000 10.2000 ;
	    RECT 97.4000 8.9000 97.8000 10.2000 ;
	    RECT 99.5000 7.9000 99.9000 10.2000 ;
	    RECT 100.6000 8.9000 101.0000 10.2000 ;
	    RECT 102.2000 8.9000 102.6000 10.2000 ;
	    RECT 104.6000 7.9000 105.0000 10.2000 ;
	    RECT 105.4000 8.9000 105.8000 10.2000 ;
	    RECT 107.0000 8.9000 107.4000 10.2000 ;
	    RECT 108.6000 8.9000 109.0000 10.2000 ;
	    RECT 111.8000 8.2000 112.3000 10.2000 ;
	    RECT 114.9000 9.9000 115.3000 10.2000 ;
	    RECT 114.9000 8.2000 115.4000 9.9000 ;
	    RECT 118.2000 7.9000 118.6000 10.2000 ;
	    RECT 119.8000 8.9000 120.2000 10.2000 ;
	    RECT 120.6000 8.9000 121.0000 10.2000 ;
	    RECT 122.2000 8.9000 122.6000 10.2000 ;
	    RECT 124.6000 7.9000 125.0000 10.2000 ;
	    RECT 126.2000 8.2000 126.7000 10.2000 ;
	    RECT 129.3000 9.9000 129.7000 10.2000 ;
	    RECT 129.3000 8.2000 129.8000 9.9000 ;
	    RECT 131.3000 7.9000 131.7000 10.2000 ;
	    RECT 133.4000 8.9000 133.8000 10.2000 ;
	    RECT 134.2000 8.9000 134.6000 10.2000 ;
	    RECT 135.8000 8.9000 136.2000 10.2000 ;
	    RECT 136.6000 7.9000 137.0000 10.2000 ;
	    RECT 139.8000 8.9000 140.2000 10.2000 ;
	    RECT 142.2000 7.9000 142.6000 10.2000 ;
	    RECT 143.8000 8.0000 144.2000 10.2000 ;
	    RECT 146.6000 8.9000 147.0000 10.2000 ;
	    RECT 148.2000 8.9000 148.7000 10.2000 ;
	    RECT 151.0000 7.9000 151.4000 10.2000 ;
	    RECT 153.4000 8.2000 153.9000 10.2000 ;
	    RECT 156.5000 9.9000 156.9000 10.2000 ;
	    RECT 156.5000 8.2000 157.0000 9.9000 ;
	    RECT 160.6000 8.0000 161.0000 10.2000 ;
	    RECT 163.4000 8.9000 163.8000 10.2000 ;
	    RECT 165.0000 8.9000 165.5000 10.2000 ;
	    RECT 167.8000 7.9000 168.2000 10.2000 ;
	    RECT 169.4000 8.9000 169.8000 10.2000 ;
	    RECT 171.0000 8.1000 171.4000 10.2000 ;
	    RECT 173.4000 8.0000 173.8000 10.2000 ;
	    RECT 176.2000 8.9000 176.6000 10.2000 ;
	    RECT 177.8000 8.9000 178.3000 10.2000 ;
	    RECT 180.6000 7.9000 181.0000 10.2000 ;
	    RECT 183.0000 7.9000 183.4000 10.2000 ;
	    RECT 185.4000 8.0000 185.8000 10.2000 ;
	    RECT 188.2000 8.9000 188.6000 10.2000 ;
	    RECT 189.8000 8.9000 190.3000 10.2000 ;
	    RECT 192.6000 7.9000 193.0000 10.2000 ;
	    RECT 194.2000 8.9000 194.6000 10.2000 ;
	    RECT 195.8000 8.9000 196.2000 10.2000 ;
	    RECT 197.4000 8.9000 197.8000 10.2000 ;
	    RECT 199.0000 7.9000 199.4000 10.2000 ;
	    RECT 200.6000 8.9000 201.0000 10.2000 ;
	    RECT 202.2000 8.9000 202.6000 10.2000 ;
	    RECT 203.8000 8.9000 204.2000 10.2000 ;
	    RECT 205.4000 7.9000 205.8000 10.2000 ;
	    RECT 208.1000 8.9000 208.6000 10.2000 ;
	    RECT 209.8000 8.9000 210.2000 10.2000 ;
	    RECT 212.6000 8.0000 213.0000 10.2000 ;
	    RECT 216.6000 7.9000 217.0000 10.2000 ;
	    RECT 218.2000 8.0000 218.6000 10.2000 ;
	    RECT 221.0000 8.9000 221.4000 10.2000 ;
	    RECT 222.6000 8.9000 223.1000 10.2000 ;
	    RECT 225.4000 7.9000 225.8000 10.2000 ;
	    RECT 227.0000 8.9000 227.4000 10.2000 ;
	    RECT 216.6000 6.8000 217.0000 7.6000 ;
	    RECT 229.2000 7.5000 229.6000 10.2000 ;
	    RECT 231.8000 7.7000 232.2000 10.2000 ;
	    RECT 233.4000 8.9000 233.8000 10.2000 ;
	    RECT 235.0000 8.9000 235.4000 10.2000 ;
	    RECT 236.6000 8.9000 237.0000 10.2000 ;
	    RECT 238.2000 8.9000 238.6000 10.2000 ;
	    RECT 239.0000 8.9000 239.4000 10.2000 ;
	    RECT 240.6000 8.9000 241.0000 10.2000 ;
	    RECT 241.4000 8.9000 241.8000 10.2000 ;
	    RECT 240.6000 7.8000 241.0000 8.6000 ;
	    RECT 245.4000 8.3000 245.8000 10.2000 ;
	    RECT 248.6000 7.9000 249.0000 10.2000 ;
	    RECT 249.4000 8.9000 249.8000 10.2000 ;
	    RECT 251.3000 7.9000 251.7000 10.2000 ;
	    RECT 253.4000 8.9000 253.8000 10.2000 ;
	    RECT 254.2000 8.9000 254.6000 10.2000 ;
	    RECT 255.8000 8.9000 256.2000 10.2000 ;
	    RECT 257.4000 8.9000 257.8000 10.2000 ;
	    RECT 258.2000 8.9000 258.6000 10.2000 ;
	    RECT 259.8000 8.9000 260.2000 10.2000 ;
	    RECT 258.2000 7.8000 258.6000 8.6000 ;
	    RECT 260.6000 7.9000 261.0000 10.2000 ;
	    RECT 263.3000 7.9000 263.7000 10.2000 ;
	    RECT 265.4000 8.9000 265.8000 10.2000 ;
	    RECT 267.0000 7.9000 267.4000 10.2000 ;
	    RECT 268.6000 8.9000 269.0000 10.2000 ;
	    RECT 260.6000 6.8000 261.0000 7.6000 ;
         LAYER metal2 ;
	    RECT 3.0000 174.8000 3.4000 175.2000 ;
	    RECT 4.6000 174.8000 5.0000 175.2000 ;
	    RECT 3.0000 172.2000 3.3000 174.8000 ;
	    RECT 3.0000 171.8000 3.4000 172.2000 ;
	    RECT 0.6000 170.8000 1.0000 171.2000 ;
	    RECT 0.6000 166.2000 0.9000 170.8000 ;
	    RECT 4.6000 170.2000 4.9000 174.8000 ;
	    RECT 7.8000 173.8000 8.2000 174.2000 ;
	    RECT 10.2000 173.8000 10.6000 174.2000 ;
	    RECT 12.6000 173.8000 13.0000 174.2000 ;
	    RECT 29.4000 173.8000 29.8000 174.2000 ;
	    RECT 7.8000 172.2000 8.1000 173.8000 ;
	    RECT 10.2000 172.2000 10.5000 173.8000 ;
	    RECT 12.6000 172.2000 12.9000 173.8000 ;
	    RECT 16.6000 172.8000 17.0000 173.2000 ;
	    RECT 7.8000 171.8000 8.2000 172.2000 ;
	    RECT 10.2000 171.8000 10.6000 172.2000 ;
	    RECT 12.6000 171.8000 13.0000 172.2000 ;
	    RECT 16.6000 171.2000 16.9000 172.8000 ;
	    RECT 29.4000 172.2000 29.7000 173.8000 ;
	    RECT 33.4000 172.8000 33.8000 173.2000 ;
	    RECT 37.4000 172.8000 37.8000 173.2000 ;
	    RECT 48.6000 172.8000 49.0000 173.2000 ;
	    RECT 29.4000 171.8000 29.8000 172.2000 ;
	    RECT 33.4000 171.2000 33.7000 172.8000 ;
	    RECT 37.4000 171.2000 37.7000 172.8000 ;
	    RECT 48.6000 171.2000 48.9000 172.8000 ;
	    RECT 16.6000 170.8000 17.0000 171.2000 ;
	    RECT 33.4000 170.8000 33.8000 171.2000 ;
	    RECT 37.4000 170.8000 37.8000 171.2000 ;
	    RECT 48.6000 170.8000 49.0000 171.2000 ;
	    RECT 108.0000 170.3000 109.6000 170.7000 ;
	    RECT 210.4000 170.3000 212.0000 170.7000 ;
	    RECT 4.6000 169.8000 5.0000 170.2000 ;
	    RECT 6.2000 169.8000 6.6000 170.2000 ;
	    RECT 15.8000 169.8000 16.2000 170.2000 ;
	    RECT 18.2000 169.8000 18.6000 170.2000 ;
	    RECT 6.2000 168.2000 6.5000 169.8000 ;
	    RECT 15.8000 168.2000 16.1000 169.8000 ;
	    RECT 18.2000 168.2000 18.5000 169.8000 ;
	    RECT 34.2000 168.8000 34.6000 169.2000 ;
	    RECT 49.4000 168.8000 49.8000 169.2000 ;
	    RECT 54.2000 168.8000 54.6000 169.2000 ;
	    RECT 59.8000 168.8000 60.2000 169.2000 ;
	    RECT 6.2000 167.8000 6.6000 168.2000 ;
	    RECT 15.8000 167.8000 16.2000 168.2000 ;
	    RECT 18.2000 167.8000 18.6000 168.2000 ;
	    RECT 34.2000 167.2000 34.5000 168.8000 ;
	    RECT 49.4000 167.2000 49.7000 168.8000 ;
	    RECT 54.2000 167.2000 54.5000 168.8000 ;
	    RECT 34.2000 166.8000 34.6000 167.2000 ;
	    RECT 49.4000 166.8000 49.8000 167.2000 ;
	    RECT 54.2000 166.8000 54.6000 167.2000 ;
	    RECT 59.8000 166.2000 60.1000 168.8000 ;
	    RECT 0.6000 165.8000 1.0000 166.2000 ;
	    RECT 59.8000 165.8000 60.2000 166.2000 ;
	    RECT 42.2000 154.8000 42.6000 155.2000 ;
	    RECT 11.0000 153.8000 11.4000 154.2000 ;
	    RECT 11.8000 153.8000 12.2000 154.2000 ;
	    RECT 0.6000 152.8000 1.0000 153.2000 ;
	    RECT 7.0000 152.8000 7.4000 153.2000 ;
	    RECT 0.6000 151.2000 0.9000 152.8000 ;
	    RECT 7.0000 151.2000 7.3000 152.8000 ;
	    RECT 11.0000 152.2000 11.3000 153.8000 ;
	    RECT 11.8000 152.2000 12.1000 153.8000 ;
	    RECT 42.2000 152.2000 42.5000 154.8000 ;
	    RECT 11.0000 151.8000 11.4000 152.2000 ;
	    RECT 11.8000 151.8000 12.2000 152.2000 ;
	    RECT 42.2000 151.8000 42.6000 152.2000 ;
	    RECT 0.6000 150.8000 1.0000 151.2000 ;
	    RECT 7.0000 150.8000 7.4000 151.2000 ;
	    RECT 108.0000 150.3000 109.6000 150.7000 ;
	    RECT 210.4000 150.3000 212.0000 150.7000 ;
	    RECT 3.8000 148.8000 4.2000 149.2000 ;
	    RECT 11.8000 148.8000 12.2000 149.2000 ;
	    RECT 19.8000 148.8000 20.2000 149.2000 ;
	    RECT 3.8000 147.2000 4.1000 148.8000 ;
	    RECT 3.8000 146.8000 4.2000 147.2000 ;
	    RECT 10.2000 146.8000 10.6000 147.2000 ;
	    RECT 10.2000 146.2000 10.5000 146.8000 ;
	    RECT 11.8000 146.2000 12.1000 148.8000 ;
	    RECT 19.8000 147.2000 20.1000 148.8000 ;
	    RECT 19.8000 146.8000 20.2000 147.2000 ;
	    RECT 10.2000 145.8000 10.6000 146.2000 ;
	    RECT 11.8000 145.8000 12.2000 146.2000 ;
	    RECT 15.0000 134.8000 15.4000 135.2000 ;
	    RECT 89.4000 134.8000 89.8000 135.2000 ;
	    RECT 147.8000 134.8000 148.2000 135.2000 ;
	    RECT 15.0000 134.2000 15.3000 134.8000 ;
	    RECT 5.4000 133.8000 5.8000 134.2000 ;
	    RECT 8.6000 133.8000 9.0000 134.2000 ;
	    RECT 15.0000 133.8000 15.4000 134.2000 ;
	    RECT 18.2000 133.8000 18.6000 134.2000 ;
	    RECT 5.4000 131.2000 5.7000 133.8000 ;
	    RECT 8.6000 132.2000 8.9000 133.8000 ;
	    RECT 11.0000 132.8000 11.4000 133.2000 ;
	    RECT 8.6000 131.8000 9.0000 132.2000 ;
	    RECT 11.0000 131.2000 11.3000 132.8000 ;
	    RECT 18.2000 132.1000 18.5000 133.8000 ;
	    RECT 19.0000 132.1000 19.4000 132.2000 ;
	    RECT 18.2000 131.8000 19.4000 132.1000 ;
	    RECT 3.0000 130.8000 3.4000 131.2000 ;
	    RECT 5.4000 130.8000 5.8000 131.2000 ;
	    RECT 11.0000 131.1000 11.4000 131.2000 ;
	    RECT 11.8000 131.1000 12.2000 131.2000 ;
	    RECT 11.0000 130.8000 12.2000 131.1000 ;
	    RECT 15.0000 130.8000 15.4000 131.2000 ;
	    RECT 3.0000 127.8000 3.3000 130.8000 ;
	    RECT 9.4000 129.8000 9.8000 130.2000 ;
	    RECT 9.4000 128.2000 9.7000 129.8000 ;
	    RECT 9.4000 127.8000 9.8000 128.2000 ;
	    RECT 15.0000 127.8000 15.3000 130.8000 ;
	    RECT 89.4000 130.2000 89.7000 134.8000 ;
	    RECT 108.0000 130.3000 109.6000 130.7000 ;
	    RECT 20.6000 129.8000 21.0000 130.2000 ;
	    RECT 27.8000 129.8000 28.2000 130.2000 ;
	    RECT 89.4000 129.8000 89.8000 130.2000 ;
	    RECT 20.6000 128.2000 20.9000 129.8000 ;
	    RECT 27.8000 128.2000 28.1000 129.8000 ;
	    RECT 147.8000 129.2000 148.1000 134.8000 ;
	    RECT 210.4000 130.3000 212.0000 130.7000 ;
	    RECT 147.8000 128.8000 148.2000 129.2000 ;
	    RECT 20.6000 127.8000 21.0000 128.2000 ;
	    RECT 27.8000 127.8000 28.2000 128.2000 ;
	    RECT 2.2000 127.5000 4.3000 127.8000 ;
	    RECT 2.2000 127.4000 2.6000 127.5000 ;
	    RECT 3.9000 127.4000 4.3000 127.5000 ;
	    RECT 15.0000 127.5000 17.1000 127.8000 ;
	    RECT 15.0000 127.4000 15.4000 127.5000 ;
	    RECT 16.7000 127.4000 17.1000 127.5000 ;
	    RECT 123.0000 114.8000 123.4000 115.2000 ;
	    RECT 13.3000 113.5000 13.7000 113.6000 ;
	    RECT 15.0000 113.5000 15.4000 113.6000 ;
	    RECT 13.3000 113.2000 15.4000 113.5000 ;
	    RECT 3.8000 112.8000 4.2000 113.2000 ;
	    RECT 7.8000 112.8000 8.2000 113.2000 ;
	    RECT 3.8000 111.2000 4.1000 112.8000 ;
	    RECT 7.8000 111.2000 8.1000 112.8000 ;
	    RECT 3.8000 110.8000 4.2000 111.2000 ;
	    RECT 4.6000 110.8000 5.0000 111.2000 ;
	    RECT 7.8000 110.8000 8.2000 111.2000 ;
	    RECT 12.6000 110.8000 13.0000 111.2000 ;
	    RECT 4.6000 110.2000 4.9000 110.8000 ;
	    RECT 4.6000 109.8000 5.0000 110.2000 ;
	    RECT 12.6000 108.1000 12.9000 110.8000 ;
	    RECT 15.0000 110.2000 15.3000 113.2000 ;
	    RECT 123.0000 113.1000 123.3000 114.8000 ;
	    RECT 122.2000 112.8000 123.3000 113.1000 ;
	    RECT 122.2000 112.7000 122.6000 112.8000 ;
	    RECT 108.0000 110.3000 109.6000 110.7000 ;
	    RECT 210.4000 110.3000 212.0000 110.7000 ;
	    RECT 15.0000 109.8000 15.4000 110.2000 ;
	    RECT 21.4000 109.8000 21.8000 110.2000 ;
	    RECT 21.4000 108.2000 21.7000 109.8000 ;
	    RECT 12.6000 107.8000 13.7000 108.1000 ;
	    RECT 21.4000 107.8000 21.8000 108.2000 ;
	    RECT 13.4000 107.2000 13.7000 107.8000 ;
	    RECT 13.4000 106.8000 13.8000 107.2000 ;
	    RECT 3.8000 106.1000 4.2000 106.2000 ;
	    RECT 3.8000 105.8000 4.9000 106.1000 ;
	    RECT 4.6000 95.2000 4.9000 105.8000 ;
	    RECT 3.0000 94.8000 3.4000 95.2000 ;
	    RECT 4.6000 94.8000 5.0000 95.2000 ;
	    RECT 3.0000 92.2000 3.3000 94.8000 ;
	    RECT 10.2000 93.8000 10.6000 94.2000 ;
	    RECT 17.4000 93.8000 17.8000 94.2000 ;
	    RECT 3.0000 91.8000 3.4000 92.2000 ;
	    RECT 10.2000 90.2000 10.5000 93.8000 ;
	    RECT 10.2000 89.8000 10.6000 90.2000 ;
	    RECT 10.2000 88.2000 10.5000 89.8000 ;
	    RECT 10.2000 87.8000 10.6000 88.2000 ;
	    RECT 10.2000 87.2000 10.5000 87.8000 ;
	    RECT 10.2000 86.8000 10.6000 87.2000 ;
	    RECT 17.4000 86.1000 17.7000 93.8000 ;
	    RECT 31.8000 92.8000 32.2000 93.2000 ;
	    RECT 31.8000 91.2000 32.1000 92.8000 ;
	    RECT 28.6000 90.8000 29.0000 91.2000 ;
	    RECT 31.8000 90.8000 32.2000 91.2000 ;
	    RECT 18.2000 88.8000 18.6000 89.2000 ;
	    RECT 18.2000 86.2000 18.5000 88.8000 ;
	    RECT 28.6000 87.8000 28.9000 90.8000 ;
	    RECT 108.0000 90.3000 109.6000 90.7000 ;
	    RECT 210.4000 90.3000 212.0000 90.7000 ;
	    RECT 36.6000 89.1000 37.0000 89.2000 ;
	    RECT 36.6000 88.8000 37.7000 89.1000 ;
	    RECT 28.5000 87.5000 30.6000 87.8000 ;
	    RECT 28.5000 87.4000 28.9000 87.5000 ;
	    RECT 30.2000 87.4000 30.6000 87.5000 ;
	    RECT 37.4000 87.2000 37.7000 88.8000 ;
	    RECT 26.2000 86.8000 26.6000 87.2000 ;
	    RECT 37.4000 86.8000 37.8000 87.2000 ;
	    RECT 26.2000 86.2000 26.5000 86.8000 ;
	    RECT 18.2000 86.1000 18.6000 86.2000 ;
	    RECT 17.4000 85.8000 18.6000 86.1000 ;
	    RECT 26.2000 85.8000 26.6000 86.2000 ;
	    RECT 7.0000 74.8000 7.4000 75.2000 ;
	    RECT 8.6000 74.8000 9.0000 75.2000 ;
	    RECT 5.4000 73.8000 5.8000 74.2000 ;
	    RECT 5.4000 72.2000 5.7000 73.8000 ;
	    RECT 5.4000 71.8000 5.8000 72.2000 ;
	    RECT 7.0000 70.2000 7.3000 74.8000 ;
	    RECT 8.6000 72.2000 8.9000 74.8000 ;
	    RECT 40.6000 73.8000 41.0000 74.2000 ;
	    RECT 11.8000 72.8000 12.2000 73.2000 ;
	    RECT 21.4000 72.8000 21.8000 73.2000 ;
	    RECT 8.6000 71.8000 9.0000 72.2000 ;
	    RECT 11.8000 71.2000 12.1000 72.8000 ;
	    RECT 21.4000 71.2000 21.7000 72.8000 ;
	    RECT 39.8000 72.1000 40.2000 72.2000 ;
	    RECT 40.6000 72.1000 40.9000 73.8000 ;
	    RECT 39.8000 71.8000 40.9000 72.1000 ;
	    RECT 11.8000 70.8000 12.2000 71.2000 ;
	    RECT 21.4000 70.8000 21.8000 71.2000 ;
	    RECT 108.0000 70.3000 109.6000 70.7000 ;
	    RECT 210.4000 70.3000 212.0000 70.7000 ;
	    RECT 6.2000 69.8000 6.6000 70.2000 ;
	    RECT 7.0000 69.8000 7.4000 70.2000 ;
	    RECT 2.2000 68.8000 2.6000 69.2000 ;
	    RECT 2.2000 67.2000 2.5000 68.8000 ;
	    RECT 6.2000 68.2000 6.5000 69.8000 ;
	    RECT 6.2000 67.8000 6.6000 68.2000 ;
	    RECT 200.6000 67.9000 201.0000 68.3000 ;
	    RECT 2.2000 66.8000 2.6000 67.2000 ;
	    RECT 200.6000 66.1000 200.9000 67.9000 ;
	    RECT 201.4000 66.1000 201.8000 66.2000 ;
	    RECT 200.6000 65.8000 201.8000 66.1000 ;
	    RECT 200.6000 55.2000 200.9000 65.8000 ;
	    RECT 152.6000 54.8000 153.0000 55.2000 ;
	    RECT 200.6000 54.8000 201.0000 55.2000 ;
	    RECT 5.4000 53.8000 5.8000 54.2000 ;
	    RECT 23.8000 53.8000 24.2000 54.2000 ;
	    RECT 4.6000 52.1000 5.0000 52.2000 ;
	    RECT 5.4000 52.1000 5.7000 53.8000 ;
	    RECT 4.6000 51.8000 5.7000 52.1000 ;
	    RECT 9.4000 52.8000 9.8000 53.2000 ;
	    RECT 16.6000 52.8000 17.0000 53.2000 ;
	    RECT 9.4000 51.2000 9.7000 52.8000 ;
	    RECT 16.6000 51.2000 16.9000 52.8000 ;
	    RECT 23.8000 52.2000 24.1000 53.8000 ;
	    RECT 42.2000 52.8000 42.6000 53.2000 ;
	    RECT 152.6000 53.1000 152.9000 54.8000 ;
	    RECT 151.8000 52.8000 152.9000 53.1000 ;
	    RECT 23.8000 51.8000 24.2000 52.2000 ;
	    RECT 42.2000 51.2000 42.5000 52.8000 ;
	    RECT 151.8000 52.7000 152.2000 52.8000 ;
	    RECT 7.8000 50.8000 8.2000 51.2000 ;
	    RECT 9.4000 50.8000 9.8000 51.2000 ;
	    RECT 16.6000 50.8000 17.0000 51.2000 ;
	    RECT 42.2000 50.8000 42.6000 51.2000 ;
	    RECT 1.4000 49.1000 1.8000 49.2000 ;
	    RECT 0.6000 48.8000 1.8000 49.1000 ;
	    RECT 0.6000 47.2000 0.9000 48.8000 ;
	    RECT 0.6000 46.8000 1.0000 47.2000 ;
	    RECT 7.8000 45.2000 8.1000 50.8000 ;
	    RECT 108.0000 50.3000 109.6000 50.7000 ;
	    RECT 210.4000 50.3000 212.0000 50.7000 ;
	    RECT 13.4000 48.8000 13.8000 49.2000 ;
	    RECT 22.2000 49.1000 22.6000 49.2000 ;
	    RECT 22.2000 48.8000 23.3000 49.1000 ;
	    RECT 13.4000 46.2000 13.7000 48.8000 ;
	    RECT 23.0000 47.2000 23.3000 48.8000 ;
	    RECT 39.0000 48.8000 39.4000 49.2000 ;
	    RECT 249.4000 48.8000 249.8000 49.2000 ;
	    RECT 259.0000 48.8000 259.4000 49.2000 ;
	    RECT 39.0000 47.2000 39.3000 48.8000 ;
	    RECT 23.0000 46.8000 23.4000 47.2000 ;
	    RECT 39.0000 46.8000 39.4000 47.2000 ;
	    RECT 249.4000 46.2000 249.7000 48.8000 ;
	    RECT 259.0000 46.2000 259.3000 48.8000 ;
	    RECT 13.4000 45.8000 13.8000 46.2000 ;
	    RECT 249.4000 45.8000 249.8000 46.2000 ;
	    RECT 251.0000 45.8000 251.4000 46.2000 ;
	    RECT 259.0000 45.8000 259.4000 46.2000 ;
	    RECT 251.0000 45.2000 251.3000 45.8000 ;
	    RECT 7.8000 44.8000 8.2000 45.2000 ;
	    RECT 251.0000 44.8000 251.4000 45.2000 ;
	    RECT 23.0000 34.8000 23.4000 35.2000 ;
	    RECT 235.0000 34.8000 235.4000 35.2000 ;
	    RECT 251.0000 34.8000 251.4000 35.2000 ;
	    RECT 5.4000 33.8000 5.8000 34.2000 ;
	    RECT 11.8000 33.8000 12.2000 34.2000 ;
	    RECT 3.8000 29.8000 4.2000 30.2000 ;
	    RECT 3.8000 28.2000 4.1000 29.8000 ;
	    RECT 4.6000 29.1000 5.0000 29.2000 ;
	    RECT 5.4000 29.1000 5.7000 33.8000 ;
	    RECT 4.6000 28.8000 5.7000 29.1000 ;
	    RECT 11.8000 33.2000 12.1000 33.8000 ;
	    RECT 11.8000 32.8000 12.2000 33.2000 ;
	    RECT 11.8000 31.2000 12.1000 32.8000 ;
	    RECT 23.0000 32.2000 23.3000 34.8000 ;
	    RECT 35.8000 33.8000 36.2000 34.2000 ;
	    RECT 23.0000 31.8000 23.4000 32.2000 ;
	    RECT 35.8000 32.1000 36.1000 33.8000 ;
	    RECT 235.0000 32.2000 235.3000 34.8000 ;
	    RECT 248.6000 33.8000 249.0000 34.2000 ;
	    RECT 241.4000 32.8000 241.8000 33.2000 ;
	    RECT 36.6000 32.1000 37.0000 32.2000 ;
	    RECT 35.8000 31.8000 37.0000 32.1000 ;
	    RECT 235.0000 31.8000 235.4000 32.2000 ;
	    RECT 241.4000 31.2000 241.7000 32.8000 ;
	    RECT 248.6000 32.2000 248.9000 33.8000 ;
	    RECT 249.4000 32.8000 249.8000 33.2000 ;
	    RECT 248.6000 31.8000 249.0000 32.2000 ;
	    RECT 249.4000 31.2000 249.7000 32.8000 ;
	    RECT 251.0000 32.2000 251.3000 34.8000 ;
	    RECT 251.0000 31.8000 251.4000 32.2000 ;
	    RECT 11.8000 30.8000 12.2000 31.2000 ;
	    RECT 15.8000 30.8000 16.2000 31.2000 ;
	    RECT 241.4000 30.8000 241.8000 31.2000 ;
	    RECT 249.4000 30.8000 249.8000 31.2000 ;
	    RECT 3.8000 27.8000 4.2000 28.2000 ;
	    RECT 4.6000 27.2000 4.9000 28.8000 ;
	    RECT 11.8000 28.2000 12.1000 30.8000 ;
	    RECT 11.8000 27.8000 12.2000 28.2000 ;
	    RECT 4.6000 26.8000 5.0000 27.2000 ;
	    RECT 15.8000 25.2000 16.1000 30.8000 ;
	    RECT 108.0000 30.3000 109.6000 30.7000 ;
	    RECT 210.4000 30.3000 212.0000 30.7000 ;
	    RECT 32.6000 29.8000 33.0000 30.2000 ;
	    RECT 223.8000 29.8000 224.2000 30.2000 ;
	    RECT 32.6000 28.2000 32.9000 29.8000 ;
	    RECT 220.6000 28.8000 221.0000 29.2000 ;
	    RECT 32.6000 27.8000 33.0000 28.2000 ;
	    RECT 220.6000 27.2000 220.9000 28.8000 ;
	    RECT 223.8000 28.2000 224.1000 29.8000 ;
	    RECT 223.8000 27.8000 224.2000 28.2000 ;
	    RECT 220.6000 26.8000 221.0000 27.2000 ;
	    RECT 15.8000 24.8000 16.2000 25.2000 ;
	    RECT 215.0000 17.8000 215.4000 18.2000 ;
	    RECT 218.2000 17.8000 218.6000 18.2000 ;
	    RECT 195.0000 15.8000 195.4000 16.2000 ;
	    RECT 27.8000 14.8000 28.2000 15.2000 ;
	    RECT 187.0000 14.8000 187.4000 15.2000 ;
	    RECT 27.8000 13.1000 28.1000 14.8000 ;
	    RECT 27.8000 12.8000 29.0000 13.1000 ;
	    RECT 28.6000 12.7000 29.0000 12.8000 ;
	    RECT 187.0000 12.2000 187.3000 14.8000 ;
	    RECT 190.2000 14.0000 190.6000 14.4000 ;
	    RECT 195.0000 14.2000 195.3000 15.8000 ;
	    RECT 215.0000 15.2000 215.3000 17.8000 ;
	    RECT 218.2000 17.2000 218.5000 17.8000 ;
	    RECT 218.2000 16.8000 218.6000 17.2000 ;
	    RECT 215.0000 14.8000 215.4000 15.2000 ;
	    RECT 259.8000 14.8000 260.2000 15.2000 ;
	    RECT 187.0000 11.8000 187.4000 12.2000 ;
	    RECT 190.2000 11.2000 190.5000 14.0000 ;
	    RECT 195.0000 13.8000 195.4000 14.2000 ;
	    RECT 196.6000 13.8000 197.0000 14.2000 ;
	    RECT 196.6000 13.2000 196.9000 13.8000 ;
	    RECT 196.6000 12.8000 197.0000 13.2000 ;
	    RECT 215.0000 12.2000 215.3000 14.8000 ;
	    RECT 249.4000 13.8000 249.8000 14.2000 ;
	    RECT 227.0000 12.8000 227.4000 13.2000 ;
	    RECT 215.0000 11.8000 215.4000 12.2000 ;
	    RECT 227.0000 11.2000 227.3000 12.8000 ;
	    RECT 249.4000 12.2000 249.7000 13.8000 ;
	    RECT 259.8000 12.2000 260.1000 14.8000 ;
	    RECT 249.4000 11.8000 249.8000 12.2000 ;
	    RECT 259.8000 11.8000 260.2000 12.2000 ;
	    RECT 187.8000 11.1000 188.2000 11.2000 ;
	    RECT 188.6000 11.1000 189.0000 11.2000 ;
	    RECT 187.8000 10.8000 189.0000 11.1000 ;
	    RECT 190.2000 10.8000 190.6000 11.2000 ;
	    RECT 227.0000 10.8000 227.4000 11.2000 ;
	    RECT 108.0000 10.3000 109.6000 10.7000 ;
	    RECT 210.4000 10.3000 212.0000 10.7000 ;
	    RECT 240.6000 9.8000 241.0000 10.2000 ;
	    RECT 258.2000 9.8000 258.6000 10.2000 ;
	    RECT 216.6000 8.8000 217.0000 9.2000 ;
	    RECT 216.6000 7.2000 216.9000 8.8000 ;
	    RECT 240.6000 8.2000 240.9000 9.8000 ;
	    RECT 258.2000 8.2000 258.5000 9.8000 ;
	    RECT 260.6000 8.8000 261.0000 9.2000 ;
	    RECT 240.6000 7.8000 241.0000 8.2000 ;
	    RECT 258.2000 7.8000 258.6000 8.2000 ;
	    RECT 260.6000 7.2000 260.9000 8.8000 ;
	    RECT 216.6000 6.8000 217.0000 7.2000 ;
	    RECT 260.6000 6.8000 261.0000 7.2000 ;
         LAYER metal3 ;
	    RECT 108.0000 170.3000 109.6000 170.7000 ;
	    RECT 210.4000 170.3000 212.0000 170.7000 ;
	    RECT 108.0000 150.3000 109.6000 150.7000 ;
	    RECT 210.4000 150.3000 212.0000 150.7000 ;
	    RECT 3.8000 147.1000 4.2000 147.2000 ;
	    RECT 10.2000 147.1000 10.6000 147.2000 ;
	    RECT 3.8000 146.8000 10.6000 147.1000 ;
	    RECT 12.6000 135.1000 13.0000 135.2000 ;
	    RECT 15.0000 135.1000 15.4000 135.2000 ;
	    RECT 12.6000 134.8000 15.4000 135.1000 ;
	    RECT 5.4000 131.1000 5.8000 131.2000 ;
	    RECT 11.8000 131.1000 12.2000 131.2000 ;
	    RECT 12.6000 131.1000 13.0000 131.2000 ;
	    RECT 5.4000 130.8000 13.0000 131.1000 ;
	    RECT 108.0000 130.3000 109.6000 130.7000 ;
	    RECT 210.4000 130.3000 212.0000 130.7000 ;
	    RECT 4.6000 110.8000 5.0000 111.2000 ;
	    RECT 4.6000 110.2000 4.9000 110.8000 ;
	    RECT 108.0000 110.3000 109.6000 110.7000 ;
	    RECT 210.4000 110.3000 212.0000 110.7000 ;
	    RECT 4.6000 109.8000 5.0000 110.2000 ;
	    RECT 3.8000 106.1000 4.2000 106.2000 ;
	    RECT 4.6000 106.1000 5.0000 106.2000 ;
	    RECT 3.8000 105.8000 5.0000 106.1000 ;
	    RECT 108.0000 90.3000 109.6000 90.7000 ;
	    RECT 210.4000 90.3000 212.0000 90.7000 ;
	    RECT 18.2000 86.1000 18.6000 86.2000 ;
	    RECT 26.2000 86.1000 26.6000 86.2000 ;
	    RECT 18.2000 85.8000 26.6000 86.1000 ;
	    RECT 108.0000 70.3000 109.6000 70.7000 ;
	    RECT 210.4000 70.3000 212.0000 70.7000 ;
	    RECT 108.0000 50.3000 109.6000 50.7000 ;
	    RECT 210.4000 50.3000 212.0000 50.7000 ;
	    RECT 251.0000 46.1000 251.4000 46.2000 ;
	    RECT 259.0000 46.1000 259.4000 46.2000 ;
	    RECT 251.0000 45.8000 259.4000 46.1000 ;
	    RECT 108.0000 30.3000 109.6000 30.7000 ;
	    RECT 210.4000 30.3000 212.0000 30.7000 ;
	    RECT 215.0000 18.1000 215.4000 18.2000 ;
	    RECT 218.2000 18.1000 218.6000 18.2000 ;
	    RECT 215.0000 17.8000 218.6000 18.1000 ;
	    RECT 195.0000 14.1000 195.4000 14.2000 ;
	    RECT 196.6000 14.1000 197.0000 14.2000 ;
	    RECT 195.0000 13.8000 197.0000 14.1000 ;
	    RECT 187.8000 11.1000 188.2000 11.2000 ;
	    RECT 190.2000 11.1000 190.6000 11.2000 ;
	    RECT 187.8000 10.8000 190.6000 11.1000 ;
	    RECT 108.0000 10.3000 109.6000 10.7000 ;
	    RECT 210.4000 10.3000 212.0000 10.7000 ;
         LAYER metal4 ;
	    RECT 108.0000 170.3000 109.6000 170.7000 ;
	    RECT 210.4000 170.3000 212.0000 170.7000 ;
	    RECT 108.0000 150.3000 109.6000 150.7000 ;
	    RECT 210.4000 150.3000 212.0000 150.7000 ;
	    RECT 12.6000 134.8000 13.0000 135.2000 ;
	    RECT 12.6000 131.2000 12.9000 134.8000 ;
	    RECT 12.6000 130.8000 13.0000 131.2000 ;
	    RECT 108.0000 130.3000 109.6000 130.7000 ;
	    RECT 210.4000 130.3000 212.0000 130.7000 ;
	    RECT 4.6000 110.8000 5.0000 111.2000 ;
	    RECT 4.6000 106.2000 4.9000 110.8000 ;
	    RECT 108.0000 110.3000 109.6000 110.7000 ;
	    RECT 210.4000 110.3000 212.0000 110.7000 ;
	    RECT 4.6000 105.8000 5.0000 106.2000 ;
	    RECT 108.0000 90.3000 109.6000 90.7000 ;
	    RECT 210.4000 90.3000 212.0000 90.7000 ;
	    RECT 108.0000 70.3000 109.6000 70.7000 ;
	    RECT 210.4000 70.3000 212.0000 70.7000 ;
	    RECT 108.0000 50.3000 109.6000 50.7000 ;
	    RECT 210.4000 50.3000 212.0000 50.7000 ;
	    RECT 108.0000 30.3000 109.6000 30.7000 ;
	    RECT 210.4000 30.3000 212.0000 30.7000 ;
	    RECT 108.0000 10.3000 109.6000 10.7000 ;
	    RECT 210.4000 10.3000 212.0000 10.7000 ;
         LAYER metal5 ;
	    RECT 108.0000 170.7000 108.6000 170.8000 ;
	    RECT 109.0000 170.7000 109.6000 170.8000 ;
	    RECT 108.0000 170.2000 109.6000 170.7000 ;
	    RECT 210.4000 170.7000 211.0000 170.8000 ;
	    RECT 211.4000 170.7000 212.0000 170.8000 ;
	    RECT 210.4000 170.2000 212.0000 170.7000 ;
	    RECT 108.0000 150.7000 108.6000 150.8000 ;
	    RECT 109.0000 150.7000 109.6000 150.8000 ;
	    RECT 108.0000 150.2000 109.6000 150.7000 ;
	    RECT 210.4000 150.7000 211.0000 150.8000 ;
	    RECT 211.4000 150.7000 212.0000 150.8000 ;
	    RECT 210.4000 150.2000 212.0000 150.7000 ;
	    RECT 108.0000 130.7000 108.6000 130.8000 ;
	    RECT 109.0000 130.7000 109.6000 130.8000 ;
	    RECT 108.0000 130.2000 109.6000 130.7000 ;
	    RECT 210.4000 130.7000 211.0000 130.8000 ;
	    RECT 211.4000 130.7000 212.0000 130.8000 ;
	    RECT 210.4000 130.2000 212.0000 130.7000 ;
	    RECT 108.0000 110.7000 108.6000 110.8000 ;
	    RECT 109.0000 110.7000 109.6000 110.8000 ;
	    RECT 108.0000 110.2000 109.6000 110.7000 ;
	    RECT 210.4000 110.7000 211.0000 110.8000 ;
	    RECT 211.4000 110.7000 212.0000 110.8000 ;
	    RECT 210.4000 110.2000 212.0000 110.7000 ;
	    RECT 108.0000 90.7000 108.6000 90.8000 ;
	    RECT 109.0000 90.7000 109.6000 90.8000 ;
	    RECT 108.0000 90.2000 109.6000 90.7000 ;
	    RECT 210.4000 90.7000 211.0000 90.8000 ;
	    RECT 211.4000 90.7000 212.0000 90.8000 ;
	    RECT 210.4000 90.2000 212.0000 90.7000 ;
	    RECT 108.0000 70.7000 108.6000 70.8000 ;
	    RECT 109.0000 70.7000 109.6000 70.8000 ;
	    RECT 108.0000 70.2000 109.6000 70.7000 ;
	    RECT 210.4000 70.7000 211.0000 70.8000 ;
	    RECT 211.4000 70.7000 212.0000 70.8000 ;
	    RECT 210.4000 70.2000 212.0000 70.7000 ;
	    RECT 108.0000 50.7000 108.6000 50.8000 ;
	    RECT 109.0000 50.7000 109.6000 50.8000 ;
	    RECT 108.0000 50.2000 109.6000 50.7000 ;
	    RECT 210.4000 50.7000 211.0000 50.8000 ;
	    RECT 211.4000 50.7000 212.0000 50.8000 ;
	    RECT 210.4000 50.2000 212.0000 50.7000 ;
	    RECT 108.0000 30.7000 108.6000 30.8000 ;
	    RECT 109.0000 30.7000 109.6000 30.8000 ;
	    RECT 108.0000 30.2000 109.6000 30.7000 ;
	    RECT 210.4000 30.7000 211.0000 30.8000 ;
	    RECT 211.4000 30.7000 212.0000 30.8000 ;
	    RECT 210.4000 30.2000 212.0000 30.7000 ;
	    RECT 108.0000 10.7000 108.6000 10.8000 ;
	    RECT 109.0000 10.7000 109.6000 10.8000 ;
	    RECT 108.0000 10.2000 109.6000 10.7000 ;
	    RECT 210.4000 10.7000 211.0000 10.8000 ;
	    RECT 211.4000 10.7000 212.0000 10.8000 ;
	    RECT 210.4000 10.2000 212.0000 10.7000 ;
         LAYER metal6 ;
	    RECT 108.0000 -3.0000 109.6000 183.0000 ;
	    RECT 210.4000 -3.0000 212.0000 183.0000 ;
      END
   END gnd
   PIN clk
      PORT
         LAYER metal1 ;
	    RECT 97.7000 134.1000 98.6000 134.5000 ;
	    RECT 98.2000 133.8000 98.6000 134.1000 ;
	    RECT 161.4000 134.1000 162.3000 134.5000 ;
	    RECT 168.6000 134.1000 169.5000 134.5000 ;
	    RECT 161.4000 133.8000 161.8000 134.1000 ;
	    RECT 168.6000 133.8000 169.0000 134.1000 ;
	    RECT 84.6000 126.9000 85.0000 127.2000 ;
	    RECT 84.6000 126.5000 85.5000 126.9000 ;
	    RECT 147.0000 94.1000 147.9000 94.5000 ;
	    RECT 147.0000 93.8000 147.4000 94.1000 ;
	    RECT 150.5000 74.1000 151.4000 74.5000 ;
	    RECT 157.7000 74.1000 158.6000 74.5000 ;
	    RECT 151.0000 73.8000 151.4000 74.1000 ;
	    RECT 158.2000 73.8000 158.6000 74.1000 ;
	    RECT 140.6000 46.9000 141.0000 47.2000 ;
	    RECT 140.1000 46.5000 141.0000 46.9000 ;
	    RECT 140.6000 46.2000 140.9000 46.5000 ;
	    RECT 140.6000 45.8000 141.0000 46.2000 ;
	    RECT 182.2000 26.9000 182.6000 27.2000 ;
	    RECT 182.2000 26.5000 183.1000 26.9000 ;
	    RECT 83.3000 14.1000 84.2000 14.5000 ;
	    RECT 83.8000 13.8000 84.2000 14.1000 ;
	    RECT 147.8000 14.1000 148.7000 14.5000 ;
	    RECT 163.8000 14.1000 164.7000 14.5000 ;
	    RECT 147.8000 13.8000 148.2000 14.1000 ;
	    RECT 163.8000 13.8000 164.2000 14.1000 ;
         LAYER metal2 ;
	    RECT 84.6000 133.8000 85.0000 134.2000 ;
	    RECT 98.2000 134.1000 98.6000 134.2000 ;
	    RECT 99.0000 134.1000 99.4000 134.2000 ;
	    RECT 98.2000 133.8000 99.4000 134.1000 ;
	    RECT 161.4000 133.8000 161.8000 134.2000 ;
	    RECT 167.8000 134.1000 168.2000 134.2000 ;
	    RECT 168.6000 134.1000 169.0000 134.2000 ;
	    RECT 167.8000 133.8000 169.0000 134.1000 ;
	    RECT 84.6000 127.2000 84.9000 133.8000 ;
	    RECT 161.4000 129.2000 161.7000 133.8000 ;
	    RECT 161.4000 128.8000 161.8000 129.2000 ;
	    RECT 84.6000 126.8000 85.0000 127.2000 ;
	    RECT 147.0000 106.8000 147.4000 107.2000 ;
	    RECT 147.0000 94.2000 147.3000 106.8000 ;
	    RECT 147.0000 93.8000 147.4000 94.2000 ;
	    RECT 147.0000 74.2000 147.3000 93.8000 ;
	    RECT 147.0000 73.8000 147.4000 74.2000 ;
	    RECT 151.0000 74.1000 151.4000 74.2000 ;
	    RECT 150.2000 73.8000 151.4000 74.1000 ;
	    RECT 157.4000 74.1000 157.8000 74.2000 ;
	    RECT 158.2000 74.1000 158.6000 74.2000 ;
	    RECT 157.4000 73.8000 158.6000 74.1000 ;
	    RECT 150.2000 47.2000 150.5000 73.8000 ;
	    RECT 140.6000 46.8000 141.0000 47.2000 ;
	    RECT 150.2000 46.8000 150.6000 47.2000 ;
	    RECT 140.6000 46.2000 140.9000 46.8000 ;
	    RECT 140.6000 45.8000 141.0000 46.2000 ;
	    RECT 182.2000 26.8000 182.6000 27.2000 ;
	    RECT 182.2000 26.2000 182.5000 26.8000 ;
	    RECT 163.8000 25.8000 164.2000 26.2000 ;
	    RECT 182.2000 25.8000 182.6000 26.2000 ;
	    RECT 83.8000 16.8000 84.2000 17.2000 ;
	    RECT 83.8000 14.2000 84.1000 16.8000 ;
	    RECT 163.8000 14.2000 164.1000 25.8000 ;
	    RECT 83.8000 13.8000 84.2000 14.2000 ;
	    RECT 147.8000 14.1000 148.2000 14.2000 ;
	    RECT 148.6000 14.1000 149.0000 14.2000 ;
	    RECT 147.8000 13.8000 149.0000 14.1000 ;
	    RECT 163.0000 14.1000 163.4000 14.2000 ;
	    RECT 163.8000 14.1000 164.2000 14.2000 ;
	    RECT 163.0000 13.8000 164.2000 14.1000 ;
	    RECT 83.8000 0.8000 84.2000 1.2000 ;
	    RECT 83.8000 -1.8000 84.1000 0.8000 ;
	    RECT 83.8000 -2.2000 84.2000 -1.8000 ;
         LAYER metal3 ;
	    RECT 84.6000 134.1000 85.0000 134.2000 ;
	    RECT 99.0000 134.1000 99.4000 134.2000 ;
	    RECT 161.4000 134.1000 161.8000 134.2000 ;
	    RECT 167.8000 134.1000 168.2000 134.2000 ;
	    RECT 84.6000 133.8000 168.2000 134.1000 ;
	    RECT 159.0000 129.1000 159.4000 129.2000 ;
	    RECT 161.4000 129.1000 161.8000 129.2000 ;
	    RECT 159.0000 128.8000 161.8000 129.1000 ;
	    RECT 147.0000 107.1000 147.4000 107.2000 ;
	    RECT 159.0000 107.1000 159.4000 107.2000 ;
	    RECT 147.0000 106.8000 159.4000 107.1000 ;
	    RECT 147.0000 74.1000 147.4000 74.2000 ;
	    RECT 151.0000 74.1000 151.4000 74.2000 ;
	    RECT 157.4000 74.1000 157.8000 74.2000 ;
	    RECT 147.0000 73.8000 157.8000 74.1000 ;
	    RECT 140.6000 47.1000 141.0000 47.2000 ;
	    RECT 147.8000 47.1000 148.2000 47.2000 ;
	    RECT 150.2000 47.1000 150.6000 47.2000 ;
	    RECT 140.6000 46.8000 150.6000 47.1000 ;
	    RECT 163.8000 26.1000 164.2000 26.2000 ;
	    RECT 182.2000 26.1000 182.6000 26.2000 ;
	    RECT 163.8000 25.8000 182.6000 26.1000 ;
	    RECT 83.8000 17.1000 84.2000 17.2000 ;
	    RECT 147.8000 17.1000 148.2000 17.2000 ;
	    RECT 83.8000 16.8000 148.2000 17.1000 ;
	    RECT 147.8000 14.1000 148.2000 14.2000 ;
	    RECT 148.6000 14.1000 149.0000 14.2000 ;
	    RECT 163.0000 14.1000 163.4000 14.2000 ;
	    RECT 147.8000 13.8000 163.4000 14.1000 ;
	    RECT 83.8000 1.8000 84.2000 2.2000 ;
	    RECT 83.8000 1.2000 84.1000 1.8000 ;
	    RECT 83.8000 0.8000 84.2000 1.2000 ;
         LAYER metal4 ;
	    RECT 159.0000 128.8000 159.4000 129.2000 ;
	    RECT 159.0000 107.2000 159.3000 128.8000 ;
	    RECT 159.0000 106.8000 159.4000 107.2000 ;
	    RECT 147.8000 46.8000 148.2000 47.2000 ;
	    RECT 147.8000 17.2000 148.1000 46.8000 ;
	    RECT 83.8000 16.8000 84.2000 17.2000 ;
	    RECT 147.8000 16.8000 148.2000 17.2000 ;
	    RECT 83.8000 2.2000 84.1000 16.8000 ;
	    RECT 147.8000 14.2000 148.1000 16.8000 ;
	    RECT 147.8000 13.8000 148.2000 14.2000 ;
	    RECT 83.8000 1.8000 84.2000 2.2000 ;
      END
   END clk
   PIN reset
      PORT
         LAYER metal1 ;
	    RECT 74.1000 154.8000 74.6000 155.2000 ;
	    RECT 74.1000 154.4000 74.5000 154.8000 ;
	    RECT 74.1000 134.8000 74.6000 135.2000 ;
	    RECT 74.1000 134.4000 74.5000 134.8000 ;
	    RECT 162.3000 126.2000 162.7000 126.6000 ;
	    RECT 159.8000 126.1000 160.2000 126.2000 ;
	    RECT 162.2000 126.1000 162.7000 126.2000 ;
	    RECT 159.8000 125.8000 162.7000 126.1000 ;
	    RECT 158.1000 115.1000 158.6000 115.2000 ;
	    RECT 159.0000 115.1000 159.4000 115.2000 ;
	    RECT 158.1000 114.8000 159.4000 115.1000 ;
	    RECT 158.1000 114.4000 158.5000 114.8000 ;
	    RECT 169.3000 66.2000 169.7000 66.6000 ;
	    RECT 170.3000 66.2000 170.7000 66.6000 ;
	    RECT 169.3000 66.1000 169.8000 66.2000 ;
	    RECT 170.2000 66.1000 170.7000 66.2000 ;
	    RECT 169.3000 65.8000 170.7000 66.1000 ;
         LAYER metal2 ;
	    RECT 74.2000 182.8000 74.6000 183.2000 ;
	    RECT 74.2000 180.2000 74.5000 182.8000 ;
	    RECT 74.2000 179.8000 74.6000 180.2000 ;
	    RECT 74.2000 154.8000 74.6000 155.2000 ;
	    RECT 74.2000 154.2000 74.5000 154.8000 ;
	    RECT 74.2000 153.8000 74.6000 154.2000 ;
	    RECT 75.0000 140.1000 75.4000 140.2000 ;
	    RECT 74.2000 139.8000 75.4000 140.1000 ;
	    RECT 74.2000 135.2000 74.5000 139.8000 ;
	    RECT 74.2000 134.8000 74.6000 135.2000 ;
	    RECT 74.2000 119.2000 74.5000 134.8000 ;
	    RECT 159.8000 126.1000 160.2000 126.2000 ;
	    RECT 159.0000 125.8000 160.2000 126.1000 ;
	    RECT 159.0000 119.2000 159.3000 125.8000 ;
	    RECT 74.2000 118.8000 74.6000 119.2000 ;
	    RECT 159.0000 118.8000 159.4000 119.2000 ;
	    RECT 159.0000 115.2000 159.3000 118.8000 ;
	    RECT 159.0000 114.8000 159.4000 115.2000 ;
	    RECT 159.0000 96.2000 159.3000 114.8000 ;
	    RECT 159.0000 95.8000 159.4000 96.2000 ;
	    RECT 169.4000 70.8000 169.8000 71.2000 ;
	    RECT 169.4000 66.2000 169.7000 70.8000 ;
	    RECT 169.4000 65.8000 169.8000 66.2000 ;
         LAYER metal3 ;
	    RECT 74.2000 179.8000 74.6000 180.2000 ;
	    RECT 74.2000 179.2000 74.5000 179.8000 ;
	    RECT 74.2000 178.8000 74.6000 179.2000 ;
	    RECT 74.2000 154.8000 74.6000 155.2000 ;
	    RECT 74.2000 154.2000 74.5000 154.8000 ;
	    RECT 74.2000 153.8000 74.6000 154.2000 ;
	    RECT 74.2000 140.1000 74.6000 140.2000 ;
	    RECT 75.0000 140.1000 75.4000 140.2000 ;
	    RECT 74.2000 139.8000 75.4000 140.1000 ;
	    RECT 74.2000 119.1000 74.6000 119.2000 ;
	    RECT 159.0000 119.1000 159.4000 119.2000 ;
	    RECT 74.2000 118.8000 159.4000 119.1000 ;
	    RECT 159.0000 96.1000 159.4000 96.2000 ;
	    RECT 162.2000 96.1000 162.6000 96.2000 ;
	    RECT 159.0000 95.8000 162.6000 96.1000 ;
	    RECT 162.2000 71.1000 162.6000 71.2000 ;
	    RECT 169.4000 71.1000 169.8000 71.2000 ;
	    RECT 162.2000 70.8000 169.8000 71.1000 ;
         LAYER metal4 ;
	    RECT 74.2000 178.8000 74.6000 179.2000 ;
	    RECT 74.2000 155.2000 74.5000 178.8000 ;
	    RECT 74.2000 154.8000 74.6000 155.2000 ;
	    RECT 74.2000 140.2000 74.5000 154.8000 ;
	    RECT 74.2000 139.8000 74.6000 140.2000 ;
	    RECT 162.2000 95.8000 162.6000 96.2000 ;
	    RECT 162.2000 71.2000 162.5000 95.8000 ;
	    RECT 162.2000 70.8000 162.6000 71.2000 ;
      END
   END reset
   PIN block0[0]
      PORT
         LAYER metal1 ;
	    RECT 256.6000 73.4000 257.0000 74.2000 ;
	    RECT 256.6000 67.8000 257.0000 68.6000 ;
         LAYER metal2 ;
	    RECT 256.6000 73.8000 257.0000 74.2000 ;
	    RECT 256.6000 69.2000 256.9000 73.8000 ;
	    RECT 256.6000 68.8000 257.0000 69.2000 ;
	    RECT 256.6000 68.2000 256.9000 68.8000 ;
	    RECT 256.6000 67.8000 257.0000 68.2000 ;
         LAYER metal3 ;
	    RECT 256.6000 69.1000 257.0000 69.2000 ;
	    RECT 256.6000 68.8000 273.7000 69.1000 ;
	    RECT 273.4000 68.2000 273.7000 68.8000 ;
	    RECT 273.4000 67.8000 273.8000 68.2000 ;
      END
   END block0[0]
   PIN block0[1]
      PORT
         LAYER metal2 ;
	    RECT 25.4000 182.8000 25.8000 183.2000 ;
      END
   END block0[1]
   PIN block0[2]
      PORT
         LAYER metal2 ;
	    RECT 59.8000 -2.2000 60.2000 -1.8000 ;
      END
   END block0[2]
   PIN block0[3]
      PORT
         LAYER metal3 ;
	    RECT 273.4000 172.8000 273.8000 173.2000 ;
      END
   END block0[3]
   PIN block0[4]
      PORT
         LAYER metal3 ;
	    RECT 273.4000 124.8000 273.8000 125.2000 ;
      END
   END block0[4]
   PIN block0[5]
      PORT
         LAYER metal3 ;
	    RECT 273.4000 86.8000 273.8000 87.2000 ;
      END
   END block0[5]
   PIN block0[6]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 167.8000 -2.2000 168.2000 ;
      END
   END block0[6]
   PIN block0[7]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 52.8000 -2.2000 53.2000 ;
      END
   END block0[7]
   PIN block1[0]
      PORT
         LAYER metal1 ;
	    RECT 269.4000 93.1000 269.8000 93.2000 ;
	    RECT 270.2000 93.1000 270.6000 93.2000 ;
	    RECT 269.4000 92.8000 270.6000 93.1000 ;
	    RECT 269.4000 92.4000 269.8000 92.8000 ;
	    RECT 270.2000 47.8000 270.6000 48.2000 ;
	    RECT 269.4000 47.1000 269.8000 47.6000 ;
	    RECT 270.2000 47.1000 270.5000 47.8000 ;
	    RECT 269.4000 46.8000 270.5000 47.1000 ;
         LAYER metal2 ;
	    RECT 270.2000 92.8000 270.6000 93.2000 ;
	    RECT 270.2000 48.2000 270.5000 92.8000 ;
	    RECT 270.2000 47.8000 270.6000 48.2000 ;
	    RECT 270.2000 47.2000 270.5000 47.8000 ;
	    RECT 270.2000 46.8000 270.6000 47.2000 ;
         LAYER metal3 ;
	    RECT 270.2000 47.1000 270.6000 47.2000 ;
	    RECT 273.4000 47.1000 273.8000 47.2000 ;
	    RECT 270.2000 46.8000 273.8000 47.1000 ;
      END
   END block1[0]
   PIN block1[1]
      PORT
         LAYER metal2 ;
	    RECT 251.8000 -2.2000 252.2000 -1.8000 ;
      END
   END block1[1]
   PIN block1[2]
      PORT
         LAYER metal2 ;
	    RECT 238.2000 182.8000 238.6000 183.2000 ;
      END
   END block1[2]
   PIN block1[3]
      PORT
         LAYER metal3 ;
	    RECT 273.4000 97.8000 273.8000 98.2000 ;
      END
   END block1[3]
   PIN block1[4]
      PORT
         LAYER metal2 ;
	    RECT 156.6000 -2.2000 157.0000 -1.8000 ;
      END
   END block1[4]
   PIN block1[5]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 71.8000 -2.2000 72.2000 ;
      END
   END block1[5]
   PIN block1[6]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 150.8000 -2.2000 151.2000 ;
      END
   END block1[6]
   PIN block1[7]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 46.8000 -2.2000 47.2000 ;
      END
   END block1[7]
   PIN block2[0]
      PORT
         LAYER metal1 ;
	    RECT 261.8000 66.8000 262.6000 67.2000 ;
	    RECT 262.6000 56.8000 263.0000 57.2000 ;
	    RECT 262.7000 56.2000 263.0000 56.8000 ;
	    RECT 262.7000 55.9000 263.4000 56.2000 ;
	    RECT 263.0000 55.8000 263.4000 55.9000 ;
	    RECT 263.8000 52.4000 264.2000 53.2000 ;
         LAYER metal2 ;
	    RECT 262.2000 66.8000 262.6000 67.2000 ;
	    RECT 262.2000 59.2000 262.5000 66.8000 ;
	    RECT 262.2000 58.8000 262.6000 59.2000 ;
	    RECT 262.2000 56.1000 262.5000 58.8000 ;
	    RECT 263.0000 56.1000 263.4000 56.2000 ;
	    RECT 262.2000 55.8000 264.1000 56.1000 ;
	    RECT 263.8000 53.2000 264.1000 55.8000 ;
	    RECT 263.8000 52.8000 264.2000 53.2000 ;
         LAYER metal3 ;
	    RECT 262.2000 59.1000 262.6000 59.2000 ;
	    RECT 273.4000 59.1000 273.8000 59.2000 ;
	    RECT 262.2000 58.8000 273.8000 59.1000 ;
      END
   END block2[0]
   PIN block2[1]
      PORT
         LAYER metal2 ;
	    RECT 4.6000 -2.2000 5.0000 -1.8000 ;
      END
   END block2[1]
   PIN block2[2]
      PORT
         LAYER metal2 ;
	    RECT 218.2000 -2.2000 218.6000 -1.8000 ;
      END
   END block2[2]
   PIN block2[3]
      PORT
         LAYER metal2 ;
	    RECT 75.8000 -2.2000 76.2000 -1.8000 ;
      END
   END block2[3]
   PIN block2[4]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 81.8000 -2.2000 82.2000 ;
      END
   END block2[4]
   PIN block2[5]
      PORT
         LAYER metal2 ;
	    RECT 176.6000 182.8000 177.0000 183.2000 ;
      END
   END block2[5]
   PIN block2[6]
      PORT
         LAYER metal3 ;
	    RECT 273.4000 166.8000 273.8000 167.2000 ;
      END
   END block2[6]
   PIN block2[7]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 2.8000 -2.2000 3.2000 ;
      END
   END block2[7]
   PIN block3[0]
      PORT
         LAYER metal1 ;
	    RECT 250.6000 73.8000 251.4000 74.2000 ;
	    RECT 266.2000 73.4000 266.6000 74.2000 ;
	    RECT 263.8000 72.4000 264.2000 73.2000 ;
         LAYER metal2 ;
	    RECT 263.8000 74.8000 264.2000 75.2000 ;
	    RECT 266.2000 74.8000 266.6000 75.2000 ;
	    RECT 263.8000 74.2000 264.1000 74.8000 ;
	    RECT 266.2000 74.2000 266.5000 74.8000 ;
	    RECT 251.0000 74.1000 251.4000 74.2000 ;
	    RECT 251.8000 74.1000 252.2000 74.2000 ;
	    RECT 251.0000 73.8000 252.2000 74.1000 ;
	    RECT 263.8000 73.8000 264.2000 74.2000 ;
	    RECT 266.2000 73.8000 266.6000 74.2000 ;
	    RECT 263.8000 73.2000 264.1000 73.8000 ;
	    RECT 263.8000 72.8000 264.2000 73.2000 ;
         LAYER metal3 ;
	    RECT 263.8000 75.1000 264.2000 75.2000 ;
	    RECT 266.2000 75.1000 266.6000 75.2000 ;
	    RECT 273.4000 75.1000 273.8000 75.2000 ;
	    RECT 263.8000 74.8000 273.8000 75.1000 ;
	    RECT 251.8000 74.1000 252.2000 74.2000 ;
	    RECT 263.8000 74.1000 264.2000 74.2000 ;
	    RECT 251.8000 73.8000 264.2000 74.1000 ;
      END
   END block3[0]
   PIN block3[1]
      PORT
         LAYER metal2 ;
	    RECT 172.6000 182.8000 173.0000 183.2000 ;
      END
   END block3[1]
   PIN block3[2]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 98.8000 -2.2000 99.2000 ;
      END
   END block3[2]
   PIN block3[3]
      PORT
         LAYER metal3 ;
	    RECT 273.4000 7.8000 273.8000 8.2000 ;
      END
   END block3[3]
   PIN block3[4]
      PORT
         LAYER metal2 ;
	    RECT 195.8000 182.8000 196.2000 183.2000 ;
      END
   END block3[4]
   PIN block3[5]
      PORT
         LAYER metal2 ;
	    RECT 73.4000 -2.2000 73.8000 -1.8000 ;
      END
   END block3[5]
   PIN block3[6]
      PORT
         LAYER metal2 ;
	    RECT 183.0000 182.8000 183.4000 183.2000 ;
      END
   END block3[6]
   PIN block3[7]
      PORT
         LAYER metal3 ;
	    RECT 273.4000 91.8000 273.8000 92.2000 ;
      END
   END block3[7]
   PIN block4[0]
      PORT
         LAYER metal1 ;
	    RECT 262.2000 94.8000 262.6000 95.2000 ;
	    RECT 262.2000 94.2000 262.5000 94.8000 ;
	    RECT 261.0000 94.1000 261.8000 94.2000 ;
	    RECT 262.2000 94.1000 263.0000 94.2000 ;
	    RECT 261.0000 93.8000 263.0000 94.1000 ;
         LAYER metal2 ;
	    RECT 262.2000 94.8000 262.6000 95.2000 ;
	    RECT 262.2000 94.2000 262.5000 94.8000 ;
	    RECT 262.2000 93.8000 262.6000 94.2000 ;
         LAYER metal3 ;
	    RECT 262.2000 94.1000 262.6000 94.2000 ;
	    RECT 273.4000 94.1000 273.8000 94.2000 ;
	    RECT 262.2000 93.8000 273.8000 94.1000 ;
      END
   END block4[0]
   PIN block4[1]
      PORT
         LAYER metal2 ;
	    RECT 82.2000 182.8000 82.6000 183.2000 ;
      END
   END block4[1]
   PIN block4[2]
      PORT
         LAYER metal2 ;
	    RECT 148.6000 -2.2000 149.0000 -1.8000 ;
      END
   END block4[2]
   PIN block4[3]
      PORT
         LAYER metal2 ;
	    RECT 10.2000 182.8000 10.6000 183.2000 ;
      END
   END block4[3]
   PIN block4[4]
      PORT
         LAYER metal3 ;
	    RECT 273.4000 110.8000 273.8000 111.2000 ;
      END
   END block4[4]
   PIN block4[5]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 12.8000 -2.2000 13.2000 ;
      END
   END block4[5]
   PIN block4[6]
      PORT
         LAYER metal3 ;
	    RECT 273.4000 61.8000 273.8000 62.2000 ;
      END
   END block4[6]
   PIN block4[7]
      PORT
         LAYER metal3 ;
	    RECT 273.4000 49.8000 273.8000 50.2000 ;
      END
   END block4[7]
   PIN block5[0]
      PORT
         LAYER metal1 ;
	    RECT 262.6000 87.1000 263.4000 87.2000 ;
	    RECT 263.8000 87.1000 264.6000 87.2000 ;
	    RECT 262.6000 86.8000 264.6000 87.1000 ;
         LAYER metal2 ;
	    RECT 263.8000 88.8000 264.2000 89.2000 ;
	    RECT 263.8000 87.2000 264.1000 88.8000 ;
	    RECT 263.8000 86.8000 264.2000 87.2000 ;
         LAYER metal3 ;
	    RECT 263.8000 89.1000 264.2000 89.2000 ;
	    RECT 273.4000 89.1000 273.8000 89.2000 ;
	    RECT 263.8000 88.8000 273.8000 89.1000 ;
      END
   END block5[0]
   PIN block5[1]
      PORT
         LAYER metal3 ;
	    RECT 273.4000 56.8000 273.8000 57.2000 ;
      END
   END block5[1]
   PIN block5[2]
      PORT
         LAYER metal2 ;
	    RECT 53.4000 -2.2000 53.8000 -1.8000 ;
      END
   END block5[2]
   PIN block5[3]
      PORT
         LAYER metal2 ;
	    RECT 29.4000 182.8000 29.8000 183.2000 ;
      END
   END block5[3]
   PIN block5[4]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 165.8000 -2.2000 166.2000 ;
      END
   END block5[4]
   PIN block5[5]
      PORT
         LAYER metal2 ;
	    RECT 233.4000 -2.2000 233.8000 -1.8000 ;
      END
   END block5[5]
   PIN block5[6]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 128.8000 -2.2000 129.2000 ;
      END
   END block5[6]
   PIN block5[7]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 29.8000 -2.2000 30.2000 ;
      END
   END block5[7]
   PIN block6[0]
      PORT
         LAYER metal1 ;
	    RECT 268.6000 114.1000 269.0000 114.2000 ;
	    RECT 270.2000 114.1000 270.6000 114.2000 ;
	    RECT 268.6000 113.8000 270.6000 114.1000 ;
	    RECT 268.6000 113.4000 269.0000 113.8000 ;
	    RECT 263.4000 107.2000 263.8000 107.4000 ;
	    RECT 260.2000 106.8000 261.0000 107.2000 ;
	    RECT 263.4000 106.9000 264.2000 107.2000 ;
	    RECT 263.8000 106.8000 264.2000 106.9000 ;
         LAYER metal2 ;
	    RECT 270.2000 114.8000 270.6000 115.2000 ;
	    RECT 270.2000 114.2000 270.5000 114.8000 ;
	    RECT 270.2000 113.8000 270.6000 114.2000 ;
	    RECT 270.2000 108.2000 270.5000 113.8000 ;
	    RECT 260.6000 107.8000 261.0000 108.2000 ;
	    RECT 263.8000 107.8000 264.2000 108.2000 ;
	    RECT 270.2000 107.8000 270.6000 108.2000 ;
	    RECT 260.6000 107.2000 260.9000 107.8000 ;
	    RECT 263.8000 107.2000 264.1000 107.8000 ;
	    RECT 260.6000 106.8000 261.0000 107.2000 ;
	    RECT 263.8000 106.8000 264.2000 107.2000 ;
         LAYER metal3 ;
	    RECT 270.2000 115.1000 270.6000 115.2000 ;
	    RECT 273.4000 115.1000 273.8000 115.2000 ;
	    RECT 270.2000 114.8000 273.8000 115.1000 ;
	    RECT 260.6000 108.1000 261.0000 108.2000 ;
	    RECT 263.8000 108.1000 264.2000 108.2000 ;
	    RECT 270.2000 108.1000 270.6000 108.2000 ;
	    RECT 260.6000 107.8000 270.6000 108.1000 ;
      END
   END block6[0]
   PIN block6[1]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 77.8000 -2.2000 78.2000 ;
      END
   END block6[1]
   PIN block6[2]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 145.8000 -2.2000 146.2000 ;
      END
   END block6[2]
   PIN block6[3]
      PORT
         LAYER metal2 ;
	    RECT 135.0000 182.8000 135.4000 183.2000 ;
      END
   END block6[3]
   PIN block6[4]
      PORT
         LAYER metal3 ;
	    RECT 273.4000 106.8000 273.8000 107.2000 ;
      END
   END block6[4]
   PIN block6[5]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 16.8000 -2.2000 17.2000 ;
      END
   END block6[5]
   PIN block6[6]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 90.8000 -2.2000 91.2000 ;
      END
   END block6[6]
   PIN block6[7]
      PORT
         LAYER metal2 ;
	    RECT 194.2000 182.8000 194.6000 183.2000 ;
      END
   END block6[7]
   PIN block7[0]
      PORT
         LAYER metal1 ;
	    RECT 255.0000 172.4000 255.4000 173.2000 ;
	    RECT 259.8000 112.4000 260.2000 113.2000 ;
	    RECT 245.8000 106.8000 246.6000 107.2000 ;
	    RECT 261.4000 54.4000 261.8000 55.2000 ;
	    RECT 269.4000 54.8000 269.8000 55.6000 ;
         LAYER metal2 ;
	    RECT 255.0000 173.1000 255.4000 173.2000 ;
	    RECT 255.8000 173.1000 256.2000 173.2000 ;
	    RECT 255.0000 172.8000 256.2000 173.1000 ;
	    RECT 259.8000 112.8000 260.2000 113.2000 ;
	    RECT 259.8000 111.2000 260.1000 112.8000 ;
	    RECT 246.2000 110.8000 246.6000 111.2000 ;
	    RECT 259.8000 110.8000 260.2000 111.2000 ;
	    RECT 246.2000 107.2000 246.5000 110.8000 ;
	    RECT 246.2000 106.8000 246.6000 107.2000 ;
	    RECT 269.4000 55.8000 269.8000 56.2000 ;
	    RECT 269.4000 55.2000 269.7000 55.8000 ;
	    RECT 261.4000 55.1000 261.8000 55.2000 ;
	    RECT 262.2000 55.1000 262.6000 55.2000 ;
	    RECT 261.4000 54.8000 262.6000 55.1000 ;
	    RECT 269.4000 54.8000 269.8000 55.2000 ;
         LAYER metal3 ;
	    RECT 253.4000 173.1000 253.8000 173.2000 ;
	    RECT 255.8000 173.1000 256.2000 173.2000 ;
	    RECT 253.4000 172.8000 256.2000 173.1000 ;
	    RECT 246.2000 111.1000 246.6000 111.2000 ;
	    RECT 253.4000 111.1000 253.8000 111.2000 ;
	    RECT 259.8000 111.1000 260.2000 111.2000 ;
	    RECT 261.4000 111.1000 261.8000 111.2000 ;
	    RECT 246.2000 110.8000 261.8000 111.1000 ;
	    RECT 269.4000 55.8000 269.8000 56.2000 ;
	    RECT 261.4000 55.1000 261.8000 55.2000 ;
	    RECT 262.2000 55.1000 262.6000 55.2000 ;
	    RECT 269.4000 55.1000 269.7000 55.8000 ;
	    RECT 273.4000 55.1000 273.8000 55.2000 ;
	    RECT 261.4000 54.8000 273.8000 55.1000 ;
         LAYER metal4 ;
	    RECT 253.4000 172.8000 253.8000 173.2000 ;
	    RECT 253.4000 111.2000 253.7000 172.8000 ;
	    RECT 253.4000 110.8000 253.8000 111.2000 ;
	    RECT 261.4000 110.8000 261.8000 111.2000 ;
	    RECT 261.4000 55.2000 261.7000 110.8000 ;
	    RECT 261.4000 54.8000 261.8000 55.2000 ;
      END
   END block7[0]
   PIN block7[1]
      PORT
         LAYER metal3 ;
	    RECT 273.4000 26.8000 273.8000 27.2000 ;
      END
   END block7[1]
   PIN block7[2]
      PORT
         LAYER metal2 ;
	    RECT 7.8000 182.8000 8.2000 183.2000 ;
      END
   END block7[2]
   PIN block7[3]
      PORT
         LAYER metal3 ;
	    RECT 273.4000 112.8000 273.8000 113.2000 ;
      END
   END block7[3]
   PIN block7[4]
      PORT
         LAYER metal3 ;
	    RECT 273.4000 133.8000 273.8000 134.2000 ;
      END
   END block7[4]
   PIN block7[5]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 64.8000 -2.2000 65.2000 ;
      END
   END block7[5]
   PIN block7[6]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 92.8000 -2.2000 93.2000 ;
      END
   END block7[6]
   PIN block7[7]
      PORT
         LAYER metal3 ;
	    RECT 273.4000 24.8000 273.8000 25.2000 ;
      END
   END block7[7]
   PIN block8[0]
      PORT
         LAYER metal1 ;
	    RECT 267.6000 154.2000 268.0000 154.6000 ;
	    RECT 267.7000 153.8000 268.2000 154.2000 ;
	    RECT 268.6000 127.1000 269.0000 127.6000 ;
	    RECT 269.4000 127.1000 269.8000 127.2000 ;
	    RECT 268.6000 126.8000 269.8000 127.1000 ;
	    RECT 236.2000 86.8000 237.0000 87.2000 ;
	    RECT 245.4000 75.1000 245.8000 75.6000 ;
	    RECT 246.2000 75.1000 246.6000 75.2000 ;
	    RECT 245.4000 74.8000 246.6000 75.1000 ;
         LAYER metal2 ;
	    RECT 267.8000 154.1000 268.2000 154.2000 ;
	    RECT 268.6000 154.1000 269.0000 154.2000 ;
	    RECT 267.8000 153.8000 269.0000 154.1000 ;
	    RECT 269.4000 127.1000 269.8000 127.2000 ;
	    RECT 270.2000 127.1000 270.6000 127.2000 ;
	    RECT 269.4000 126.8000 270.6000 127.1000 ;
	    RECT 236.6000 87.8000 237.0000 88.2000 ;
	    RECT 246.2000 87.8000 246.6000 88.2000 ;
	    RECT 236.6000 87.2000 236.9000 87.8000 ;
	    RECT 236.6000 86.8000 237.0000 87.2000 ;
	    RECT 246.2000 75.2000 246.5000 87.8000 ;
	    RECT 246.2000 74.8000 246.6000 75.2000 ;
         LAYER metal3 ;
	    RECT 267.8000 154.1000 268.2000 154.2000 ;
	    RECT 268.6000 154.1000 269.0000 154.2000 ;
	    RECT 267.8000 153.8000 269.0000 154.1000 ;
	    RECT 267.8000 127.1000 268.2000 127.2000 ;
	    RECT 270.2000 127.1000 270.6000 127.2000 ;
	    RECT 273.4000 127.1000 273.8000 127.2000 ;
	    RECT 267.8000 126.8000 273.8000 127.1000 ;
	    RECT 236.6000 88.1000 237.0000 88.2000 ;
	    RECT 246.2000 88.1000 246.6000 88.2000 ;
	    RECT 267.8000 88.1000 268.2000 88.2000 ;
	    RECT 236.6000 87.8000 268.2000 88.1000 ;
         LAYER metal4 ;
	    RECT 267.8000 153.8000 268.2000 154.2000 ;
	    RECT 267.8000 127.2000 268.1000 153.8000 ;
	    RECT 267.8000 126.8000 268.2000 127.2000 ;
	    RECT 267.8000 88.2000 268.1000 126.8000 ;
	    RECT 267.8000 87.8000 268.2000 88.2000 ;
      END
   END block8[0]
   PIN block8[1]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 50.8000 -2.2000 51.2000 ;
      END
   END block8[1]
   PIN block8[2]
      PORT
         LAYER metal3 ;
	    RECT 273.4000 44.8000 273.8000 45.2000 ;
      END
   END block8[2]
   PIN block8[3]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 156.8000 -2.2000 157.2000 ;
      END
   END block8[3]
   PIN block8[4]
      PORT
         LAYER metal2 ;
	    RECT 240.6000 -2.2000 241.0000 -1.8000 ;
      END
   END block8[4]
   PIN block8[5]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 174.8000 -2.2000 175.2000 ;
      END
   END block8[5]
   PIN block8[6]
      PORT
         LAYER metal3 ;
	    RECT 273.4000 163.8000 273.8000 164.2000 ;
      END
   END block8[6]
   PIN block8[7]
      PORT
         LAYER metal2 ;
	    RECT 4.6000 182.8000 5.0000 183.2000 ;
      END
   END block8[7]
   PIN block9[0]
      PORT
         LAYER metal1 ;
	    RECT 238.2000 127.8000 238.6000 128.6000 ;
	    RECT 250.2000 127.8000 250.6000 128.6000 ;
	    RECT 255.8000 94.8000 256.2000 95.6000 ;
	    RECT 220.2000 93.8000 221.0000 94.2000 ;
         LAYER metal2 ;
	    RECT 238.2000 127.8000 238.6000 128.2000 ;
	    RECT 250.2000 128.1000 250.6000 128.2000 ;
	    RECT 249.4000 127.8000 250.6000 128.1000 ;
	    RECT 238.2000 127.2000 238.5000 127.8000 ;
	    RECT 249.4000 127.2000 249.7000 127.8000 ;
	    RECT 238.2000 126.8000 238.6000 127.2000 ;
	    RECT 249.4000 126.8000 249.8000 127.2000 ;
	    RECT 220.6000 98.8000 221.0000 99.2000 ;
	    RECT 255.8000 98.8000 256.2000 99.2000 ;
	    RECT 220.6000 94.2000 220.9000 98.8000 ;
	    RECT 255.8000 96.2000 256.1000 98.8000 ;
	    RECT 255.8000 95.8000 256.2000 96.2000 ;
	    RECT 255.8000 95.2000 256.1000 95.8000 ;
	    RECT 255.8000 94.8000 256.2000 95.2000 ;
	    RECT 220.6000 93.8000 221.0000 94.2000 ;
         LAYER metal3 ;
	    RECT 238.2000 127.1000 238.6000 127.2000 ;
	    RECT 249.4000 127.1000 249.8000 127.2000 ;
	    RECT 238.2000 126.8000 249.8000 127.1000 ;
	    RECT 220.6000 99.1000 221.0000 99.2000 ;
	    RECT 249.4000 99.1000 249.8000 99.2000 ;
	    RECT 255.8000 99.1000 256.2000 99.2000 ;
	    RECT 220.6000 98.8000 256.2000 99.1000 ;
	    RECT 255.8000 96.1000 256.2000 96.2000 ;
	    RECT 273.4000 96.1000 273.8000 96.2000 ;
	    RECT 255.8000 95.8000 273.8000 96.1000 ;
         LAYER metal4 ;
	    RECT 249.4000 126.8000 249.8000 127.2000 ;
	    RECT 249.4000 99.2000 249.7000 126.8000 ;
	    RECT 249.4000 98.8000 249.8000 99.2000 ;
      END
   END block9[0]
   PIN block9[1]
      PORT
         LAYER metal2 ;
	    RECT 208.6000 182.8000 209.0000 183.2000 ;
      END
   END block9[1]
   PIN block9[2]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 9.8000 -2.2000 10.2000 ;
      END
   END block9[2]
   PIN block9[3]
      PORT
         LAYER metal2 ;
	    RECT 61.4000 -2.2000 61.8000 -1.8000 ;
      END
   END block9[3]
   PIN block9[4]
      PORT
         LAYER metal2 ;
	    RECT 175.0000 182.8000 175.4000 183.2000 ;
      END
   END block9[4]
   PIN block9[5]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 169.8000 -2.2000 170.2000 ;
      END
   END block9[5]
   PIN block9[6]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 163.8000 -2.2000 164.2000 ;
      END
   END block9[6]
   PIN block9[7]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 114.8000 -2.2000 115.2000 ;
      END
   END block9[7]
   PIN block10[0]
      PORT
         LAYER metal1 ;
	    RECT 266.6000 167.1000 267.4000 167.2000 ;
	    RECT 266.3000 167.0000 267.4000 167.1000 ;
	    RECT 265.2000 166.8000 267.4000 167.0000 ;
	    RECT 265.2000 166.7000 266.6000 166.8000 ;
	    RECT 265.2000 166.6000 265.6000 166.7000 ;
	    RECT 264.6000 134.8000 265.0000 135.2000 ;
	    RECT 264.6000 134.4000 264.9000 134.8000 ;
	    RECT 264.4000 134.1000 264.9000 134.4000 ;
	    RECT 264.4000 134.0000 264.8000 134.1000 ;
	    RECT 262.2000 132.4000 262.6000 133.2000 ;
	    RECT 258.2000 87.1000 259.0000 87.2000 ;
	    RECT 258.2000 87.0000 259.3000 87.1000 ;
	    RECT 258.2000 86.8000 260.4000 87.0000 ;
	    RECT 259.0000 86.7000 260.4000 86.8000 ;
	    RECT 260.0000 86.6000 260.4000 86.7000 ;
         LAYER metal2 ;
	    RECT 267.0000 168.8000 267.4000 169.2000 ;
	    RECT 267.0000 167.2000 267.3000 168.8000 ;
	    RECT 267.0000 166.8000 267.4000 167.2000 ;
	    RECT 264.6000 134.8000 265.0000 135.2000 ;
	    RECT 264.6000 133.2000 264.9000 134.8000 ;
	    RECT 262.2000 133.1000 262.6000 133.2000 ;
	    RECT 263.0000 133.1000 263.4000 133.2000 ;
	    RECT 262.2000 132.8000 263.4000 133.1000 ;
	    RECT 264.6000 132.8000 265.0000 133.2000 ;
	    RECT 258.2000 86.8000 258.6000 87.2000 ;
	    RECT 258.2000 86.2000 258.5000 86.8000 ;
	    RECT 258.2000 85.8000 258.6000 86.2000 ;
         LAYER metal3 ;
	    RECT 267.0000 169.1000 267.4000 169.2000 ;
	    RECT 270.2000 169.1000 270.6000 169.2000 ;
	    RECT 273.4000 169.1000 273.8000 169.2000 ;
	    RECT 267.0000 168.8000 273.8000 169.1000 ;
	    RECT 262.2000 133.1000 262.6000 133.2000 ;
	    RECT 263.0000 133.1000 263.4000 133.2000 ;
	    RECT 264.6000 133.1000 265.0000 133.2000 ;
	    RECT 270.2000 133.1000 270.6000 133.2000 ;
	    RECT 262.2000 132.8000 270.6000 133.1000 ;
	    RECT 262.2000 87.1000 262.6000 87.2000 ;
	    RECT 258.2000 86.8000 262.6000 87.1000 ;
	    RECT 258.2000 86.2000 258.5000 86.8000 ;
	    RECT 258.2000 85.8000 258.6000 86.2000 ;
         LAYER metal4 ;
	    RECT 270.2000 168.8000 270.6000 169.2000 ;
	    RECT 270.2000 133.2000 270.5000 168.8000 ;
	    RECT 262.2000 132.8000 262.6000 133.2000 ;
	    RECT 270.2000 132.8000 270.6000 133.2000 ;
	    RECT 262.2000 87.2000 262.5000 132.8000 ;
	    RECT 262.2000 86.8000 262.6000 87.2000 ;
      END
   END block10[0]
   PIN block10[1]
      PORT
         LAYER metal2 ;
	    RECT 258.2000 182.8000 258.6000 183.2000 ;
      END
   END block10[1]
   PIN block10[2]
      PORT
         LAYER metal2 ;
	    RECT 127.8000 182.8000 128.2000 183.2000 ;
      END
   END block10[2]
   PIN block10[3]
      PORT
         LAYER metal2 ;
	    RECT 198.2000 182.8000 198.6000 183.2000 ;
      END
   END block10[3]
   PIN block10[4]
      PORT
         LAYER metal2 ;
	    RECT 63.8000 182.8000 64.2000 183.2000 ;
      END
   END block10[4]
   PIN block10[5]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 158.8000 -2.2000 159.2000 ;
      END
   END block10[5]
   PIN block10[6]
      PORT
         LAYER metal3 ;
	    RECT 273.4000 2.8000 273.8000 3.2000 ;
      END
   END block10[6]
   PIN block10[7]
      PORT
         LAYER metal2 ;
	    RECT 86.2000 182.8000 86.6000 183.2000 ;
      END
   END block10[7]
   PIN block11[0]
      PORT
         LAYER metal1 ;
	    RECT 203.0000 133.4000 203.4000 134.2000 ;
	    RECT 246.2000 134.1000 246.6000 134.2000 ;
	    RECT 245.8000 133.8000 246.6000 134.1000 ;
	    RECT 245.8000 133.6000 246.2000 133.8000 ;
	    RECT 247.8000 127.8000 248.2000 128.6000 ;
	    RECT 255.8000 107.1000 256.6000 107.2000 ;
	    RECT 255.8000 107.0000 256.9000 107.1000 ;
	    RECT 255.8000 106.8000 258.0000 107.0000 ;
	    RECT 256.6000 106.7000 258.0000 106.8000 ;
	    RECT 257.6000 106.6000 258.0000 106.7000 ;
         LAYER metal2 ;
	    RECT 203.0000 134.8000 203.4000 135.2000 ;
	    RECT 203.0000 134.2000 203.3000 134.8000 ;
	    RECT 203.0000 133.8000 203.4000 134.2000 ;
	    RECT 246.2000 133.8000 246.6000 134.2000 ;
	    RECT 247.8000 133.8000 248.2000 134.2000 ;
	    RECT 246.2000 133.2000 246.5000 133.8000 ;
	    RECT 246.2000 132.8000 246.6000 133.2000 ;
	    RECT 247.8000 128.2000 248.1000 133.8000 ;
	    RECT 247.8000 127.8000 248.2000 128.2000 ;
	    RECT 247.8000 120.1000 248.1000 127.8000 ;
	    RECT 248.6000 120.1000 249.0000 120.2000 ;
	    RECT 247.8000 119.8000 249.0000 120.1000 ;
	    RECT 255.8000 109.8000 256.2000 110.2000 ;
	    RECT 255.8000 107.2000 256.1000 109.8000 ;
	    RECT 255.8000 106.8000 256.2000 107.2000 ;
         LAYER metal3 ;
	    RECT 203.0000 134.8000 203.4000 135.2000 ;
	    RECT 203.0000 134.1000 203.3000 134.8000 ;
	    RECT 208.6000 134.1000 209.0000 134.2000 ;
	    RECT 247.8000 134.1000 248.2000 134.2000 ;
	    RECT 203.0000 133.8000 209.0000 134.1000 ;
	    RECT 234.2000 133.8000 248.2000 134.1000 ;
	    RECT 234.2000 133.2000 234.5000 133.8000 ;
	    RECT 246.2000 133.2000 246.5000 133.8000 ;
	    RECT 234.2000 132.8000 234.6000 133.2000 ;
	    RECT 246.2000 132.8000 246.6000 133.2000 ;
	    RECT 247.8000 120.1000 248.2000 120.2000 ;
	    RECT 248.6000 120.1000 249.0000 120.2000 ;
	    RECT 247.8000 119.8000 249.0000 120.1000 ;
	    RECT 247.8000 110.1000 248.2000 110.2000 ;
	    RECT 255.8000 110.1000 256.2000 110.2000 ;
	    RECT 247.8000 109.8000 273.7000 110.1000 ;
	    RECT 273.4000 109.2000 273.7000 109.8000 ;
	    RECT 273.4000 108.8000 273.8000 109.2000 ;
         LAYER metal4 ;
	    RECT 208.6000 134.1000 209.0000 134.2000 ;
	    RECT 209.4000 134.1000 209.8000 134.2000 ;
	    RECT 208.6000 133.8000 209.8000 134.1000 ;
	    RECT 234.2000 133.8000 234.6000 134.2000 ;
	    RECT 234.2000 133.2000 234.5000 133.8000 ;
	    RECT 234.2000 132.8000 234.6000 133.2000 ;
	    RECT 247.8000 119.8000 248.2000 120.2000 ;
	    RECT 247.8000 110.2000 248.1000 119.8000 ;
	    RECT 247.8000 109.8000 248.2000 110.2000 ;
         LAYER metal5 ;
	    RECT 209.4000 134.1000 209.8000 134.2000 ;
	    RECT 234.2000 134.1000 234.6000 134.2000 ;
	    RECT 209.4000 133.8000 234.6000 134.1000 ;
      END
   END block11[0]
   PIN block11[1]
      PORT
         LAYER metal2 ;
	    RECT 183.8000 -2.2000 184.2000 -1.8000 ;
      END
   END block11[1]
   PIN block11[2]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 14.8000 -2.2000 15.2000 ;
      END
   END block11[2]
   PIN block11[3]
      PORT
         LAYER metal3 ;
	    RECT -2.6000 94.8000 -2.2000 95.2000 ;
      END
   END block11[3]
   PIN block11[4]
      PORT
         LAYER metal2 ;
	    RECT 205.4000 -2.2000 205.8000 -1.8000 ;
      END
   END block11[4]
   PIN block11[5]
      PORT
         LAYER metal2 ;
	    RECT 193.4000 -2.2000 193.8000 -1.8000 ;
      END
   END block11[5]
   PIN block11[6]
      PORT
         LAYER metal2 ;
	    RECT 123.8000 -2.2000 124.2000 -1.8000 ;
      END
   END block11[6]
   PIN block11[7]
      PORT
         LAYER metal2 ;
	    RECT 59.8000 182.8000 60.2000 183.2000 ;
      END
   END block11[7]
   PIN start
      PORT
         LAYER metal1 ;
	    RECT 92.2000 156.8000 92.6000 157.2000 ;
	    RECT 92.3000 156.2000 92.6000 156.8000 ;
	    RECT 92.3000 155.9000 93.0000 156.2000 ;
	    RECT 92.6000 155.8000 93.0000 155.9000 ;
	    RECT 86.2000 154.4000 86.6000 155.2000 ;
	    RECT 107.0000 154.1000 107.4000 154.2000 ;
	    RECT 106.6000 153.8000 107.4000 154.1000 ;
	    RECT 109.4000 154.1000 109.8000 154.2000 ;
	    RECT 111.0000 154.1000 111.4000 154.2000 ;
	    RECT 109.4000 153.8000 111.4000 154.1000 ;
	    RECT 106.6000 153.6000 107.0000 153.8000 ;
	    RECT 109.4000 153.4000 109.8000 153.8000 ;
	    RECT 89.4000 152.4000 89.8000 153.2000 ;
	    RECT 120.6000 127.8000 121.0000 128.6000 ;
	    RECT 124.2000 127.2000 124.6000 127.4000 ;
	    RECT 123.8000 126.9000 124.6000 127.2000 ;
	    RECT 123.8000 126.8000 124.2000 126.9000 ;
	    RECT 143.0000 95.1000 143.4000 95.2000 ;
	    RECT 144.6000 95.1000 145.0000 95.2000 ;
	    RECT 143.0000 94.8000 145.0000 95.1000 ;
	    RECT 144.6000 94.4000 145.0000 94.8000 ;
	    RECT 143.0000 94.1000 143.4000 94.2000 ;
	    RECT 142.6000 93.8000 143.4000 94.1000 ;
	    RECT 142.6000 93.6000 143.0000 93.8000 ;
	    RECT 140.6000 75.1000 141.0000 75.2000 ;
	    RECT 142.2000 75.1000 142.6000 75.2000 ;
	    RECT 140.6000 74.8000 142.6000 75.1000 ;
	    RECT 142.2000 74.4000 142.6000 74.8000 ;
	    RECT 156.6000 54.1000 157.0000 54.2000 ;
	    RECT 156.6000 53.8000 157.4000 54.1000 ;
	    RECT 157.0000 53.6000 157.4000 53.8000 ;
         LAYER metal2 ;
	    RECT 93.4000 183.1000 93.8000 183.2000 ;
	    RECT 93.4000 182.8000 94.5000 183.1000 ;
	    RECT 92.6000 155.8000 93.0000 156.2000 ;
	    RECT 92.6000 155.2000 92.9000 155.8000 ;
	    RECT 94.2000 155.2000 94.5000 182.8000 ;
	    RECT 86.2000 155.1000 86.6000 155.2000 ;
	    RECT 87.0000 155.1000 87.4000 155.2000 ;
	    RECT 86.2000 154.8000 87.4000 155.1000 ;
	    RECT 89.4000 154.8000 89.8000 155.2000 ;
	    RECT 92.6000 154.8000 93.0000 155.2000 ;
	    RECT 94.2000 154.8000 94.6000 155.2000 ;
	    RECT 107.0000 154.8000 107.4000 155.2000 ;
	    RECT 109.4000 154.8000 109.8000 155.2000 ;
	    RECT 89.4000 153.2000 89.7000 154.8000 ;
	    RECT 107.0000 154.2000 107.3000 154.8000 ;
	    RECT 109.4000 154.2000 109.7000 154.8000 ;
	    RECT 107.0000 153.8000 107.4000 154.2000 ;
	    RECT 109.4000 153.8000 109.8000 154.2000 ;
	    RECT 111.0000 153.8000 111.4000 154.2000 ;
	    RECT 89.4000 152.8000 89.8000 153.2000 ;
	    RECT 111.0000 137.2000 111.3000 153.8000 ;
	    RECT 111.0000 136.8000 111.4000 137.2000 ;
	    RECT 120.6000 136.8000 121.0000 137.2000 ;
	    RECT 120.6000 128.2000 120.9000 136.8000 ;
	    RECT 120.6000 127.8000 121.0000 128.2000 ;
	    RECT 123.8000 127.8000 124.2000 128.2000 ;
	    RECT 123.8000 127.2000 124.1000 127.8000 ;
	    RECT 123.8000 126.8000 124.2000 127.2000 ;
	    RECT 140.6000 94.8000 141.0000 95.2000 ;
	    RECT 143.0000 94.8000 143.4000 95.2000 ;
	    RECT 140.6000 75.2000 140.9000 94.8000 ;
	    RECT 143.0000 94.2000 143.3000 94.8000 ;
	    RECT 143.0000 93.8000 143.4000 94.2000 ;
	    RECT 140.6000 74.8000 141.0000 75.2000 ;
	    RECT 140.6000 70.2000 140.9000 74.8000 ;
	    RECT 140.6000 69.8000 141.0000 70.2000 ;
	    RECT 156.6000 69.8000 157.0000 70.2000 ;
	    RECT 156.6000 54.2000 156.9000 69.8000 ;
	    RECT 156.6000 53.8000 157.0000 54.2000 ;
         LAYER metal3 ;
	    RECT 87.0000 155.1000 87.4000 155.2000 ;
	    RECT 89.4000 155.1000 89.8000 155.2000 ;
	    RECT 92.6000 155.1000 93.0000 155.2000 ;
	    RECT 94.2000 155.1000 94.6000 155.2000 ;
	    RECT 107.0000 155.1000 107.4000 155.2000 ;
	    RECT 109.4000 155.1000 109.8000 155.2000 ;
	    RECT 87.0000 154.8000 109.8000 155.1000 ;
	    RECT 111.0000 137.1000 111.4000 137.2000 ;
	    RECT 120.6000 137.1000 121.0000 137.2000 ;
	    RECT 111.0000 136.8000 121.0000 137.1000 ;
	    RECT 120.6000 128.1000 121.0000 128.2000 ;
	    RECT 123.8000 128.1000 124.2000 128.2000 ;
	    RECT 125.4000 128.1000 125.8000 128.2000 ;
	    RECT 120.6000 127.8000 125.8000 128.1000 ;
	    RECT 125.4000 95.1000 125.8000 95.2000 ;
	    RECT 140.6000 95.1000 141.0000 95.2000 ;
	    RECT 143.0000 95.1000 143.4000 95.2000 ;
	    RECT 125.4000 94.8000 143.4000 95.1000 ;
	    RECT 140.6000 70.1000 141.0000 70.2000 ;
	    RECT 156.6000 70.1000 157.0000 70.2000 ;
	    RECT 140.6000 69.8000 157.0000 70.1000 ;
         LAYER metal4 ;
	    RECT 125.4000 127.8000 125.8000 128.2000 ;
	    RECT 125.4000 95.2000 125.7000 127.8000 ;
	    RECT 125.4000 94.8000 125.8000 95.2000 ;
      END
   END start
   PIN target[0]
      PORT
         LAYER metal1 ;
	    RECT 24.6000 54.1000 25.4000 54.2000 ;
	    RECT 24.6000 53.8000 26.3000 54.1000 ;
	    RECT 26.0000 53.6000 26.3000 53.8000 ;
	    RECT 28.0000 53.8000 28.4000 54.2000 ;
	    RECT 28.0000 53.6000 28.3000 53.8000 ;
	    RECT 26.0000 53.3000 27.0000 53.6000 ;
	    RECT 26.2000 53.2000 27.0000 53.3000 ;
	    RECT 27.9000 53.2000 28.3000 53.6000 ;
	    RECT 33.4000 52.4000 33.8000 53.2000 ;
	    RECT 23.8000 47.8000 24.2000 48.6000 ;
	    RECT 27.8000 47.8000 28.2000 48.6000 ;
	    RECT 33.4000 47.7000 34.2000 47.8000 ;
	    RECT 33.2000 47.4000 34.2000 47.7000 ;
	    RECT 35.1000 47.4000 35.5000 47.8000 ;
	    RECT 33.2000 47.2000 33.5000 47.4000 ;
	    RECT 31.8000 46.9000 33.5000 47.2000 ;
	    RECT 35.2000 47.2000 35.5000 47.4000 ;
	    RECT 31.8000 46.8000 32.6000 46.9000 ;
	    RECT 35.2000 46.8000 35.6000 47.2000 ;
	    RECT 28.6000 32.4000 29.0000 33.2000 ;
         LAYER metal2 ;
	    RECT 24.6000 53.8000 25.0000 54.2000 ;
	    RECT 24.6000 50.2000 24.9000 53.8000 ;
	    RECT 26.2000 53.5000 26.6000 53.6000 ;
	    RECT 27.9000 53.5000 28.3000 53.6000 ;
	    RECT 26.2000 53.2000 28.3000 53.5000 ;
	    RECT 33.4000 52.8000 33.8000 53.2000 ;
	    RECT 24.6000 49.8000 25.0000 50.2000 ;
	    RECT 23.8000 47.8000 24.2000 48.2000 ;
	    RECT 23.8000 46.2000 24.1000 47.8000 ;
	    RECT 24.6000 46.2000 24.9000 49.8000 ;
	    RECT 27.8000 48.1000 28.2000 48.2000 ;
	    RECT 27.8000 47.8000 28.9000 48.1000 ;
	    RECT 28.6000 46.2000 28.9000 47.8000 ;
	    RECT 33.4000 47.8000 33.7000 52.8000 ;
	    RECT 33.4000 47.5000 35.5000 47.8000 ;
	    RECT 33.4000 47.4000 33.8000 47.5000 ;
	    RECT 35.1000 47.4000 35.5000 47.5000 ;
	    RECT 31.8000 46.8000 32.2000 47.2000 ;
	    RECT 31.8000 46.2000 32.1000 46.8000 ;
	    RECT 23.8000 45.8000 24.2000 46.2000 ;
	    RECT 24.6000 45.8000 25.0000 46.2000 ;
	    RECT 28.6000 45.8000 29.0000 46.2000 ;
	    RECT 31.8000 45.8000 32.2000 46.2000 ;
	    RECT 28.6000 33.2000 28.9000 45.8000 ;
	    RECT 28.6000 32.8000 29.0000 33.2000 ;
         LAYER metal3 ;
	    RECT 24.6000 50.1000 25.0000 50.2000 ;
	    RECT -2.6000 49.8000 25.0000 50.1000 ;
	    RECT -2.6000 49.2000 -2.3000 49.8000 ;
	    RECT -2.6000 48.8000 -2.2000 49.2000 ;
	    RECT 23.8000 46.1000 24.2000 46.2000 ;
	    RECT 24.6000 46.1000 25.0000 46.2000 ;
	    RECT 28.6000 46.1000 29.0000 46.2000 ;
	    RECT 31.8000 46.1000 32.2000 46.2000 ;
	    RECT 23.8000 45.8000 32.2000 46.1000 ;
      END
   END target[0]
   PIN target[1]
      PORT
         LAYER metal1 ;
	    RECT 15.0000 52.4000 15.4000 53.2000 ;
	    RECT 41.4000 47.8000 41.8000 48.6000 ;
	    RECT 19.8000 47.7000 20.6000 47.8000 ;
	    RECT 19.6000 47.4000 20.6000 47.7000 ;
	    RECT 21.5000 47.4000 21.9000 47.8000 ;
	    RECT 19.6000 47.2000 19.9000 47.4000 ;
	    RECT 18.2000 46.9000 19.9000 47.2000 ;
	    RECT 21.6000 47.2000 21.9000 47.4000 ;
	    RECT 18.2000 46.8000 19.0000 46.9000 ;
	    RECT 21.6000 46.8000 22.0000 47.2000 ;
	    RECT 40.6000 47.1000 41.0000 47.2000 ;
	    RECT 41.4000 47.1000 41.7000 47.8000 ;
	    RECT 40.6000 46.8000 41.7000 47.1000 ;
	    RECT 13.4000 33.4000 13.8000 34.2000 ;
	    RECT 37.2000 33.8000 37.6000 34.2000 ;
	    RECT 40.2000 34.1000 41.0000 34.2000 ;
	    RECT 37.3000 33.6000 37.6000 33.8000 ;
	    RECT 39.3000 33.8000 41.0000 34.1000 ;
	    RECT 39.3000 33.6000 39.6000 33.8000 ;
	    RECT 37.3000 33.2000 37.7000 33.6000 ;
	    RECT 38.6000 33.3000 39.6000 33.6000 ;
	    RECT 38.6000 33.2000 39.4000 33.3000 ;
	    RECT 17.4000 32.4000 17.8000 33.2000 ;
	    RECT 28.6000 27.8000 29.0000 28.6000 ;
	    RECT 28.6000 27.1000 28.9000 27.8000 ;
	    RECT 29.4000 27.1000 29.8000 27.6000 ;
	    RECT 28.6000 26.8000 29.8000 27.1000 ;
         LAYER metal2 ;
	    RECT 15.0000 52.8000 15.4000 53.2000 ;
	    RECT 18.2000 52.8000 18.6000 53.2000 ;
	    RECT 15.0000 52.2000 15.3000 52.8000 ;
	    RECT 15.0000 51.8000 15.4000 52.2000 ;
	    RECT 18.2000 47.2000 18.5000 52.8000 ;
	    RECT 19.8000 47.5000 21.9000 47.8000 ;
	    RECT 19.8000 47.4000 20.2000 47.5000 ;
	    RECT 21.5000 47.4000 21.9000 47.5000 ;
	    RECT 18.2000 46.8000 18.6000 47.2000 ;
	    RECT 40.6000 46.8000 41.0000 47.2000 ;
	    RECT 18.2000 45.1000 18.5000 46.8000 ;
	    RECT 17.4000 44.8000 18.5000 45.1000 ;
	    RECT 13.4000 35.8000 13.8000 36.2000 ;
	    RECT 13.4000 34.2000 13.7000 35.8000 ;
	    RECT 13.4000 33.8000 13.8000 34.2000 ;
	    RECT 13.4000 31.2000 13.7000 33.8000 ;
	    RECT 17.4000 33.2000 17.7000 44.8000 ;
	    RECT 40.6000 34.2000 40.9000 46.8000 ;
	    RECT 40.6000 33.8000 41.0000 34.2000 ;
	    RECT 37.3000 33.5000 37.7000 33.6000 ;
	    RECT 39.0000 33.5000 39.4000 33.6000 ;
	    RECT 37.3000 33.2000 39.4000 33.5000 ;
	    RECT 17.4000 32.8000 17.8000 33.2000 ;
	    RECT 17.4000 31.2000 17.7000 32.8000 ;
	    RECT 40.6000 31.2000 40.9000 33.8000 ;
	    RECT 13.4000 30.8000 13.8000 31.2000 ;
	    RECT 17.4000 30.8000 17.8000 31.2000 ;
	    RECT 28.6000 30.8000 29.0000 31.2000 ;
	    RECT 40.6000 30.8000 41.0000 31.2000 ;
	    RECT 28.6000 28.2000 28.9000 30.8000 ;
	    RECT 28.6000 27.8000 29.0000 28.2000 ;
         LAYER metal3 ;
	    RECT 18.2000 53.1000 18.6000 53.2000 ;
	    RECT 15.0000 52.8000 18.6000 53.1000 ;
	    RECT 15.0000 52.2000 15.3000 52.8000 ;
	    RECT 15.0000 51.8000 15.4000 52.2000 ;
	    RECT -2.6000 36.1000 -2.2000 36.2000 ;
	    RECT 13.4000 36.1000 13.8000 36.2000 ;
	    RECT -2.6000 35.8000 13.8000 36.1000 ;
	    RECT 13.4000 31.1000 13.8000 31.2000 ;
	    RECT 17.4000 31.1000 17.8000 31.2000 ;
	    RECT 28.6000 31.1000 29.0000 31.2000 ;
	    RECT 40.6000 31.1000 41.0000 31.2000 ;
	    RECT 13.4000 30.8000 41.0000 31.1000 ;
      END
   END target[1]
   PIN target[2]
      PORT
         LAYER metal1 ;
	    RECT 0.6000 54.1000 1.4000 54.2000 ;
	    RECT 0.6000 53.8000 2.3000 54.1000 ;
	    RECT 2.0000 53.6000 2.3000 53.8000 ;
	    RECT 4.0000 53.8000 4.4000 54.2000 ;
	    RECT 4.0000 53.6000 4.3000 53.8000 ;
	    RECT 2.0000 53.3000 3.0000 53.6000 ;
	    RECT 2.2000 53.2000 3.0000 53.3000 ;
	    RECT 3.9000 53.2000 4.3000 53.6000 ;
	    RECT 6.2000 52.4000 6.6000 53.2000 ;
	    RECT 5.0000 47.1000 5.8000 47.2000 ;
	    RECT 4.7000 47.0000 5.8000 47.1000 ;
	    RECT 3.6000 46.8000 5.8000 47.0000 ;
	    RECT 3.6000 46.7000 5.0000 46.8000 ;
	    RECT 3.6000 46.6000 4.0000 46.7000 ;
	    RECT 6.2000 34.8000 6.6000 35.2000 ;
	    RECT 6.2000 34.2000 6.5000 34.8000 ;
	    RECT 8.0000 34.3000 8.4000 34.4000 ;
	    RECT 7.0000 34.2000 8.4000 34.3000 ;
	    RECT 0.6000 34.1000 1.4000 34.2000 ;
	    RECT 0.6000 33.8000 2.3000 34.1000 ;
	    RECT 2.0000 33.6000 2.3000 33.8000 ;
	    RECT 4.0000 33.8000 4.4000 34.2000 ;
	    RECT 6.2000 34.0000 8.4000 34.2000 ;
	    RECT 6.2000 33.9000 7.3000 34.0000 ;
	    RECT 6.2000 33.8000 7.0000 33.9000 ;
	    RECT 4.0000 33.6000 4.3000 33.8000 ;
	    RECT 2.0000 33.3000 3.0000 33.6000 ;
	    RECT 2.2000 33.2000 3.0000 33.3000 ;
	    RECT 3.9000 33.2000 4.3000 33.6000 ;
	    RECT 0.6000 27.8000 1.0000 28.6000 ;
         LAYER metal2 ;
	    RECT 0.6000 53.8000 1.0000 54.2000 ;
	    RECT 0.6000 53.2000 0.9000 53.8000 ;
	    RECT 2.2000 53.5000 2.6000 53.6000 ;
	    RECT 3.9000 53.5000 4.3000 53.6000 ;
	    RECT 2.2000 53.2000 4.3000 53.5000 ;
	    RECT 0.6000 52.8000 1.0000 53.2000 ;
	    RECT 6.2000 52.8000 6.6000 53.2000 ;
	    RECT 6.2000 51.1000 6.5000 52.8000 ;
	    RECT 5.4000 50.8000 6.5000 51.1000 ;
	    RECT 5.4000 47.2000 5.7000 50.8000 ;
	    RECT 5.4000 46.8000 5.8000 47.2000 ;
	    RECT 0.6000 34.8000 1.0000 35.2000 ;
	    RECT 5.4000 35.1000 5.7000 46.8000 ;
	    RECT 6.2000 35.1000 6.6000 35.2000 ;
	    RECT 5.4000 34.8000 6.6000 35.1000 ;
	    RECT 0.6000 34.2000 0.9000 34.8000 ;
	    RECT 6.2000 34.2000 6.5000 34.8000 ;
	    RECT 0.6000 33.8000 1.0000 34.2000 ;
	    RECT 6.2000 33.8000 6.6000 34.2000 ;
	    RECT 0.6000 28.2000 0.9000 33.8000 ;
	    RECT 2.2000 33.5000 2.6000 33.6000 ;
	    RECT 3.9000 33.5000 4.3000 33.6000 ;
	    RECT 2.2000 33.2000 4.3000 33.5000 ;
	    RECT 0.6000 27.8000 1.0000 28.2000 ;
         LAYER metal3 ;
	    RECT 0.6000 53.1000 1.0000 53.2000 ;
	    RECT 6.2000 53.1000 6.6000 53.2000 ;
	    RECT 0.6000 52.8000 6.6000 53.1000 ;
	    RECT 0.6000 34.8000 1.0000 35.2000 ;
	    RECT 0.6000 34.1000 0.9000 34.8000 ;
	    RECT 6.2000 34.1000 6.6000 34.2000 ;
	    RECT 0.6000 33.8000 6.6000 34.1000 ;
	    RECT -2.6000 28.1000 -2.2000 28.2000 ;
	    RECT 0.6000 28.1000 1.0000 28.2000 ;
	    RECT -2.6000 27.8000 1.0000 28.1000 ;
      END
   END target[2]
   PIN target[3]
      PORT
         LAYER metal1 ;
	    RECT 0.6000 67.8000 1.0000 68.6000 ;
	    RECT 15.0000 47.8000 15.4000 48.6000 ;
	    RECT 6.2000 46.8000 6.6000 47.6000 ;
	    RECT 21.4000 32.4000 21.8000 33.2000 ;
	    RECT 13.4000 27.8000 13.8000 28.6000 ;
	    RECT 13.4000 27.1000 13.7000 27.8000 ;
	    RECT 14.2000 27.1000 14.6000 27.6000 ;
	    RECT 13.4000 26.8000 14.6000 27.1000 ;
         LAYER metal2 ;
	    RECT 0.6000 67.8000 1.0000 68.2000 ;
	    RECT 0.6000 67.2000 0.9000 67.8000 ;
	    RECT 0.6000 66.8000 1.0000 67.2000 ;
	    RECT 7.0000 66.8000 7.4000 67.2000 ;
	    RECT 7.0000 47.2000 7.3000 66.8000 ;
	    RECT 14.2000 48.1000 14.6000 48.2000 ;
	    RECT 15.0000 48.1000 15.4000 48.2000 ;
	    RECT 14.2000 47.8000 15.4000 48.1000 ;
	    RECT 6.2000 47.1000 6.6000 47.2000 ;
	    RECT 7.0000 47.1000 7.4000 47.2000 ;
	    RECT 6.2000 46.8000 7.4000 47.1000 ;
	    RECT 21.4000 32.8000 21.8000 33.2000 ;
	    RECT 21.4000 32.2000 21.7000 32.8000 ;
	    RECT 14.2000 31.8000 14.6000 32.2000 ;
	    RECT 21.4000 31.8000 21.8000 32.2000 ;
	    RECT 14.2000 27.2000 14.5000 31.8000 ;
	    RECT 14.2000 26.8000 14.6000 27.2000 ;
         LAYER metal3 ;
	    RECT -2.6000 67.1000 -2.2000 67.2000 ;
	    RECT 0.6000 67.1000 1.0000 67.2000 ;
	    RECT 7.0000 67.1000 7.4000 67.2000 ;
	    RECT -2.6000 66.8000 7.4000 67.1000 ;
	    RECT 14.2000 47.8000 14.6000 48.2000 ;
	    RECT 14.2000 47.2000 14.5000 47.8000 ;
	    RECT 7.0000 47.1000 7.4000 47.2000 ;
	    RECT 14.2000 47.1000 14.6000 47.2000 ;
	    RECT 7.0000 46.8000 14.6000 47.1000 ;
	    RECT 14.2000 32.1000 14.6000 32.2000 ;
	    RECT 21.4000 32.1000 21.8000 32.2000 ;
	    RECT 14.2000 31.8000 21.8000 32.1000 ;
         LAYER metal4 ;
	    RECT 14.2000 46.8000 14.6000 47.2000 ;
	    RECT 14.2000 32.2000 14.5000 46.8000 ;
	    RECT 14.2000 31.8000 14.6000 32.2000 ;
      END
   END target[3]
   PIN target[4]
      PORT
         LAYER metal1 ;
	    RECT 6.2000 92.4000 6.6000 93.2000 ;
	    RECT 8.6000 85.4000 9.0000 86.2000 ;
	    RECT 13.4000 74.8000 13.8000 75.6000 ;
	    RECT 0.6000 72.4000 1.0000 73.2000 ;
         LAYER metal2 ;
	    RECT 6.2000 92.8000 6.6000 93.2000 ;
	    RECT 6.2000 92.2000 6.5000 92.8000 ;
	    RECT 6.2000 91.8000 6.6000 92.2000 ;
	    RECT 8.6000 91.8000 9.0000 92.2000 ;
	    RECT 8.6000 86.2000 8.9000 91.8000 ;
	    RECT 8.6000 86.1000 9.0000 86.2000 ;
	    RECT 8.6000 85.8000 9.7000 86.1000 ;
	    RECT 9.4000 76.2000 9.7000 85.8000 ;
	    RECT 0.6000 75.8000 1.0000 76.2000 ;
	    RECT 9.4000 75.8000 9.8000 76.2000 ;
	    RECT 13.4000 75.8000 13.8000 76.2000 ;
	    RECT 0.6000 73.2000 0.9000 75.8000 ;
	    RECT 13.4000 75.2000 13.7000 75.8000 ;
	    RECT 13.4000 74.8000 13.8000 75.2000 ;
	    RECT 0.6000 72.8000 1.0000 73.2000 ;
         LAYER metal3 ;
	    RECT 6.2000 92.1000 6.6000 92.2000 ;
	    RECT 8.6000 92.1000 9.0000 92.2000 ;
	    RECT 6.2000 91.8000 9.0000 92.1000 ;
	    RECT -2.6000 76.1000 -2.2000 76.2000 ;
	    RECT 0.6000 76.1000 1.0000 76.2000 ;
	    RECT 9.4000 76.1000 9.8000 76.2000 ;
	    RECT 13.4000 76.1000 13.8000 76.2000 ;
	    RECT -2.6000 75.8000 13.8000 76.1000 ;
      END
   END target[4]
   PIN target[5]
      PORT
         LAYER metal1 ;
	    RECT 0.6000 92.4000 1.0000 93.2000 ;
	    RECT 2.2000 86.1000 2.6000 86.6000 ;
	    RECT 6.2000 86.4000 6.6000 87.2000 ;
	    RECT 3.0000 86.1000 3.4000 86.2000 ;
	    RECT 2.2000 85.8000 3.4000 86.1000 ;
	    RECT 15.8000 73.8000 16.2000 74.6000 ;
	    RECT 19.0000 74.4000 19.4000 75.2000 ;
	    RECT 11.0000 72.4000 11.4000 73.2000 ;
         LAYER metal2 ;
	    RECT 0.6000 93.8000 1.0000 94.2000 ;
	    RECT 0.6000 93.2000 0.9000 93.8000 ;
	    RECT 0.6000 92.8000 1.0000 93.2000 ;
	    RECT 0.6000 87.2000 0.9000 92.8000 ;
	    RECT 0.6000 86.8000 1.0000 87.2000 ;
	    RECT 3.0000 86.8000 3.4000 87.2000 ;
	    RECT 6.2000 86.8000 6.6000 87.2000 ;
	    RECT 3.0000 86.2000 3.3000 86.8000 ;
	    RECT 3.0000 85.8000 3.4000 86.2000 ;
	    RECT 3.0000 82.2000 3.3000 85.8000 ;
	    RECT 6.2000 82.2000 6.5000 86.8000 ;
	    RECT 3.0000 81.8000 3.4000 82.2000 ;
	    RECT 6.2000 81.8000 6.6000 82.2000 ;
	    RECT 11.0000 81.8000 11.4000 82.2000 ;
	    RECT 11.0000 75.2000 11.3000 81.8000 ;
	    RECT 11.0000 74.8000 11.4000 75.2000 ;
	    RECT 15.8000 74.8000 16.2000 75.2000 ;
	    RECT 18.2000 75.1000 18.6000 75.2000 ;
	    RECT 19.0000 75.1000 19.4000 75.2000 ;
	    RECT 18.2000 74.8000 19.4000 75.1000 ;
	    RECT 11.0000 73.2000 11.3000 74.8000 ;
	    RECT 15.8000 74.2000 16.1000 74.8000 ;
	    RECT 15.8000 73.8000 16.2000 74.2000 ;
	    RECT 11.0000 72.8000 11.4000 73.2000 ;
         LAYER metal3 ;
	    RECT -2.6000 97.1000 -2.2000 97.2000 ;
	    RECT 0.6000 97.1000 1.0000 97.2000 ;
	    RECT -2.6000 96.8000 1.0000 97.1000 ;
	    RECT 0.6000 94.8000 1.0000 95.2000 ;
	    RECT 0.6000 94.2000 0.9000 94.8000 ;
	    RECT 0.6000 93.8000 1.0000 94.2000 ;
	    RECT 0.6000 87.1000 1.0000 87.2000 ;
	    RECT 3.0000 87.1000 3.4000 87.2000 ;
	    RECT 0.6000 86.8000 3.4000 87.1000 ;
	    RECT 3.0000 82.1000 3.4000 82.2000 ;
	    RECT 6.2000 82.1000 6.6000 82.2000 ;
	    RECT 11.0000 82.1000 11.4000 82.2000 ;
	    RECT 3.0000 81.8000 11.4000 82.1000 ;
	    RECT 11.0000 75.1000 11.4000 75.2000 ;
	    RECT 15.8000 75.1000 16.2000 75.2000 ;
	    RECT 18.2000 75.1000 18.6000 75.2000 ;
	    RECT 11.0000 74.8000 18.6000 75.1000 ;
         LAYER metal4 ;
	    RECT 0.6000 96.8000 1.0000 97.2000 ;
	    RECT 0.6000 95.2000 0.9000 96.8000 ;
	    RECT 0.6000 94.8000 1.0000 95.2000 ;
      END
   END target[5]
   PIN target[6]
      PORT
         LAYER metal1 ;
	    RECT 0.6000 112.4000 1.0000 113.2000 ;
	    RECT 19.8000 107.8000 20.2000 108.6000 ;
	    RECT 15.7000 107.4000 16.1000 107.8000 ;
	    RECT 17.0000 107.7000 17.8000 107.8000 ;
	    RECT 17.0000 107.4000 18.0000 107.7000 ;
	    RECT 15.7000 107.2000 16.0000 107.4000 ;
	    RECT 15.6000 106.8000 16.0000 107.2000 ;
	    RECT 17.7000 107.2000 18.0000 107.4000 ;
	    RECT 17.7000 107.1000 19.4000 107.2000 ;
	    RECT 19.8000 107.1000 20.2000 107.2000 ;
	    RECT 17.7000 106.9000 20.2000 107.1000 ;
	    RECT 18.6000 106.8000 20.2000 106.9000 ;
	    RECT 20.4000 94.3000 20.8000 94.4000 ;
	    RECT 20.4000 94.2000 21.8000 94.3000 ;
	    RECT 20.4000 94.0000 22.6000 94.2000 ;
	    RECT 21.5000 93.9000 22.6000 94.0000 ;
	    RECT 21.8000 93.8000 22.6000 93.9000 ;
	    RECT 23.0000 87.7000 23.8000 87.8000 ;
	    RECT 22.8000 87.4000 23.8000 87.7000 ;
	    RECT 24.7000 87.4000 25.1000 87.8000 ;
	    RECT 22.8000 87.2000 23.1000 87.4000 ;
	    RECT 21.4000 86.9000 23.1000 87.2000 ;
	    RECT 24.8000 87.2000 25.1000 87.4000 ;
	    RECT 21.4000 86.8000 22.2000 86.9000 ;
	    RECT 24.8000 86.8000 25.2000 87.2000 ;
	    RECT 32.6000 87.1000 33.4000 87.2000 ;
	    RECT 32.6000 87.0000 33.7000 87.1000 ;
	    RECT 32.6000 86.8000 34.8000 87.0000 ;
	    RECT 32.6000 86.2000 32.9000 86.8000 ;
	    RECT 33.4000 86.7000 34.8000 86.8000 ;
	    RECT 34.4000 86.6000 34.8000 86.7000 ;
	    RECT 32.6000 85.8000 33.0000 86.2000 ;
         LAYER metal2 ;
	    RECT 0.6000 116.8000 1.0000 117.2000 ;
	    RECT 16.6000 116.8000 17.0000 117.2000 ;
	    RECT 0.6000 113.2000 0.9000 116.8000 ;
	    RECT 0.6000 112.8000 1.0000 113.2000 ;
	    RECT 16.6000 107.8000 16.9000 116.8000 ;
	    RECT 19.8000 107.8000 20.2000 108.2000 ;
	    RECT 15.7000 107.5000 17.8000 107.8000 ;
	    RECT 15.7000 107.4000 16.1000 107.5000 ;
	    RECT 17.4000 107.4000 17.8000 107.5000 ;
	    RECT 19.8000 107.2000 20.1000 107.8000 ;
	    RECT 19.8000 106.8000 20.2000 107.2000 ;
	    RECT 19.8000 105.2000 20.1000 106.8000 ;
	    RECT 19.8000 104.8000 20.2000 105.2000 ;
	    RECT 22.2000 104.8000 22.6000 105.2000 ;
	    RECT 22.2000 94.2000 22.5000 104.8000 ;
	    RECT 22.2000 93.8000 22.6000 94.2000 ;
	    RECT 22.2000 92.1000 22.5000 93.8000 ;
	    RECT 21.4000 91.8000 22.5000 92.1000 ;
	    RECT 21.4000 88.2000 21.7000 91.8000 ;
	    RECT 21.4000 87.8000 21.8000 88.2000 ;
	    RECT 21.4000 87.2000 21.7000 87.8000 ;
	    RECT 23.0000 87.5000 25.1000 87.8000 ;
	    RECT 23.0000 87.4000 23.4000 87.5000 ;
	    RECT 24.7000 87.4000 25.1000 87.5000 ;
	    RECT 21.4000 86.8000 21.8000 87.2000 ;
	    RECT 32.6000 86.8000 33.0000 87.2000 ;
	    RECT 32.6000 86.2000 32.9000 86.8000 ;
	    RECT 32.6000 85.8000 33.0000 86.2000 ;
         LAYER metal3 ;
	    RECT -2.6000 117.1000 -2.2000 117.2000 ;
	    RECT 0.6000 117.1000 1.0000 117.2000 ;
	    RECT 16.6000 117.1000 17.0000 117.2000 ;
	    RECT -2.6000 116.8000 17.0000 117.1000 ;
	    RECT 19.8000 105.1000 20.2000 105.2000 ;
	    RECT 22.2000 105.1000 22.6000 105.2000 ;
	    RECT 19.8000 104.8000 22.6000 105.1000 ;
	    RECT 21.4000 87.8000 21.8000 88.2000 ;
	    RECT 21.4000 87.1000 21.7000 87.8000 ;
	    RECT 32.6000 87.1000 33.0000 87.2000 ;
	    RECT 21.4000 86.8000 33.0000 87.1000 ;
      END
   END target[6]
   PIN target[7]
      PORT
         LAYER metal1 ;
	    RECT 11.8000 113.8000 12.6000 114.2000 ;
	    RECT 11.0000 112.4000 11.4000 113.2000 ;
	    RECT 35.0000 92.4000 35.4000 93.2000 ;
	    RECT 15.4000 86.8000 16.2000 87.2000 ;
	    RECT 27.0000 86.8000 27.8000 87.2000 ;
	    RECT 35.8000 73.8000 36.6000 74.2000 ;
         LAYER metal2 ;
	    RECT 11.8000 113.8000 12.2000 114.2000 ;
	    RECT 11.8000 113.2000 12.1000 113.8000 ;
	    RECT 11.0000 113.1000 11.4000 113.2000 ;
	    RECT 11.8000 113.1000 12.2000 113.2000 ;
	    RECT 11.0000 112.8000 12.2000 113.1000 ;
	    RECT 35.0000 92.8000 35.4000 93.2000 ;
	    RECT 35.0000 92.2000 35.3000 92.8000 ;
	    RECT 35.0000 91.8000 35.4000 92.2000 ;
	    RECT 15.8000 86.8000 16.2000 87.2000 ;
	    RECT 27.0000 86.8000 27.4000 87.2000 ;
	    RECT 15.8000 85.2000 16.1000 86.8000 ;
	    RECT 27.0000 85.2000 27.3000 86.8000 ;
	    RECT 15.8000 84.8000 16.2000 85.2000 ;
	    RECT 27.0000 84.8000 27.4000 85.2000 ;
	    RECT 35.8000 84.8000 36.2000 85.2000 ;
	    RECT 35.8000 74.2000 36.1000 84.8000 ;
	    RECT 35.8000 73.8000 36.2000 74.2000 ;
         LAYER metal3 ;
	    RECT -2.6000 113.1000 -2.2000 113.2000 ;
	    RECT 11.0000 113.1000 11.4000 113.2000 ;
	    RECT 11.8000 113.1000 12.2000 113.2000 ;
	    RECT -2.6000 112.8000 12.2000 113.1000 ;
	    RECT 35.0000 92.8000 35.4000 93.2000 ;
	    RECT 35.0000 92.2000 35.3000 92.8000 ;
	    RECT 35.0000 91.8000 35.4000 92.2000 ;
	    RECT 11.0000 85.1000 11.4000 85.2000 ;
	    RECT 15.8000 85.1000 16.2000 85.2000 ;
	    RECT 27.0000 85.1000 27.4000 85.2000 ;
	    RECT 35.0000 85.1000 35.4000 85.2000 ;
	    RECT 35.8000 85.1000 36.2000 85.2000 ;
	    RECT 11.0000 84.8000 36.2000 85.1000 ;
         LAYER metal4 ;
	    RECT 11.0000 112.8000 11.4000 113.2000 ;
	    RECT 11.0000 85.2000 11.3000 112.8000 ;
	    RECT 35.0000 92.8000 35.4000 93.2000 ;
	    RECT 35.0000 85.2000 35.3000 92.8000 ;
	    RECT 11.0000 84.8000 11.4000 85.2000 ;
	    RECT 35.0000 84.8000 35.4000 85.2000 ;
      END
   END target[7]
   PIN target[8]
      PORT
         LAYER metal1 ;
	    RECT 11.8000 172.4000 12.2000 173.2000 ;
	    RECT 14.2000 165.4000 14.6000 166.2000 ;
	    RECT 2.2000 154.8000 2.6000 155.6000 ;
	    RECT 7.8000 152.4000 8.2000 153.2000 ;
         LAYER metal2 ;
	    RECT 11.8000 172.8000 12.2000 173.2000 ;
	    RECT 11.8000 171.2000 12.1000 172.8000 ;
	    RECT 11.8000 170.8000 12.2000 171.2000 ;
	    RECT 14.2000 170.8000 14.6000 171.2000 ;
	    RECT 14.2000 166.2000 14.5000 170.8000 ;
	    RECT 14.2000 165.8000 14.6000 166.2000 ;
	    RECT 14.2000 158.2000 14.5000 165.8000 ;
	    RECT 7.8000 157.8000 8.2000 158.2000 ;
	    RECT 14.2000 157.8000 14.6000 158.2000 ;
	    RECT 7.8000 155.2000 8.1000 157.8000 ;
	    RECT 2.2000 155.1000 2.6000 155.2000 ;
	    RECT 3.0000 155.1000 3.4000 155.2000 ;
	    RECT 2.2000 154.8000 3.4000 155.1000 ;
	    RECT 7.8000 154.8000 8.2000 155.2000 ;
	    RECT 7.8000 153.2000 8.1000 154.8000 ;
	    RECT 7.8000 152.8000 8.2000 153.2000 ;
         LAYER metal3 ;
	    RECT 11.8000 171.1000 12.2000 171.2000 ;
	    RECT 14.2000 171.1000 14.6000 171.2000 ;
	    RECT 11.8000 170.8000 14.6000 171.1000 ;
	    RECT 7.8000 158.1000 8.2000 158.2000 ;
	    RECT 14.2000 158.1000 14.6000 158.2000 ;
	    RECT 7.8000 157.8000 14.6000 158.1000 ;
	    RECT -2.6000 155.1000 -2.2000 155.2000 ;
	    RECT 3.0000 155.1000 3.4000 155.2000 ;
	    RECT 7.8000 155.1000 8.2000 155.2000 ;
	    RECT -2.6000 154.8000 8.2000 155.1000 ;
      END
   END target[8]
   PIN target[9]
      PORT
         LAYER metal1 ;
	    RECT 0.6000 172.4000 1.0000 173.2000 ;
	    RECT 4.6000 166.1000 5.0000 166.6000 ;
	    RECT 11.8000 166.4000 12.2000 167.2000 ;
	    RECT 5.4000 166.1000 5.8000 166.2000 ;
	    RECT 4.6000 165.8000 5.8000 166.1000 ;
	    RECT 4.6000 153.8000 5.0000 154.6000 ;
	    RECT 13.4000 147.8000 13.8000 148.6000 ;
	    RECT 5.4000 146.1000 5.8000 146.2000 ;
	    RECT 7.0000 146.1000 7.4000 146.6000 ;
	    RECT 5.4000 145.8000 7.4000 146.1000 ;
         LAYER metal2 ;
	    RECT 0.6000 173.8000 1.0000 174.2000 ;
	    RECT 0.6000 173.2000 0.9000 173.8000 ;
	    RECT 0.6000 172.8000 1.0000 173.2000 ;
	    RECT 5.4000 172.8000 5.8000 173.2000 ;
	    RECT 5.4000 166.2000 5.7000 172.8000 ;
	    RECT 11.8000 166.8000 12.2000 167.2000 ;
	    RECT 11.8000 166.2000 12.1000 166.8000 ;
	    RECT 5.4000 165.8000 5.8000 166.2000 ;
	    RECT 11.8000 165.8000 12.2000 166.2000 ;
	    RECT 4.6000 154.1000 5.0000 154.2000 ;
	    RECT 5.4000 154.1000 5.7000 165.8000 ;
	    RECT 4.6000 153.8000 5.7000 154.1000 ;
	    RECT 4.6000 147.1000 4.9000 153.8000 ;
	    RECT 5.4000 147.8000 5.8000 148.2000 ;
	    RECT 12.6000 148.1000 13.0000 148.2000 ;
	    RECT 13.4000 148.1000 13.8000 148.2000 ;
	    RECT 12.6000 147.8000 13.8000 148.1000 ;
	    RECT 5.4000 147.1000 5.7000 147.8000 ;
	    RECT 4.6000 146.8000 5.7000 147.1000 ;
	    RECT 5.4000 146.2000 5.7000 146.8000 ;
	    RECT 5.4000 145.8000 5.8000 146.2000 ;
         LAYER metal3 ;
	    RECT 0.6000 173.8000 1.0000 174.2000 ;
	    RECT -2.6000 173.1000 -2.2000 173.2000 ;
	    RECT 0.6000 173.1000 0.9000 173.8000 ;
	    RECT 5.4000 173.1000 5.8000 173.2000 ;
	    RECT -2.6000 172.8000 5.8000 173.1000 ;
	    RECT 5.4000 166.1000 5.8000 166.2000 ;
	    RECT 11.8000 166.1000 12.2000 166.2000 ;
	    RECT 5.4000 165.8000 12.2000 166.1000 ;
	    RECT 5.4000 148.1000 5.8000 148.2000 ;
	    RECT 12.6000 148.1000 13.0000 148.2000 ;
	    RECT 5.4000 147.8000 13.0000 148.1000 ;
      END
   END target[9]
   PIN target[10]
      PORT
         LAYER metal1 ;
	    RECT 12.6000 134.1000 13.0000 134.2000 ;
	    RECT 13.4000 134.1000 13.8000 134.2000 ;
	    RECT 12.6000 133.8000 13.8000 134.1000 ;
	    RECT 12.6000 133.4000 13.0000 133.8000 ;
	    RECT 13.4000 133.4000 13.8000 133.8000 ;
         LAYER metal2 ;
	    RECT 12.6000 134.1000 13.0000 134.2000 ;
	    RECT 13.4000 134.1000 13.8000 134.2000 ;
	    RECT 12.6000 133.8000 13.8000 134.1000 ;
         LAYER metal3 ;
	    RECT -2.6000 134.8000 -2.2000 135.2000 ;
	    RECT -2.6000 134.1000 -2.3000 134.8000 ;
	    RECT 13.4000 134.1000 13.8000 134.2000 ;
	    RECT -2.6000 133.8000 13.8000 134.1000 ;
      END
   END target[10]
   PIN target[11]
      PORT
         LAYER metal1 ;
	    RECT 12.6000 127.8000 13.0000 128.6000 ;
	    RECT 24.6000 127.8000 25.0000 128.6000 ;
	    RECT 5.0000 126.8000 5.8000 127.2000 ;
	    RECT 17.8000 127.1000 18.6000 127.2000 ;
	    RECT 19.0000 127.1000 19.4000 127.2000 ;
	    RECT 17.8000 126.8000 19.4000 127.1000 ;
         LAYER metal2 ;
	    RECT 12.6000 127.8000 13.0000 128.2000 ;
	    RECT 24.6000 127.8000 25.0000 128.2000 ;
	    RECT 12.6000 127.2000 12.9000 127.8000 ;
	    RECT 24.6000 127.2000 24.9000 127.8000 ;
	    RECT 5.4000 127.1000 5.8000 127.2000 ;
	    RECT 6.2000 127.1000 6.6000 127.2000 ;
	    RECT 5.4000 126.8000 6.6000 127.1000 ;
	    RECT 12.6000 126.8000 13.0000 127.2000 ;
	    RECT 18.2000 127.1000 18.6000 127.2000 ;
	    RECT 19.0000 127.1000 19.4000 127.2000 ;
	    RECT 18.2000 126.8000 19.4000 127.1000 ;
	    RECT 24.6000 126.8000 25.0000 127.2000 ;
	    RECT 5.4000 125.2000 5.7000 126.8000 ;
	    RECT 5.4000 124.8000 5.8000 125.2000 ;
         LAYER metal3 ;
	    RECT 6.2000 127.1000 6.6000 127.2000 ;
	    RECT 12.6000 127.1000 13.0000 127.2000 ;
	    RECT 18.2000 127.1000 18.6000 127.2000 ;
	    RECT 24.6000 127.1000 25.0000 127.2000 ;
	    RECT 6.2000 126.8000 25.0000 127.1000 ;
	    RECT -2.6000 125.1000 -2.2000 125.2000 ;
	    RECT 5.4000 125.1000 5.8000 125.2000 ;
	    RECT -2.6000 124.8000 5.8000 125.1000 ;
      END
   END target[11]
   PIN target[12]
      PORT
         LAYER metal1 ;
	    RECT 18.2000 174.8000 18.6000 175.6000 ;
	    RECT 17.4000 167.8000 17.8000 168.6000 ;
	    RECT 31.0000 167.8000 31.4000 168.6000 ;
	    RECT 19.8000 165.4000 20.2000 166.2000 ;
         LAYER metal2 ;
	    RECT 18.2000 182.8000 18.6000 183.2000 ;
	    RECT 18.2000 175.2000 18.5000 182.8000 ;
	    RECT 18.2000 174.8000 18.6000 175.2000 ;
	    RECT 18.2000 171.1000 18.5000 174.8000 ;
	    RECT 17.4000 170.8000 18.5000 171.1000 ;
	    RECT 17.4000 168.2000 17.7000 170.8000 ;
	    RECT 17.4000 167.8000 17.8000 168.2000 ;
	    RECT 31.0000 167.8000 31.4000 168.2000 ;
	    RECT 17.4000 166.2000 17.7000 167.8000 ;
	    RECT 31.0000 167.2000 31.3000 167.8000 ;
	    RECT 19.8000 166.8000 20.2000 167.2000 ;
	    RECT 31.0000 166.8000 31.4000 167.2000 ;
	    RECT 19.8000 166.2000 20.1000 166.8000 ;
	    RECT 17.4000 165.8000 17.8000 166.2000 ;
	    RECT 19.0000 166.1000 19.4000 166.2000 ;
	    RECT 19.8000 166.1000 20.2000 166.2000 ;
	    RECT 19.0000 165.8000 20.2000 166.1000 ;
         LAYER metal3 ;
	    RECT 19.8000 167.1000 20.2000 167.2000 ;
	    RECT 31.0000 167.1000 31.4000 167.2000 ;
	    RECT 19.8000 166.8000 31.4000 167.1000 ;
	    RECT 17.4000 166.1000 17.8000 166.2000 ;
	    RECT 19.0000 166.1000 19.4000 166.2000 ;
	    RECT 17.4000 165.8000 19.4000 166.1000 ;
      END
   END target[12]
   PIN target[13]
      PORT
         LAYER metal1 ;
	    RECT 20.6000 174.1000 21.0000 174.6000 ;
	    RECT 21.4000 174.1000 21.8000 174.2000 ;
	    RECT 20.6000 173.8000 21.8000 174.1000 ;
	    RECT 15.8000 172.4000 16.2000 173.2000 ;
	    RECT 25.4000 173.1000 25.8000 173.2000 ;
	    RECT 26.2000 173.1000 26.6000 173.2000 ;
	    RECT 25.4000 172.8000 26.6000 173.1000 ;
	    RECT 25.4000 172.4000 25.8000 172.8000 ;
	    RECT 26.2000 172.4000 26.6000 172.8000 ;
	    RECT 23.8000 167.8000 24.2000 168.6000 ;
	    RECT 22.2000 167.1000 22.6000 167.2000 ;
	    RECT 23.8000 167.1000 24.1000 167.8000 ;
	    RECT 22.2000 166.8000 24.1000 167.1000 ;
	    RECT 22.2000 166.4000 22.6000 166.8000 ;
         LAYER metal2 ;
	    RECT 22.2000 183.1000 22.6000 183.2000 ;
	    RECT 21.4000 182.8000 22.6000 183.1000 ;
	    RECT 21.4000 174.2000 21.7000 182.8000 ;
	    RECT 15.8000 173.8000 16.2000 174.2000 ;
	    RECT 21.4000 173.8000 21.8000 174.2000 ;
	    RECT 15.8000 173.2000 16.1000 173.8000 ;
	    RECT 21.4000 173.2000 21.7000 173.8000 ;
	    RECT 15.8000 172.8000 16.2000 173.2000 ;
	    RECT 21.4000 172.8000 21.8000 173.2000 ;
	    RECT 23.8000 172.8000 24.2000 173.2000 ;
	    RECT 24.6000 173.1000 25.0000 173.2000 ;
	    RECT 25.4000 173.1000 25.8000 173.2000 ;
	    RECT 24.6000 172.8000 25.8000 173.1000 ;
	    RECT 23.8000 168.2000 24.1000 172.8000 ;
	    RECT 23.8000 167.8000 24.2000 168.2000 ;
         LAYER metal3 ;
	    RECT 15.8000 173.8000 16.2000 174.2000 ;
	    RECT 15.8000 173.1000 16.1000 173.8000 ;
	    RECT 21.4000 173.1000 21.8000 173.2000 ;
	    RECT 23.8000 173.1000 24.2000 173.2000 ;
	    RECT 24.6000 173.1000 25.0000 173.2000 ;
	    RECT 15.8000 172.8000 25.0000 173.1000 ;
      END
   END target[13]
   PIN target[14]
      PORT
         LAYER metal1 ;
	    RECT 40.6000 173.4000 41.0000 174.2000 ;
	    RECT 45.4000 173.4000 45.8000 174.2000 ;
	    RECT 38.2000 167.8000 38.6000 168.6000 ;
	    RECT 44.6000 167.8000 45.0000 168.6000 ;
         LAYER metal2 ;
	    RECT 40.6000 182.8000 41.0000 183.2000 ;
	    RECT 40.6000 174.2000 40.9000 182.8000 ;
	    RECT 40.6000 173.8000 41.0000 174.2000 ;
	    RECT 45.4000 173.8000 45.8000 174.2000 ;
	    RECT 40.6000 173.2000 40.9000 173.8000 ;
	    RECT 45.4000 173.2000 45.7000 173.8000 ;
	    RECT 38.2000 172.8000 38.6000 173.2000 ;
	    RECT 40.6000 172.8000 41.0000 173.2000 ;
	    RECT 45.4000 172.8000 45.8000 173.2000 ;
	    RECT 38.2000 168.2000 38.5000 172.8000 ;
	    RECT 38.2000 167.8000 38.6000 168.2000 ;
	    RECT 44.6000 168.1000 45.0000 168.2000 ;
	    RECT 45.4000 168.1000 45.7000 172.8000 ;
	    RECT 44.6000 167.8000 45.7000 168.1000 ;
         LAYER metal3 ;
	    RECT 38.2000 173.1000 38.6000 173.2000 ;
	    RECT 40.6000 173.1000 41.0000 173.2000 ;
	    RECT 45.4000 173.1000 45.8000 173.2000 ;
	    RECT 38.2000 172.8000 45.8000 173.1000 ;
      END
   END target[14]
   PIN target[15]
      PORT
         LAYER metal1 ;
	    RECT 44.6000 174.8000 45.0000 175.2000 ;
	    RECT 44.6000 174.2000 44.9000 174.8000 ;
	    RECT 36.6000 173.4000 37.0000 174.2000 ;
	    RECT 44.6000 173.4000 45.0000 174.2000 ;
	    RECT 39.8000 166.8000 40.2000 167.6000 ;
	    RECT 50.2000 166.8000 50.6000 167.6000 ;
         LAYER metal2 ;
	    RECT 36.6000 182.8000 37.0000 183.2000 ;
	    RECT 36.6000 174.2000 36.9000 182.8000 ;
	    RECT 44.6000 174.8000 45.0000 175.2000 ;
	    RECT 44.6000 174.2000 44.9000 174.8000 ;
	    RECT 36.6000 174.1000 37.0000 174.2000 ;
	    RECT 37.4000 174.1000 37.8000 174.2000 ;
	    RECT 36.6000 173.8000 37.8000 174.1000 ;
	    RECT 39.8000 173.8000 40.2000 174.2000 ;
	    RECT 44.6000 173.8000 45.0000 174.2000 ;
	    RECT 50.2000 173.8000 50.6000 174.2000 ;
	    RECT 39.8000 167.2000 40.1000 173.8000 ;
	    RECT 50.2000 167.2000 50.5000 173.8000 ;
	    RECT 39.8000 166.8000 40.2000 167.2000 ;
	    RECT 50.2000 166.8000 50.6000 167.2000 ;
         LAYER metal3 ;
	    RECT 37.4000 174.1000 37.8000 174.2000 ;
	    RECT 39.8000 174.1000 40.2000 174.2000 ;
	    RECT 44.6000 174.1000 45.0000 174.2000 ;
	    RECT 50.2000 174.1000 50.6000 174.2000 ;
	    RECT 37.4000 173.8000 50.6000 174.1000 ;
      END
   END target[15]
   PIN nonce0[0]
      PORT
         LAYER metal1 ;
	    RECT 151.8000 175.9000 152.2000 179.9000 ;
	    RECT 151.8000 174.8000 152.1000 175.9000 ;
	    RECT 151.8000 171.1000 152.2000 174.8000 ;
         LAYER metal2 ;
	    RECT 152.6000 183.1000 153.0000 183.2000 ;
	    RECT 151.8000 182.8000 153.0000 183.1000 ;
	    RECT 151.8000 179.2000 152.1000 182.8000 ;
	    RECT 151.8000 178.8000 152.2000 179.2000 ;
      END
   END nonce0[0]
   PIN nonce0[1]
      PORT
         LAYER metal1 ;
	    RECT 156.6000 155.9000 157.0000 159.9000 ;
	    RECT 156.7000 154.8000 157.0000 155.9000 ;
	    RECT 156.6000 151.1000 157.0000 154.8000 ;
         LAYER metal2 ;
	    RECT 155.8000 182.8000 156.2000 183.2000 ;
	    RECT 155.8000 171.1000 156.1000 182.8000 ;
	    RECT 155.8000 170.8000 156.9000 171.1000 ;
	    RECT 156.6000 159.2000 156.9000 170.8000 ;
	    RECT 156.6000 158.8000 157.0000 159.2000 ;
      END
   END nonce0[1]
   PIN nonce0[2]
      PORT
         LAYER metal1 ;
	    RECT 76.6000 175.9000 77.0000 179.9000 ;
	    RECT 76.7000 174.8000 77.0000 175.9000 ;
	    RECT 76.6000 171.1000 77.0000 174.8000 ;
         LAYER metal2 ;
	    RECT 77.4000 183.1000 77.8000 183.2000 ;
	    RECT 76.6000 182.8000 77.8000 183.1000 ;
	    RECT 76.6000 179.2000 76.9000 182.8000 ;
	    RECT 76.6000 178.8000 77.0000 179.2000 ;
      END
   END nonce0[2]
   PIN nonce0[3]
      PORT
         LAYER metal1 ;
	    RECT 113.4000 175.9000 113.8000 179.9000 ;
	    RECT 113.5000 174.8000 113.8000 175.9000 ;
	    RECT 113.4000 171.1000 113.8000 174.8000 ;
         LAYER metal2 ;
	    RECT 112.6000 183.1000 113.0000 183.2000 ;
	    RECT 112.6000 182.8000 113.7000 183.1000 ;
	    RECT 113.4000 179.2000 113.7000 182.8000 ;
	    RECT 113.4000 178.8000 113.8000 179.2000 ;
      END
   END nonce0[3]
   PIN nonce0[4]
      PORT
         LAYER metal1 ;
	    RECT 79.0000 175.9000 79.4000 179.9000 ;
	    RECT 79.1000 174.8000 79.4000 175.9000 ;
	    RECT 79.0000 171.1000 79.4000 174.8000 ;
         LAYER metal2 ;
	    RECT 83.8000 182.8000 84.2000 183.2000 ;
	    RECT 83.8000 180.2000 84.1000 182.8000 ;
	    RECT 79.0000 179.8000 79.4000 180.2000 ;
	    RECT 83.8000 179.8000 84.2000 180.2000 ;
	    RECT 79.0000 179.2000 79.3000 179.8000 ;
	    RECT 79.0000 178.8000 79.4000 179.2000 ;
         LAYER metal3 ;
	    RECT 79.0000 180.1000 79.4000 180.2000 ;
	    RECT 83.8000 180.1000 84.2000 180.2000 ;
	    RECT 79.0000 179.8000 84.2000 180.1000 ;
      END
   END nonce0[4]
   PIN nonce0[5]
      PORT
         LAYER metal1 ;
	    RECT 74.2000 175.9000 74.6000 179.9000 ;
	    RECT 74.3000 174.8000 74.6000 175.9000 ;
	    RECT 74.2000 171.1000 74.6000 174.8000 ;
         LAYER metal2 ;
	    RECT 75.8000 182.8000 76.2000 183.2000 ;
	    RECT 75.8000 178.2000 76.1000 182.8000 ;
	    RECT 74.2000 177.8000 74.6000 178.2000 ;
	    RECT 75.8000 177.8000 76.2000 178.2000 ;
	    RECT 74.2000 177.2000 74.5000 177.8000 ;
	    RECT 74.2000 176.8000 74.6000 177.2000 ;
         LAYER metal3 ;
	    RECT 75.8000 178.1000 76.2000 178.2000 ;
	    RECT 74.2000 177.8000 76.2000 178.1000 ;
	    RECT 74.2000 177.2000 74.5000 177.8000 ;
	    RECT 74.2000 176.8000 74.6000 177.2000 ;
      END
   END nonce0[5]
   PIN nonce0[6]
      PORT
         LAYER metal1 ;
	    RECT 148.6000 175.9000 149.0000 179.9000 ;
	    RECT 148.7000 174.8000 149.0000 175.9000 ;
	    RECT 148.6000 171.1000 149.0000 174.8000 ;
         LAYER metal2 ;
	    RECT 147.8000 183.1000 148.2000 183.2000 ;
	    RECT 147.8000 182.8000 148.9000 183.1000 ;
	    RECT 148.6000 179.2000 148.9000 182.8000 ;
	    RECT 148.6000 178.8000 149.0000 179.2000 ;
      END
   END nonce0[6]
   PIN nonce0[7]
      PORT
         LAYER metal1 ;
	    RECT 51.0000 175.9000 51.4000 179.9000 ;
	    RECT 51.1000 174.8000 51.4000 175.9000 ;
	    RECT 51.0000 171.1000 51.4000 174.8000 ;
         LAYER metal2 ;
	    RECT 50.2000 183.1000 50.6000 183.2000 ;
	    RECT 50.2000 182.8000 51.3000 183.1000 ;
	    RECT 51.0000 179.2000 51.3000 182.8000 ;
	    RECT 51.0000 178.8000 51.4000 179.2000 ;
      END
   END nonce0[7]
   PIN nonce1[0]
      PORT
         LAYER metal1 ;
	    RECT 109.4000 179.1000 109.8000 179.9000 ;
	    RECT 110.2000 179.1000 110.6000 179.2000 ;
	    RECT 109.4000 178.8000 110.6000 179.1000 ;
	    RECT 109.4000 175.9000 109.8000 178.8000 ;
	    RECT 109.5000 174.8000 109.8000 175.9000 ;
	    RECT 109.4000 171.1000 109.8000 174.8000 ;
         LAYER metal2 ;
	    RECT 110.2000 182.8000 110.6000 183.2000 ;
	    RECT 110.2000 179.2000 110.5000 182.8000 ;
	    RECT 110.2000 178.8000 110.6000 179.2000 ;
      END
   END nonce1[0]
   PIN nonce1[1]
      PORT
         LAYER metal1 ;
	    RECT 44.6000 155.9000 45.0000 159.9000 ;
	    RECT 44.6000 154.8000 44.9000 155.9000 ;
	    RECT 44.6000 151.1000 45.0000 154.8000 ;
         LAYER metal2 ;
	    RECT 45.4000 182.8000 45.8000 183.2000 ;
	    RECT 45.4000 180.2000 45.7000 182.8000 ;
	    RECT 45.4000 179.8000 45.8000 180.2000 ;
	    RECT 44.6000 166.8000 45.0000 167.2000 ;
	    RECT 44.6000 159.2000 44.9000 166.8000 ;
	    RECT 44.6000 158.8000 45.0000 159.2000 ;
         LAYER metal3 ;
	    RECT 44.6000 180.1000 45.0000 180.2000 ;
	    RECT 45.4000 180.1000 45.8000 180.2000 ;
	    RECT 44.6000 179.8000 45.8000 180.1000 ;
	    RECT 44.6000 167.1000 45.0000 167.2000 ;
	    RECT 45.4000 167.1000 45.8000 167.2000 ;
	    RECT 44.6000 166.8000 45.8000 167.1000 ;
         LAYER metal4 ;
	    RECT 44.6000 180.1000 45.0000 180.2000 ;
	    RECT 44.6000 179.8000 45.7000 180.1000 ;
	    RECT 45.4000 167.2000 45.7000 179.8000 ;
	    RECT 45.4000 166.8000 45.8000 167.2000 ;
      END
   END nonce1[1]
   PIN nonce1[2]
      PORT
         LAYER metal1 ;
	    RECT 52.6000 6.2000 53.0000 9.9000 ;
	    RECT 52.7000 5.1000 53.0000 6.2000 ;
	    RECT 52.6000 1.1000 53.0000 5.1000 ;
         LAYER metal2 ;
	    RECT 52.6000 1.8000 53.0000 2.2000 ;
	    RECT 52.6000 1.2000 52.9000 1.8000 ;
	    RECT 52.6000 0.8000 53.0000 1.2000 ;
	    RECT 55.0000 0.8000 55.4000 1.2000 ;
	    RECT 55.0000 -1.8000 55.3000 0.8000 ;
	    RECT 55.0000 -2.2000 55.4000 -1.8000 ;
         LAYER metal3 ;
	    RECT 52.6000 1.1000 53.0000 1.2000 ;
	    RECT 55.0000 1.1000 55.4000 1.2000 ;
	    RECT 52.6000 0.8000 55.4000 1.1000 ;
      END
   END nonce1[2]
   PIN nonce1[3]
      PORT
         LAYER metal1 ;
	    RECT 97.4000 175.9000 97.8000 179.9000 ;
	    RECT 97.5000 174.8000 97.8000 175.9000 ;
	    RECT 97.4000 171.1000 97.8000 174.8000 ;
         LAYER metal2 ;
	    RECT 96.6000 183.1000 97.0000 183.2000 ;
	    RECT 96.6000 182.8000 97.7000 183.1000 ;
	    RECT 97.4000 179.2000 97.7000 182.8000 ;
	    RECT 97.4000 178.8000 97.8000 179.2000 ;
      END
   END nonce1[3]
   PIN nonce1[4]
      PORT
         LAYER metal1 ;
	    RECT 171.0000 15.9000 171.4000 19.9000 ;
	    RECT 171.0000 14.8000 171.3000 15.9000 ;
	    RECT 171.0000 11.1000 171.4000 14.8000 ;
         LAYER metal2 ;
	    RECT 171.0000 11.8000 171.4000 12.2000 ;
	    RECT 171.0000 -1.9000 171.3000 11.8000 ;
	    RECT 171.8000 -1.9000 172.2000 -1.8000 ;
	    RECT 171.0000 -2.2000 172.2000 -1.9000 ;
      END
   END nonce1[4]
   PIN nonce1[5]
      PORT
         LAYER metal1 ;
	    RECT 269.4000 175.9000 269.8000 179.9000 ;
	    RECT 269.5000 174.8000 269.8000 175.9000 ;
	    RECT 269.4000 171.1000 269.8000 174.8000 ;
         LAYER metal2 ;
	    RECT 268.6000 183.1000 269.0000 183.2000 ;
	    RECT 268.6000 182.8000 269.7000 183.1000 ;
	    RECT 269.4000 179.2000 269.7000 182.8000 ;
	    RECT 269.4000 178.8000 269.8000 179.2000 ;
      END
   END nonce1[5]
   PIN nonce1[6]
      PORT
         LAYER metal1 ;
	    RECT 189.4000 175.9000 189.8000 179.9000 ;
	    RECT 189.5000 174.8000 189.8000 175.9000 ;
	    RECT 189.4000 171.1000 189.8000 174.8000 ;
         LAYER metal2 ;
	    RECT 188.6000 183.1000 189.0000 183.2000 ;
	    RECT 188.6000 182.8000 189.7000 183.1000 ;
	    RECT 189.4000 179.2000 189.7000 182.8000 ;
	    RECT 189.4000 178.8000 189.8000 179.2000 ;
      END
   END nonce1[6]
   PIN nonce1[7]
      PORT
         LAYER metal1 ;
	    RECT 266.2000 6.2000 266.6000 9.9000 ;
	    RECT 266.2000 5.1000 266.5000 6.2000 ;
	    RECT 266.2000 1.1000 266.6000 5.1000 ;
         LAYER metal2 ;
	    RECT 266.2000 1.8000 266.6000 2.2000 ;
	    RECT 266.2000 -1.9000 266.5000 1.8000 ;
	    RECT 267.0000 -1.9000 267.4000 -1.8000 ;
	    RECT 266.2000 -2.2000 267.4000 -1.9000 ;
      END
   END nonce1[7]
   PIN nonce2[0]
      PORT
         LAYER metal1 ;
	    RECT 151.0000 175.9000 151.4000 179.9000 ;
	    RECT 151.1000 174.8000 151.4000 175.9000 ;
	    RECT 151.0000 171.1000 151.4000 174.8000 ;
         LAYER metal2 ;
	    RECT 150.2000 183.1000 150.6000 183.2000 ;
	    RECT 150.2000 182.8000 151.3000 183.1000 ;
	    RECT 151.0000 179.2000 151.3000 182.8000 ;
	    RECT 151.0000 178.8000 151.4000 179.2000 ;
      END
   END nonce2[0]
   PIN nonce2[1]
      PORT
         LAYER metal1 ;
	    RECT 199.8000 6.2000 200.2000 9.9000 ;
	    RECT 199.9000 5.1000 200.2000 6.2000 ;
	    RECT 199.8000 1.1000 200.2000 5.1000 ;
         LAYER metal2 ;
	    RECT 199.8000 1.8000 200.2000 2.2000 ;
	    RECT 199.0000 -1.9000 199.4000 -1.8000 ;
	    RECT 199.8000 -1.9000 200.1000 1.8000 ;
	    RECT 199.0000 -2.2000 200.1000 -1.9000 ;
      END
   END nonce2[1]
   PIN nonce2[2]
      PORT
         LAYER metal1 ;
	    RECT 169.4000 175.9000 169.8000 179.9000 ;
	    RECT 169.4000 174.8000 169.7000 175.9000 ;
	    RECT 169.4000 171.1000 169.8000 174.8000 ;
         LAYER metal2 ;
	    RECT 170.2000 183.1000 170.6000 183.2000 ;
	    RECT 169.4000 182.8000 170.6000 183.1000 ;
	    RECT 169.4000 179.2000 169.7000 182.8000 ;
	    RECT 169.4000 178.8000 169.8000 179.2000 ;
      END
   END nonce2[2]
   PIN nonce2[3]
      PORT
         LAYER metal1 ;
	    RECT 123.8000 175.9000 124.2000 179.9000 ;
	    RECT 123.8000 174.8000 124.1000 175.9000 ;
	    RECT 123.8000 171.1000 124.2000 174.8000 ;
         LAYER metal2 ;
	    RECT 124.6000 183.1000 125.0000 183.2000 ;
	    RECT 123.8000 182.8000 125.0000 183.1000 ;
	    RECT 123.8000 179.2000 124.1000 182.8000 ;
	    RECT 123.8000 178.8000 124.2000 179.2000 ;
      END
   END nonce2[3]
   PIN nonce2[4]
      PORT
         LAYER metal1 ;
	    RECT 131.8000 175.9000 132.2000 179.9000 ;
	    RECT 131.9000 174.8000 132.2000 175.9000 ;
	    RECT 131.8000 171.1000 132.2000 174.8000 ;
         LAYER metal2 ;
	    RECT 131.0000 183.1000 131.4000 183.2000 ;
	    RECT 131.0000 182.8000 132.1000 183.1000 ;
	    RECT 131.8000 179.2000 132.1000 182.8000 ;
	    RECT 131.8000 178.8000 132.2000 179.2000 ;
      END
   END nonce2[4]
   PIN nonce2[5]
      PORT
         LAYER metal1 ;
	    RECT 0.6000 6.2000 1.0000 9.9000 ;
	    RECT 0.6000 5.1000 0.9000 6.2000 ;
	    RECT 0.6000 1.1000 1.0000 5.1000 ;
         LAYER metal2 ;
	    RECT 0.6000 7.8000 1.0000 8.2000 ;
	    RECT 0.6000 7.2000 0.9000 7.8000 ;
	    RECT 0.6000 6.8000 1.0000 7.2000 ;
         LAYER metal3 ;
	    RECT 0.6000 7.8000 1.0000 8.2000 ;
	    RECT -2.6000 7.1000 -2.2000 7.2000 ;
	    RECT 0.6000 7.1000 0.9000 7.8000 ;
	    RECT -2.6000 6.8000 0.9000 7.1000 ;
      END
   END nonce2[5]
   PIN nonce2[6]
      PORT
         LAYER metal1 ;
	    RECT 95.0000 175.9000 95.4000 179.9000 ;
	    RECT 95.1000 174.8000 95.4000 175.9000 ;
	    RECT 95.0000 171.1000 95.4000 174.8000 ;
         LAYER metal2 ;
	    RECT 95.0000 182.8000 95.4000 183.2000 ;
	    RECT 95.0000 179.2000 95.3000 182.8000 ;
	    RECT 95.0000 178.8000 95.4000 179.2000 ;
      END
   END nonce2[6]
   PIN nonce2[7]
      PORT
         LAYER metal1 ;
	    RECT 146.2000 175.9000 146.6000 179.9000 ;
	    RECT 146.3000 174.8000 146.6000 175.9000 ;
	    RECT 146.2000 171.1000 146.6000 174.8000 ;
         LAYER metal2 ;
	    RECT 145.4000 183.1000 145.8000 183.2000 ;
	    RECT 145.4000 182.8000 146.5000 183.1000 ;
	    RECT 146.2000 179.2000 146.5000 182.8000 ;
	    RECT 146.2000 178.8000 146.6000 179.2000 ;
      END
   END nonce2[7]
   PIN nonce3[0]
      PORT
         LAYER metal1 ;
	    RECT 143.8000 175.9000 144.2000 179.9000 ;
	    RECT 143.9000 174.8000 144.2000 175.9000 ;
	    RECT 143.8000 171.1000 144.2000 174.8000 ;
         LAYER metal2 ;
	    RECT 143.0000 183.1000 143.4000 183.2000 ;
	    RECT 143.0000 182.8000 144.1000 183.1000 ;
	    RECT 143.8000 179.2000 144.1000 182.8000 ;
	    RECT 143.8000 178.8000 144.2000 179.2000 ;
      END
   END nonce3[0]
   PIN nonce3[1]
      PORT
         LAYER metal1 ;
	    RECT 76.6000 155.9000 77.0000 159.9000 ;
	    RECT 76.7000 154.8000 77.0000 155.9000 ;
	    RECT 76.6000 151.1000 77.0000 154.8000 ;
         LAYER metal2 ;
	    RECT 79.0000 183.1000 79.4000 183.2000 ;
	    RECT 78.2000 182.8000 79.4000 183.1000 ;
	    RECT 78.2000 178.2000 78.5000 182.8000 ;
	    RECT 76.6000 177.8000 77.0000 178.2000 ;
	    RECT 78.2000 177.8000 78.6000 178.2000 ;
	    RECT 76.6000 159.2000 76.9000 177.8000 ;
	    RECT 76.6000 158.8000 77.0000 159.2000 ;
         LAYER metal3 ;
	    RECT 76.6000 178.1000 77.0000 178.2000 ;
	    RECT 78.2000 178.1000 78.6000 178.2000 ;
	    RECT 76.6000 177.8000 78.6000 178.1000 ;
      END
   END nonce3[1]
   PIN nonce3[2]
      PORT
         LAYER metal1 ;
	    RECT 168.6000 175.9000 169.0000 179.9000 ;
	    RECT 168.7000 174.8000 169.0000 175.9000 ;
	    RECT 168.6000 171.1000 169.0000 174.8000 ;
         LAYER metal2 ;
	    RECT 167.8000 183.1000 168.2000 183.2000 ;
	    RECT 167.8000 182.8000 168.9000 183.1000 ;
	    RECT 168.6000 179.2000 168.9000 182.8000 ;
	    RECT 168.6000 178.8000 169.0000 179.2000 ;
      END
   END nonce3[2]
   PIN nonce3[3]
      PORT
         LAYER metal1 ;
	    RECT 182.2000 6.2000 182.6000 9.9000 ;
	    RECT 182.2000 5.1000 182.5000 6.2000 ;
	    RECT 182.2000 1.1000 182.6000 5.1000 ;
         LAYER metal2 ;
	    RECT 182.2000 1.8000 182.6000 2.2000 ;
	    RECT 182.2000 -1.8000 182.5000 1.8000 ;
	    RECT 182.2000 -2.2000 182.6000 -1.8000 ;
      END
   END nonce3[3]
   PIN nonce3[4]
      PORT
         LAYER metal1 ;
	    RECT 3.0000 6.2000 3.4000 9.9000 ;
	    RECT 3.0000 5.1000 3.3000 6.2000 ;
	    RECT 3.0000 1.1000 3.4000 5.1000 ;
         LAYER metal2 ;
	    RECT 3.0000 6.8000 3.4000 7.2000 ;
	    RECT 3.0000 5.2000 3.3000 6.8000 ;
	    RECT 3.0000 4.8000 3.4000 5.2000 ;
         LAYER metal3 ;
	    RECT -2.6000 5.1000 -2.2000 5.2000 ;
	    RECT 3.0000 5.1000 3.4000 5.2000 ;
	    RECT -2.6000 4.8000 3.4000 5.1000 ;
      END
   END nonce3[4]
   PIN nonce3[5]
      PORT
         LAYER metal1 ;
	    RECT 173.4000 175.9000 173.8000 179.9000 ;
	    RECT 173.5000 174.8000 173.8000 175.9000 ;
	    RECT 173.4000 171.1000 173.8000 174.8000 ;
         LAYER metal2 ;
	    RECT 178.2000 182.8000 178.6000 183.2000 ;
	    RECT 178.2000 180.2000 178.5000 182.8000 ;
	    RECT 173.4000 179.8000 173.8000 180.2000 ;
	    RECT 178.2000 179.8000 178.6000 180.2000 ;
	    RECT 173.4000 179.2000 173.7000 179.8000 ;
	    RECT 173.4000 178.8000 173.8000 179.2000 ;
         LAYER metal3 ;
	    RECT 173.4000 180.1000 173.8000 180.2000 ;
	    RECT 178.2000 180.1000 178.6000 180.2000 ;
	    RECT 173.4000 179.8000 178.6000 180.1000 ;
      END
   END nonce3[5]
   PIN nonce3[6]
      PORT
         LAYER metal1 ;
	    RECT 36.6000 6.2000 37.0000 9.9000 ;
	    RECT 36.7000 5.1000 37.0000 6.2000 ;
	    RECT 36.6000 1.1000 37.0000 5.1000 ;
         LAYER metal2 ;
	    RECT 36.6000 1.8000 37.0000 2.2000 ;
	    RECT 35.8000 -1.9000 36.2000 -1.8000 ;
	    RECT 36.6000 -1.9000 36.9000 1.8000 ;
	    RECT 35.8000 -2.2000 36.9000 -1.9000 ;
      END
   END nonce3[6]
   PIN nonce3[7]
      PORT
         LAYER metal1 ;
	    RECT 19.0000 6.2000 19.4000 9.9000 ;
	    RECT 19.0000 5.1000 19.3000 6.2000 ;
	    RECT 19.0000 1.1000 19.4000 5.1000 ;
         LAYER metal2 ;
	    RECT 19.0000 1.8000 19.4000 2.2000 ;
	    RECT 19.0000 -1.9000 19.3000 1.8000 ;
	    RECT 19.8000 -1.9000 20.2000 -1.8000 ;
	    RECT 19.0000 -2.2000 20.2000 -1.9000 ;
      END
   END nonce3[7]
   PIN finish
      PORT
         LAYER metal1 ;
	    RECT 121.4000 155.9000 121.8000 159.9000 ;
	    RECT 121.4000 154.8000 121.7000 155.9000 ;
	    RECT 121.4000 151.1000 121.8000 154.8000 ;
         LAYER metal2 ;
	    RECT 122.2000 182.8000 122.6000 183.2000 ;
	    RECT 122.2000 168.1000 122.5000 182.8000 ;
	    RECT 121.4000 167.8000 122.5000 168.1000 ;
	    RECT 121.4000 159.2000 121.7000 167.8000 ;
	    RECT 121.4000 158.8000 121.8000 159.2000 ;
      END
   END finish
   OBS
         LAYER metal1 ;
	    RECT 0.6000 176.1000 1.0000 176.2000 ;
	    RECT 1.4000 176.1000 1.8000 179.9000 ;
	    RECT 0.6000 175.8000 1.8000 176.1000 ;
	    RECT 3.5000 175.9000 4.5000 179.9000 ;
	    RECT 1.4000 174.1000 1.8000 175.8000 ;
	    RECT 3.8000 174.2000 4.1000 175.9000 ;
	    RECT 6.2000 175.8000 6.6000 176.6000 ;
	    RECT 2.2000 174.1000 2.6000 174.2000 ;
	    RECT 3.8000 174.1000 4.2000 174.2000 ;
	    RECT 1.4000 173.8000 3.0000 174.1000 ;
	    RECT 3.8000 173.8000 5.0000 174.1000 ;
	    RECT 5.4000 173.8000 5.8000 174.6000 ;
	    RECT 1.4000 171.1000 1.8000 173.8000 ;
	    RECT 2.6000 173.6000 3.0000 173.8000 ;
	    RECT 2.3000 173.1000 4.1000 173.3000 ;
	    RECT 4.7000 173.1000 5.0000 173.8000 ;
	    RECT 7.0000 173.1000 7.4000 179.9000 ;
	    RECT 8.6000 175.8000 9.0000 176.6000 ;
	    RECT 9.4000 173.1000 9.8000 179.9000 ;
	    RECT 10.2000 176.8000 10.6000 177.2000 ;
	    RECT 10.2000 176.1000 10.5000 176.8000 ;
	    RECT 11.0000 176.1000 11.4000 179.9000 ;
	    RECT 10.2000 175.8000 11.4000 176.1000 ;
	    RECT 2.2000 173.0000 4.2000 173.1000 ;
	    RECT 2.2000 171.1000 2.6000 173.0000 ;
	    RECT 3.8000 171.4000 4.2000 173.0000 ;
	    RECT 4.6000 171.7000 5.0000 173.1000 ;
	    RECT 5.4000 171.4000 5.8000 173.1000 ;
	    RECT 3.8000 171.1000 5.8000 171.4000 ;
	    RECT 6.5000 172.8000 7.4000 173.1000 ;
	    RECT 8.9000 172.8000 9.8000 173.1000 ;
	    RECT 6.5000 172.2000 6.9000 172.8000 ;
	    RECT 8.9000 172.2000 9.3000 172.8000 ;
	    RECT 6.5000 171.8000 7.4000 172.2000 ;
	    RECT 8.6000 171.8000 9.3000 172.2000 ;
	    RECT 6.5000 171.1000 6.9000 171.8000 ;
	    RECT 8.9000 171.1000 9.3000 171.8000 ;
	    RECT 11.0000 171.1000 11.4000 175.8000 ;
	    RECT 13.4000 173.1000 13.8000 179.9000 ;
	    RECT 14.2000 176.1000 14.6000 176.6000 ;
	    RECT 15.0000 176.1000 15.4000 179.9000 ;
	    RECT 14.2000 175.8000 15.4000 176.1000 ;
	    RECT 13.4000 172.8000 14.3000 173.1000 ;
	    RECT 13.9000 172.2000 14.3000 172.8000 ;
	    RECT 13.9000 171.8000 14.6000 172.2000 ;
	    RECT 13.9000 171.1000 14.3000 171.8000 ;
	    RECT 15.0000 171.1000 15.4000 175.8000 ;
	    RECT 17.4000 174.1000 17.8000 179.9000 ;
	    RECT 18.2000 179.6000 20.2000 179.9000 ;
	    RECT 18.2000 175.9000 18.6000 179.6000 ;
	    RECT 19.0000 175.9000 19.4000 179.3000 ;
	    RECT 19.8000 176.2000 20.2000 179.6000 ;
	    RECT 21.4000 176.2000 21.8000 179.9000 ;
	    RECT 19.8000 175.9000 21.8000 176.2000 ;
	    RECT 19.1000 175.6000 19.4000 175.9000 ;
	    RECT 19.1000 175.3000 20.1000 175.6000 ;
	    RECT 19.8000 175.2000 20.1000 175.3000 ;
	    RECT 21.0000 175.2000 21.4000 175.4000 ;
	    RECT 19.8000 174.8000 20.2000 175.2000 ;
	    RECT 21.0000 175.1000 21.8000 175.2000 ;
	    RECT 22.2000 175.1000 22.6000 179.9000 ;
	    RECT 24.1000 176.3000 24.5000 179.9000 ;
	    RECT 24.1000 175.9000 25.0000 176.3000 ;
	    RECT 27.0000 176.1000 27.4000 179.9000 ;
	    RECT 27.8000 176.1000 28.2000 176.6000 ;
	    RECT 23.8000 175.1000 24.2000 175.6000 ;
	    RECT 21.0000 174.9000 24.2000 175.1000 ;
	    RECT 21.4000 174.8000 24.2000 174.9000 ;
	    RECT 19.1000 174.4000 19.5000 174.8000 ;
	    RECT 19.1000 174.2000 19.4000 174.4000 ;
	    RECT 19.0000 174.1000 19.4000 174.2000 ;
	    RECT 17.4000 173.8000 19.4000 174.1000 ;
	    RECT 17.4000 171.1000 17.8000 173.8000 ;
	    RECT 19.8000 173.1000 20.1000 174.8000 ;
	    RECT 19.5000 171.1000 20.3000 173.1000 ;
	    RECT 22.2000 171.1000 22.6000 174.8000 ;
	    RECT 24.6000 174.2000 24.9000 175.9000 ;
	    RECT 27.0000 175.8000 28.2000 176.1000 ;
	    RECT 24.6000 174.1000 25.0000 174.2000 ;
	    RECT 25.4000 174.1000 25.8000 174.2000 ;
	    RECT 24.6000 173.8000 25.8000 174.1000 ;
	    RECT 24.6000 172.1000 24.9000 173.8000 ;
	    RECT 24.6000 171.1000 25.0000 172.1000 ;
	    RECT 27.0000 171.1000 27.4000 175.8000 ;
	    RECT 28.6000 173.1000 29.0000 179.9000 ;
	    RECT 30.2000 175.6000 30.6000 179.9000 ;
	    RECT 32.3000 176.2000 32.7000 179.9000 ;
	    RECT 32.3000 175.9000 33.0000 176.2000 ;
	    RECT 30.2000 175.4000 32.2000 175.6000 ;
	    RECT 30.2000 175.3000 32.3000 175.4000 ;
	    RECT 31.9000 175.0000 32.3000 175.3000 ;
	    RECT 32.7000 175.2000 33.0000 175.9000 ;
	    RECT 31.2000 174.2000 31.6000 174.6000 ;
	    RECT 31.0000 173.8000 31.5000 174.2000 ;
	    RECT 32.0000 173.5000 32.3000 175.0000 ;
	    RECT 32.6000 174.8000 33.0000 175.2000 ;
	    RECT 31.1000 173.2000 32.3000 173.5000 ;
	    RECT 28.1000 172.8000 29.0000 173.1000 ;
	    RECT 28.1000 172.2000 28.5000 172.8000 ;
	    RECT 30.2000 172.4000 30.6000 173.2000 ;
	    RECT 27.8000 171.8000 28.5000 172.2000 ;
	    RECT 31.1000 172.1000 31.4000 173.2000 ;
	    RECT 32.7000 173.1000 33.0000 174.8000 ;
	    RECT 28.1000 171.1000 28.5000 171.8000 ;
	    RECT 31.0000 171.1000 31.4000 172.1000 ;
	    RECT 32.6000 171.1000 33.0000 173.1000 ;
	    RECT 34.2000 176.1000 34.6000 179.9000 ;
	    RECT 35.0000 176.1000 35.4000 176.6000 ;
	    RECT 34.2000 175.8000 35.4000 176.1000 ;
	    RECT 34.2000 171.1000 34.6000 175.8000 ;
	    RECT 35.8000 173.1000 36.2000 179.9000 ;
	    RECT 35.3000 172.8000 36.2000 173.1000 ;
	    RECT 38.2000 176.1000 38.6000 179.9000 ;
	    RECT 39.0000 176.1000 39.4000 176.6000 ;
	    RECT 38.2000 175.8000 39.4000 176.1000 ;
	    RECT 35.3000 172.2000 35.7000 172.8000 ;
	    RECT 35.0000 171.8000 35.7000 172.2000 ;
	    RECT 35.3000 171.1000 35.7000 171.8000 ;
	    RECT 38.2000 171.1000 38.6000 175.8000 ;
	    RECT 39.8000 173.1000 40.2000 179.9000 ;
	    RECT 39.3000 172.8000 40.2000 173.1000 ;
	    RECT 42.2000 176.1000 42.6000 179.9000 ;
	    RECT 43.0000 176.1000 43.4000 176.6000 ;
	    RECT 42.2000 175.8000 43.4000 176.1000 ;
	    RECT 39.3000 172.2000 39.7000 172.8000 ;
	    RECT 39.0000 171.8000 39.7000 172.2000 ;
	    RECT 39.3000 171.1000 39.7000 171.8000 ;
	    RECT 42.2000 171.1000 42.6000 175.8000 ;
	    RECT 43.8000 173.1000 44.2000 179.9000 ;
	    RECT 43.3000 172.8000 44.2000 173.1000 ;
	    RECT 46.2000 173.1000 46.6000 179.9000 ;
	    RECT 47.0000 176.1000 47.4000 176.6000 ;
	    RECT 47.8000 176.1000 48.2000 179.9000 ;
	    RECT 47.0000 175.8000 48.2000 176.1000 ;
	    RECT 49.4000 176.2000 49.8000 179.9000 ;
	    RECT 49.4000 175.9000 50.5000 176.2000 ;
	    RECT 46.2000 172.8000 47.1000 173.1000 ;
	    RECT 43.3000 172.2000 43.7000 172.8000 ;
	    RECT 46.7000 172.2000 47.1000 172.8000 ;
	    RECT 43.3000 171.8000 44.2000 172.2000 ;
	    RECT 46.7000 171.8000 47.4000 172.2000 ;
	    RECT 43.3000 171.1000 43.7000 171.8000 ;
	    RECT 46.7000 171.1000 47.1000 171.8000 ;
	    RECT 47.8000 171.1000 48.2000 175.8000 ;
	    RECT 50.2000 175.6000 50.5000 175.9000 ;
	    RECT 51.8000 175.6000 52.2000 179.9000 ;
	    RECT 53.9000 177.9000 54.5000 179.9000 ;
	    RECT 56.2000 177.9000 56.6000 179.9000 ;
	    RECT 58.4000 178.2000 58.8000 179.9000 ;
	    RECT 58.4000 177.9000 59.4000 178.2000 ;
	    RECT 54.2000 177.5000 54.6000 177.9000 ;
	    RECT 56.3000 177.6000 56.6000 177.9000 ;
	    RECT 55.9000 177.3000 57.7000 177.6000 ;
	    RECT 59.0000 177.5000 59.4000 177.9000 ;
	    RECT 55.9000 177.2000 56.3000 177.3000 ;
	    RECT 57.3000 177.2000 57.7000 177.3000 ;
	    RECT 53.8000 176.6000 54.5000 177.0000 ;
	    RECT 54.2000 176.1000 54.5000 176.6000 ;
	    RECT 55.3000 176.5000 56.4000 176.8000 ;
	    RECT 55.3000 176.4000 55.7000 176.5000 ;
	    RECT 54.2000 175.8000 55.4000 176.1000 ;
	    RECT 50.2000 175.2000 50.8000 175.6000 ;
	    RECT 51.8000 175.3000 53.9000 175.6000 ;
	    RECT 49.4000 174.4000 49.8000 175.2000 ;
	    RECT 50.2000 173.7000 50.5000 175.2000 ;
	    RECT 49.4000 173.4000 50.5000 173.7000 ;
	    RECT 51.8000 173.6000 52.2000 175.3000 ;
	    RECT 53.5000 175.2000 53.9000 175.3000 ;
	    RECT 52.7000 174.9000 53.1000 175.0000 ;
	    RECT 52.7000 174.6000 54.6000 174.9000 ;
	    RECT 54.2000 174.5000 54.6000 174.6000 ;
	    RECT 55.1000 174.2000 55.4000 175.8000 ;
	    RECT 56.1000 175.9000 56.4000 176.5000 ;
	    RECT 56.7000 176.5000 57.1000 176.6000 ;
	    RECT 59.0000 176.5000 59.4000 176.6000 ;
	    RECT 56.7000 176.2000 59.4000 176.5000 ;
	    RECT 56.1000 175.7000 58.5000 175.9000 ;
	    RECT 60.6000 175.7000 61.0000 179.9000 ;
	    RECT 56.1000 175.6000 61.0000 175.7000 ;
	    RECT 58.1000 175.5000 61.0000 175.6000 ;
	    RECT 58.2000 175.4000 61.0000 175.5000 ;
	    RECT 63.0000 175.7000 63.4000 179.9000 ;
	    RECT 65.2000 178.2000 65.6000 179.9000 ;
	    RECT 64.6000 177.9000 65.6000 178.2000 ;
	    RECT 67.4000 177.9000 67.8000 179.9000 ;
	    RECT 69.5000 177.9000 70.1000 179.9000 ;
	    RECT 64.6000 177.5000 65.0000 177.9000 ;
	    RECT 67.4000 177.6000 67.7000 177.9000 ;
	    RECT 66.3000 177.3000 68.1000 177.6000 ;
	    RECT 69.4000 177.5000 69.8000 177.9000 ;
	    RECT 66.3000 177.2000 66.7000 177.3000 ;
	    RECT 67.7000 177.2000 68.1000 177.3000 ;
	    RECT 64.6000 176.5000 65.0000 176.6000 ;
	    RECT 66.9000 176.5000 67.3000 176.6000 ;
	    RECT 64.6000 176.2000 67.3000 176.5000 ;
	    RECT 67.6000 176.5000 68.7000 176.8000 ;
	    RECT 67.6000 175.9000 67.9000 176.5000 ;
	    RECT 68.3000 176.4000 68.7000 176.5000 ;
	    RECT 69.5000 176.6000 70.2000 177.0000 ;
	    RECT 69.5000 176.1000 69.8000 176.6000 ;
	    RECT 65.5000 175.7000 67.9000 175.9000 ;
	    RECT 63.0000 175.6000 67.9000 175.7000 ;
	    RECT 68.6000 175.8000 69.8000 176.1000 ;
	    RECT 63.0000 175.5000 65.9000 175.6000 ;
	    RECT 63.0000 175.4000 65.8000 175.5000 ;
	    RECT 57.4000 175.1000 57.8000 175.2000 ;
	    RECT 66.2000 175.1000 66.6000 175.2000 ;
	    RECT 67.8000 175.1000 68.2000 175.2000 ;
	    RECT 57.4000 174.8000 59.9000 175.1000 ;
	    RECT 58.2000 174.7000 58.6000 174.8000 ;
	    RECT 59.5000 174.7000 59.9000 174.8000 ;
	    RECT 64.1000 174.8000 68.2000 175.1000 ;
	    RECT 64.1000 174.7000 64.5000 174.8000 ;
	    RECT 58.7000 174.2000 59.1000 174.3000 ;
	    RECT 64.9000 174.2000 65.3000 174.3000 ;
	    RECT 68.6000 174.2000 68.9000 175.8000 ;
	    RECT 71.8000 175.6000 72.2000 179.9000 ;
	    RECT 72.6000 176.2000 73.0000 179.9000 ;
	    RECT 75.0000 176.2000 75.4000 179.9000 ;
	    RECT 77.4000 176.2000 77.8000 179.9000 ;
	    RECT 72.6000 175.9000 73.7000 176.2000 ;
	    RECT 75.0000 175.9000 76.1000 176.2000 ;
	    RECT 77.4000 175.9000 78.5000 176.2000 ;
	    RECT 70.1000 175.3000 72.2000 175.6000 ;
	    RECT 70.1000 175.2000 70.5000 175.3000 ;
	    RECT 71.8000 175.1000 72.2000 175.3000 ;
	    RECT 73.4000 175.6000 73.7000 175.9000 ;
	    RECT 75.8000 175.6000 76.1000 175.9000 ;
	    RECT 78.2000 175.6000 78.5000 175.9000 ;
	    RECT 79.8000 175.7000 80.2000 179.9000 ;
	    RECT 82.0000 178.2000 82.4000 179.9000 ;
	    RECT 81.4000 177.9000 82.4000 178.2000 ;
	    RECT 84.2000 177.9000 84.6000 179.9000 ;
	    RECT 86.3000 177.9000 86.9000 179.9000 ;
	    RECT 81.4000 177.5000 81.8000 177.9000 ;
	    RECT 84.2000 177.6000 84.5000 177.9000 ;
	    RECT 83.1000 177.3000 84.9000 177.6000 ;
	    RECT 86.2000 177.5000 86.6000 177.9000 ;
	    RECT 83.1000 177.2000 83.5000 177.3000 ;
	    RECT 84.5000 177.2000 84.9000 177.3000 ;
	    RECT 81.4000 176.5000 81.8000 176.6000 ;
	    RECT 83.7000 176.5000 84.1000 176.6000 ;
	    RECT 81.4000 176.2000 84.1000 176.5000 ;
	    RECT 84.4000 176.5000 85.5000 176.8000 ;
	    RECT 84.4000 175.9000 84.7000 176.5000 ;
	    RECT 85.1000 176.4000 85.5000 176.5000 ;
	    RECT 86.3000 176.6000 87.0000 177.0000 ;
	    RECT 86.3000 176.1000 86.6000 176.6000 ;
	    RECT 82.3000 175.7000 84.7000 175.9000 ;
	    RECT 79.8000 175.6000 84.7000 175.7000 ;
	    RECT 85.4000 175.8000 86.6000 176.1000 ;
	    RECT 88.6000 176.1000 89.0000 179.9000 ;
	    RECT 89.4000 176.8000 89.8000 177.2000 ;
	    RECT 89.4000 176.1000 89.7000 176.8000 ;
	    RECT 88.6000 175.8000 89.7000 176.1000 ;
	    RECT 73.4000 175.2000 74.0000 175.6000 ;
	    RECT 75.8000 175.2000 76.4000 175.6000 ;
	    RECT 78.2000 175.2000 78.8000 175.6000 ;
	    RECT 79.8000 175.5000 82.7000 175.6000 ;
	    RECT 79.8000 175.4000 82.6000 175.5000 ;
	    RECT 72.6000 175.1000 73.0000 175.2000 ;
	    RECT 70.9000 174.9000 71.3000 175.0000 ;
	    RECT 69.4000 174.6000 71.3000 174.9000 ;
	    RECT 71.8000 174.8000 73.0000 175.1000 ;
	    RECT 69.4000 174.5000 69.8000 174.6000 ;
	    RECT 55.1000 174.1000 60.6000 174.2000 ;
	    RECT 63.4000 174.1000 68.9000 174.2000 ;
	    RECT 55.1000 173.9000 68.9000 174.1000 ;
	    RECT 55.3000 173.8000 55.7000 173.9000 ;
	    RECT 49.4000 171.1000 49.8000 173.4000 ;
	    RECT 51.8000 173.3000 53.7000 173.6000 ;
	    RECT 51.8000 171.1000 52.2000 173.3000 ;
	    RECT 53.3000 173.2000 53.7000 173.3000 ;
	    RECT 58.2000 172.8000 58.5000 173.9000 ;
	    RECT 59.8000 173.8000 64.2000 173.9000 ;
	    RECT 57.3000 172.7000 57.7000 172.8000 ;
	    RECT 54.2000 172.1000 54.6000 172.5000 ;
	    RECT 56.3000 172.4000 57.7000 172.7000 ;
	    RECT 58.2000 172.4000 58.6000 172.8000 ;
	    RECT 56.3000 172.1000 56.6000 172.4000 ;
	    RECT 59.0000 172.1000 59.4000 172.5000 ;
	    RECT 53.9000 171.8000 54.6000 172.1000 ;
	    RECT 53.9000 171.1000 54.5000 171.8000 ;
	    RECT 56.2000 171.1000 56.6000 172.1000 ;
	    RECT 58.4000 171.8000 59.4000 172.1000 ;
	    RECT 58.4000 171.1000 58.8000 171.8000 ;
	    RECT 60.6000 171.1000 61.0000 173.5000 ;
	    RECT 63.0000 171.1000 63.4000 173.5000 ;
	    RECT 65.5000 172.8000 65.8000 173.9000 ;
	    RECT 66.2000 173.8000 66.6000 173.9000 ;
	    RECT 68.3000 173.8000 68.7000 173.9000 ;
	    RECT 71.8000 173.6000 72.2000 174.8000 ;
	    RECT 72.6000 174.4000 73.0000 174.8000 ;
	    RECT 73.4000 173.7000 73.7000 175.2000 ;
	    RECT 75.0000 174.4000 75.4000 175.2000 ;
	    RECT 75.8000 173.7000 76.1000 175.2000 ;
	    RECT 77.4000 174.4000 77.8000 175.2000 ;
	    RECT 78.2000 173.7000 78.5000 175.2000 ;
	    RECT 83.0000 175.1000 83.4000 175.2000 ;
	    RECT 80.9000 174.8000 83.4000 175.1000 ;
	    RECT 80.9000 174.7000 81.3000 174.8000 ;
	    RECT 81.7000 174.2000 82.1000 174.3000 ;
	    RECT 85.4000 174.2000 85.7000 175.8000 ;
	    RECT 88.6000 175.6000 89.0000 175.8000 ;
	    RECT 86.9000 175.3000 89.0000 175.6000 ;
	    RECT 86.9000 175.2000 87.3000 175.3000 ;
	    RECT 87.7000 174.9000 88.1000 175.0000 ;
	    RECT 86.2000 174.6000 88.1000 174.9000 ;
	    RECT 86.2000 174.5000 86.6000 174.6000 ;
	    RECT 80.2000 173.9000 85.7000 174.2000 ;
	    RECT 80.2000 173.8000 81.0000 173.9000 ;
	    RECT 70.3000 173.3000 72.2000 173.6000 ;
	    RECT 70.3000 173.2000 70.7000 173.3000 ;
	    RECT 64.6000 172.1000 65.0000 172.5000 ;
	    RECT 65.4000 172.4000 65.8000 172.8000 ;
	    RECT 66.3000 172.7000 66.7000 172.8000 ;
	    RECT 66.3000 172.4000 67.7000 172.7000 ;
	    RECT 67.4000 172.1000 67.7000 172.4000 ;
	    RECT 69.4000 172.1000 69.8000 172.5000 ;
	    RECT 64.6000 171.8000 65.6000 172.1000 ;
	    RECT 65.2000 171.1000 65.6000 171.8000 ;
	    RECT 67.4000 171.1000 67.8000 172.1000 ;
	    RECT 69.4000 171.8000 70.1000 172.1000 ;
	    RECT 69.5000 171.1000 70.1000 171.8000 ;
	    RECT 71.8000 171.1000 72.2000 173.3000 ;
	    RECT 72.6000 173.4000 73.7000 173.7000 ;
	    RECT 75.0000 173.4000 76.1000 173.7000 ;
	    RECT 77.4000 173.4000 78.5000 173.7000 ;
	    RECT 72.6000 171.1000 73.0000 173.4000 ;
	    RECT 75.0000 171.1000 75.4000 173.4000 ;
	    RECT 77.4000 171.1000 77.8000 173.4000 ;
	    RECT 79.8000 171.1000 80.2000 173.5000 ;
	    RECT 82.3000 173.2000 82.6000 173.9000 ;
	    RECT 85.1000 173.8000 85.5000 173.9000 ;
	    RECT 88.6000 173.6000 89.0000 175.3000 ;
	    RECT 87.1000 173.3000 89.0000 173.6000 ;
	    RECT 87.1000 173.2000 87.5000 173.3000 ;
	    RECT 81.4000 172.1000 81.8000 172.5000 ;
	    RECT 82.2000 172.4000 82.6000 173.2000 ;
	    RECT 88.6000 173.1000 89.0000 173.3000 ;
	    RECT 89.4000 173.1000 89.8000 173.2000 ;
	    RECT 88.6000 172.8000 89.8000 173.1000 ;
	    RECT 83.1000 172.7000 83.5000 172.8000 ;
	    RECT 83.1000 172.4000 84.5000 172.7000 ;
	    RECT 84.2000 172.1000 84.5000 172.4000 ;
	    RECT 86.2000 172.1000 86.6000 172.5000 ;
	    RECT 81.4000 171.8000 82.4000 172.1000 ;
	    RECT 82.0000 171.1000 82.4000 171.8000 ;
	    RECT 84.2000 171.1000 84.6000 172.1000 ;
	    RECT 86.2000 171.8000 86.9000 172.1000 ;
	    RECT 86.3000 171.1000 86.9000 171.8000 ;
	    RECT 88.6000 171.1000 89.0000 172.8000 ;
	    RECT 89.4000 172.4000 89.8000 172.8000 ;
	    RECT 90.2000 173.1000 90.6000 179.9000 ;
	    RECT 92.3000 176.3000 92.7000 179.9000 ;
	    RECT 91.8000 175.9000 92.7000 176.3000 ;
	    RECT 93.4000 176.2000 93.8000 179.9000 ;
	    RECT 95.8000 176.2000 96.2000 179.9000 ;
	    RECT 93.4000 175.9000 94.5000 176.2000 ;
	    RECT 95.8000 175.9000 96.9000 176.2000 ;
	    RECT 91.9000 175.1000 92.2000 175.9000 ;
	    RECT 94.2000 175.6000 94.5000 175.9000 ;
	    RECT 96.6000 175.6000 96.9000 175.9000 ;
	    RECT 98.2000 175.7000 98.6000 179.9000 ;
	    RECT 100.4000 178.2000 100.8000 179.9000 ;
	    RECT 99.8000 177.9000 100.8000 178.2000 ;
	    RECT 102.6000 177.9000 103.0000 179.9000 ;
	    RECT 104.7000 177.9000 105.3000 179.9000 ;
	    RECT 99.8000 177.5000 100.2000 177.9000 ;
	    RECT 102.6000 177.6000 102.9000 177.9000 ;
	    RECT 101.5000 177.3000 103.3000 177.6000 ;
	    RECT 104.6000 177.5000 105.0000 177.9000 ;
	    RECT 101.5000 177.2000 101.9000 177.3000 ;
	    RECT 102.9000 177.2000 103.3000 177.3000 ;
	    RECT 99.8000 176.5000 100.2000 176.6000 ;
	    RECT 102.1000 176.5000 102.5000 176.6000 ;
	    RECT 99.8000 176.2000 102.5000 176.5000 ;
	    RECT 102.8000 176.5000 103.9000 176.8000 ;
	    RECT 102.8000 175.9000 103.1000 176.5000 ;
	    RECT 103.5000 176.4000 103.9000 176.5000 ;
	    RECT 104.7000 176.6000 105.4000 177.0000 ;
	    RECT 104.7000 176.1000 105.0000 176.6000 ;
	    RECT 100.7000 175.7000 103.1000 175.9000 ;
	    RECT 98.2000 175.6000 103.1000 175.7000 ;
	    RECT 103.8000 175.8000 105.0000 176.1000 ;
	    RECT 91.0000 174.8000 92.2000 175.1000 ;
	    RECT 92.6000 174.8000 93.0000 175.6000 ;
	    RECT 94.2000 175.2000 94.8000 175.6000 ;
	    RECT 96.6000 175.2000 97.2000 175.6000 ;
	    RECT 98.2000 175.5000 101.1000 175.6000 ;
	    RECT 98.2000 175.4000 101.0000 175.5000 ;
	    RECT 91.0000 174.2000 91.3000 174.8000 ;
	    RECT 91.9000 174.2000 92.2000 174.8000 ;
	    RECT 93.4000 174.4000 93.8000 175.2000 ;
	    RECT 91.0000 173.8000 91.4000 174.2000 ;
	    RECT 91.8000 173.8000 92.2000 174.2000 ;
	    RECT 91.0000 173.1000 91.4000 173.2000 ;
	    RECT 90.2000 172.8000 91.4000 173.1000 ;
	    RECT 90.2000 171.1000 90.6000 172.8000 ;
	    RECT 91.0000 172.4000 91.4000 172.8000 ;
	    RECT 91.9000 172.1000 92.2000 173.8000 ;
	    RECT 94.2000 173.7000 94.5000 175.2000 ;
	    RECT 95.8000 174.4000 96.2000 175.2000 ;
	    RECT 96.6000 173.7000 96.9000 175.2000 ;
	    RECT 101.4000 175.1000 101.8000 175.2000 ;
	    RECT 99.3000 174.8000 101.8000 175.1000 ;
	    RECT 99.3000 174.7000 99.7000 174.8000 ;
	    RECT 100.1000 174.2000 100.5000 174.3000 ;
	    RECT 103.8000 174.2000 104.1000 175.8000 ;
	    RECT 107.0000 175.6000 107.4000 179.9000 ;
	    RECT 107.8000 176.2000 108.2000 179.9000 ;
	    RECT 111.8000 176.2000 112.2000 179.9000 ;
	    RECT 107.8000 175.9000 108.9000 176.2000 ;
	    RECT 111.8000 175.9000 112.9000 176.2000 ;
	    RECT 105.3000 175.3000 107.4000 175.6000 ;
	    RECT 105.3000 175.2000 105.7000 175.3000 ;
	    RECT 106.1000 174.9000 106.5000 175.0000 ;
	    RECT 104.6000 174.6000 106.5000 174.9000 ;
	    RECT 104.6000 174.5000 105.0000 174.6000 ;
	    RECT 98.6000 173.9000 104.2000 174.2000 ;
	    RECT 98.6000 173.8000 99.4000 173.9000 ;
	    RECT 91.8000 171.1000 92.2000 172.1000 ;
	    RECT 93.4000 173.4000 94.5000 173.7000 ;
	    RECT 95.8000 173.4000 96.9000 173.7000 ;
	    RECT 93.4000 171.1000 93.8000 173.4000 ;
	    RECT 95.8000 171.1000 96.2000 173.4000 ;
	    RECT 98.2000 171.1000 98.6000 173.5000 ;
	    RECT 100.7000 172.8000 101.0000 173.9000 ;
	    RECT 103.5000 173.8000 104.2000 173.9000 ;
	    RECT 107.0000 173.6000 107.4000 175.3000 ;
	    RECT 108.6000 175.6000 108.9000 175.9000 ;
	    RECT 112.6000 175.6000 112.9000 175.9000 ;
	    RECT 114.2000 175.6000 114.6000 179.9000 ;
	    RECT 116.3000 177.9000 116.9000 179.9000 ;
	    RECT 118.6000 177.9000 119.0000 179.9000 ;
	    RECT 120.8000 178.2000 121.2000 179.9000 ;
	    RECT 120.8000 177.9000 121.8000 178.2000 ;
	    RECT 116.6000 177.5000 117.0000 177.9000 ;
	    RECT 118.7000 177.6000 119.0000 177.9000 ;
	    RECT 118.3000 177.3000 120.1000 177.6000 ;
	    RECT 121.4000 177.5000 121.8000 177.9000 ;
	    RECT 118.3000 177.2000 118.7000 177.3000 ;
	    RECT 119.7000 177.2000 120.1000 177.3000 ;
	    RECT 116.2000 176.6000 116.9000 177.0000 ;
	    RECT 116.6000 176.1000 116.9000 176.6000 ;
	    RECT 117.7000 176.5000 118.8000 176.8000 ;
	    RECT 117.7000 176.4000 118.1000 176.5000 ;
	    RECT 116.6000 175.8000 117.8000 176.1000 ;
	    RECT 108.6000 175.2000 109.2000 175.6000 ;
	    RECT 112.6000 175.2000 113.2000 175.6000 ;
	    RECT 114.2000 175.3000 116.3000 175.6000 ;
	    RECT 107.8000 174.4000 108.2000 175.2000 ;
	    RECT 108.6000 173.7000 108.9000 175.2000 ;
	    RECT 111.8000 174.4000 112.2000 175.2000 ;
	    RECT 112.6000 173.7000 112.9000 175.2000 ;
	    RECT 105.5000 173.3000 107.4000 173.6000 ;
	    RECT 105.5000 173.2000 105.9000 173.3000 ;
	    RECT 99.8000 172.1000 100.2000 172.5000 ;
	    RECT 100.6000 172.4000 101.0000 172.8000 ;
	    RECT 101.5000 172.7000 101.9000 172.8000 ;
	    RECT 101.5000 172.4000 102.9000 172.7000 ;
	    RECT 102.6000 172.1000 102.9000 172.4000 ;
	    RECT 104.6000 172.1000 105.0000 172.5000 ;
	    RECT 99.8000 171.8000 100.8000 172.1000 ;
	    RECT 100.4000 171.1000 100.8000 171.8000 ;
	    RECT 102.6000 171.1000 103.0000 172.1000 ;
	    RECT 104.6000 171.8000 105.3000 172.1000 ;
	    RECT 104.7000 171.1000 105.3000 171.8000 ;
	    RECT 107.0000 171.1000 107.4000 173.3000 ;
	    RECT 107.8000 173.4000 108.9000 173.7000 ;
	    RECT 111.8000 173.4000 112.9000 173.7000 ;
	    RECT 114.2000 173.6000 114.6000 175.3000 ;
	    RECT 115.9000 175.2000 116.3000 175.3000 ;
	    RECT 115.1000 174.9000 115.5000 175.0000 ;
	    RECT 115.1000 174.6000 117.0000 174.9000 ;
	    RECT 116.6000 174.5000 117.0000 174.6000 ;
	    RECT 117.5000 174.2000 117.8000 175.8000 ;
	    RECT 118.5000 175.9000 118.8000 176.5000 ;
	    RECT 119.1000 176.5000 119.5000 176.6000 ;
	    RECT 121.4000 176.5000 121.8000 176.6000 ;
	    RECT 119.1000 176.2000 121.8000 176.5000 ;
	    RECT 118.5000 175.7000 120.9000 175.9000 ;
	    RECT 123.0000 175.7000 123.4000 179.9000 ;
	    RECT 125.4000 176.2000 125.8000 179.9000 ;
	    RECT 118.5000 175.6000 123.4000 175.7000 ;
	    RECT 124.7000 175.9000 125.8000 176.2000 ;
	    RECT 126.5000 176.3000 126.9000 179.9000 ;
	    RECT 126.5000 175.9000 127.4000 176.3000 ;
	    RECT 124.7000 175.6000 125.0000 175.9000 ;
	    RECT 120.5000 175.5000 123.4000 175.6000 ;
	    RECT 120.6000 175.4000 123.4000 175.5000 ;
	    RECT 124.4000 175.2000 125.0000 175.6000 ;
	    RECT 119.8000 175.1000 120.2000 175.2000 ;
	    RECT 119.8000 174.8000 122.3000 175.1000 ;
	    RECT 120.6000 174.7000 121.0000 174.8000 ;
	    RECT 121.9000 174.7000 122.3000 174.8000 ;
	    RECT 121.1000 174.2000 121.5000 174.3000 ;
	    RECT 117.5000 173.9000 123.0000 174.2000 ;
	    RECT 117.7000 173.8000 118.1000 173.9000 ;
	    RECT 107.8000 171.1000 108.2000 173.4000 ;
	    RECT 111.8000 171.1000 112.2000 173.4000 ;
	    RECT 114.2000 173.3000 116.1000 173.6000 ;
	    RECT 114.2000 171.1000 114.6000 173.3000 ;
	    RECT 115.7000 173.2000 116.1000 173.3000 ;
	    RECT 120.6000 173.2000 120.9000 173.9000 ;
	    RECT 122.2000 173.8000 123.0000 173.9000 ;
	    RECT 124.7000 173.7000 125.0000 175.2000 ;
	    RECT 125.4000 174.4000 125.8000 175.2000 ;
	    RECT 126.2000 174.8000 126.6000 175.6000 ;
	    RECT 127.0000 174.2000 127.3000 175.9000 ;
	    RECT 127.0000 174.1000 127.4000 174.2000 ;
	    RECT 127.8000 174.1000 128.2000 174.2000 ;
	    RECT 127.0000 173.8000 128.2000 174.1000 ;
	    RECT 119.7000 172.7000 120.1000 172.8000 ;
	    RECT 116.6000 172.1000 117.0000 172.5000 ;
	    RECT 118.7000 172.4000 120.1000 172.7000 ;
	    RECT 120.6000 172.4000 121.0000 173.2000 ;
	    RECT 118.7000 172.1000 119.0000 172.4000 ;
	    RECT 121.4000 172.1000 121.8000 172.5000 ;
	    RECT 116.3000 171.8000 117.0000 172.1000 ;
	    RECT 116.3000 171.1000 116.9000 171.8000 ;
	    RECT 118.6000 171.1000 119.0000 172.1000 ;
	    RECT 120.8000 171.8000 121.8000 172.1000 ;
	    RECT 120.8000 171.1000 121.2000 171.8000 ;
	    RECT 123.0000 171.1000 123.4000 173.5000 ;
	    RECT 124.7000 173.4000 125.8000 173.7000 ;
	    RECT 125.4000 171.1000 125.8000 173.4000 ;
	    RECT 127.0000 172.1000 127.3000 173.8000 ;
	    RECT 127.8000 173.1000 128.2000 173.2000 ;
	    RECT 128.6000 173.1000 129.0000 179.9000 ;
	    RECT 130.2000 176.2000 130.6000 179.9000 ;
	    RECT 130.2000 175.9000 131.3000 176.2000 ;
	    RECT 131.0000 175.6000 131.3000 175.9000 ;
	    RECT 132.6000 175.7000 133.0000 179.9000 ;
	    RECT 134.8000 178.2000 135.2000 179.9000 ;
	    RECT 134.2000 177.9000 135.2000 178.2000 ;
	    RECT 137.0000 177.9000 137.4000 179.9000 ;
	    RECT 139.1000 177.9000 139.7000 179.9000 ;
	    RECT 134.2000 177.5000 134.6000 177.9000 ;
	    RECT 137.0000 177.6000 137.3000 177.9000 ;
	    RECT 135.9000 177.3000 137.7000 177.6000 ;
	    RECT 139.0000 177.5000 139.4000 177.9000 ;
	    RECT 135.9000 177.2000 136.3000 177.3000 ;
	    RECT 137.3000 177.2000 137.7000 177.3000 ;
	    RECT 134.2000 176.5000 134.6000 176.6000 ;
	    RECT 136.5000 176.5000 136.9000 176.6000 ;
	    RECT 134.2000 176.2000 136.9000 176.5000 ;
	    RECT 137.2000 176.5000 138.3000 176.8000 ;
	    RECT 137.2000 175.9000 137.5000 176.5000 ;
	    RECT 137.9000 176.4000 138.3000 176.5000 ;
	    RECT 139.1000 176.6000 139.8000 177.0000 ;
	    RECT 139.1000 176.1000 139.4000 176.6000 ;
	    RECT 135.1000 175.7000 137.5000 175.9000 ;
	    RECT 132.6000 175.6000 137.5000 175.7000 ;
	    RECT 138.2000 175.8000 139.4000 176.1000 ;
	    RECT 131.0000 175.2000 131.6000 175.6000 ;
	    RECT 132.6000 175.5000 135.5000 175.6000 ;
	    RECT 132.6000 175.4000 135.4000 175.5000 ;
	    RECT 129.4000 175.1000 129.8000 175.2000 ;
	    RECT 130.2000 175.1000 130.6000 175.2000 ;
	    RECT 129.4000 174.8000 130.6000 175.1000 ;
	    RECT 130.2000 174.4000 130.6000 174.8000 ;
	    RECT 131.0000 173.7000 131.3000 175.2000 ;
	    RECT 135.8000 175.1000 136.2000 175.2000 ;
	    RECT 133.7000 174.8000 136.2000 175.1000 ;
	    RECT 133.7000 174.7000 134.1000 174.8000 ;
	    RECT 134.5000 174.2000 134.9000 174.3000 ;
	    RECT 138.2000 174.2000 138.5000 175.8000 ;
	    RECT 141.4000 175.6000 141.8000 179.9000 ;
	    RECT 142.2000 176.2000 142.6000 179.9000 ;
	    RECT 144.6000 176.2000 145.0000 179.9000 ;
	    RECT 147.0000 176.2000 147.4000 179.9000 ;
	    RECT 149.4000 176.2000 149.8000 179.9000 ;
	    RECT 153.4000 176.2000 153.8000 179.9000 ;
	    RECT 142.2000 175.9000 143.3000 176.2000 ;
	    RECT 144.6000 175.9000 145.7000 176.2000 ;
	    RECT 147.0000 175.9000 148.1000 176.2000 ;
	    RECT 149.4000 175.9000 150.5000 176.2000 ;
	    RECT 139.7000 175.3000 141.8000 175.6000 ;
	    RECT 139.7000 175.2000 140.1000 175.3000 ;
	    RECT 140.5000 174.9000 140.9000 175.0000 ;
	    RECT 139.0000 174.6000 140.9000 174.9000 ;
	    RECT 139.0000 174.5000 139.4000 174.6000 ;
	    RECT 133.0000 173.9000 138.5000 174.2000 ;
	    RECT 133.0000 173.8000 133.8000 173.9000 ;
	    RECT 130.2000 173.4000 131.3000 173.7000 ;
	    RECT 127.8000 172.8000 129.0000 173.1000 ;
	    RECT 127.8000 172.4000 128.2000 172.8000 ;
	    RECT 127.0000 171.1000 127.4000 172.1000 ;
	    RECT 128.6000 171.1000 129.0000 172.8000 ;
	    RECT 129.4000 172.4000 129.8000 173.2000 ;
	    RECT 130.2000 171.1000 130.6000 173.4000 ;
	    RECT 132.6000 171.1000 133.0000 173.5000 ;
	    RECT 135.1000 172.8000 135.4000 173.9000 ;
	    RECT 137.9000 173.8000 138.3000 173.9000 ;
	    RECT 141.4000 173.6000 141.8000 175.3000 ;
	    RECT 143.0000 175.6000 143.3000 175.9000 ;
	    RECT 145.4000 175.6000 145.7000 175.9000 ;
	    RECT 147.8000 175.6000 148.1000 175.9000 ;
	    RECT 150.2000 175.6000 150.5000 175.9000 ;
	    RECT 152.7000 175.9000 153.8000 176.2000 ;
	    RECT 152.7000 175.6000 153.0000 175.9000 ;
	    RECT 143.0000 175.2000 143.6000 175.6000 ;
	    RECT 145.4000 175.2000 146.0000 175.6000 ;
	    RECT 147.8000 175.2000 148.4000 175.6000 ;
	    RECT 150.2000 175.2000 150.8000 175.6000 ;
	    RECT 152.4000 175.2000 153.0000 175.6000 ;
	    RECT 154.2000 175.6000 154.6000 179.9000 ;
	    RECT 156.3000 177.9000 156.9000 179.9000 ;
	    RECT 158.6000 177.9000 159.0000 179.9000 ;
	    RECT 160.8000 178.2000 161.2000 179.9000 ;
	    RECT 160.8000 177.9000 161.8000 178.2000 ;
	    RECT 156.6000 177.5000 157.0000 177.9000 ;
	    RECT 158.7000 177.6000 159.0000 177.9000 ;
	    RECT 158.3000 177.3000 160.1000 177.6000 ;
	    RECT 161.4000 177.5000 161.8000 177.9000 ;
	    RECT 158.3000 177.2000 158.7000 177.3000 ;
	    RECT 159.7000 177.2000 160.1000 177.3000 ;
	    RECT 156.2000 176.6000 156.9000 177.0000 ;
	    RECT 156.6000 176.1000 156.9000 176.6000 ;
	    RECT 157.7000 176.5000 158.8000 176.8000 ;
	    RECT 157.7000 176.4000 158.1000 176.5000 ;
	    RECT 156.6000 175.8000 157.8000 176.1000 ;
	    RECT 154.2000 175.3000 156.3000 175.6000 ;
	    RECT 142.2000 174.4000 142.6000 175.2000 ;
	    RECT 143.0000 173.7000 143.3000 175.2000 ;
	    RECT 144.6000 174.4000 145.0000 175.2000 ;
	    RECT 145.4000 173.7000 145.7000 175.2000 ;
	    RECT 147.0000 174.4000 147.4000 175.2000 ;
	    RECT 147.8000 173.7000 148.1000 175.2000 ;
	    RECT 149.4000 174.4000 149.8000 175.2000 ;
	    RECT 150.2000 173.7000 150.5000 175.2000 ;
	    RECT 139.9000 173.3000 141.8000 173.6000 ;
	    RECT 139.9000 173.2000 140.3000 173.3000 ;
	    RECT 134.2000 172.1000 134.6000 172.5000 ;
	    RECT 135.0000 172.4000 135.4000 172.8000 ;
	    RECT 135.9000 172.7000 136.3000 172.8000 ;
	    RECT 135.9000 172.4000 137.3000 172.7000 ;
	    RECT 137.0000 172.1000 137.3000 172.4000 ;
	    RECT 139.0000 172.1000 139.4000 172.5000 ;
	    RECT 134.2000 171.8000 135.2000 172.1000 ;
	    RECT 134.8000 171.1000 135.2000 171.8000 ;
	    RECT 137.0000 171.1000 137.4000 172.1000 ;
	    RECT 139.0000 171.8000 139.7000 172.1000 ;
	    RECT 139.1000 171.1000 139.7000 171.8000 ;
	    RECT 141.4000 171.1000 141.8000 173.3000 ;
	    RECT 142.2000 173.4000 143.3000 173.7000 ;
	    RECT 144.6000 173.4000 145.7000 173.7000 ;
	    RECT 147.0000 173.4000 148.1000 173.7000 ;
	    RECT 149.4000 173.4000 150.5000 173.7000 ;
	    RECT 152.7000 173.7000 153.0000 175.2000 ;
	    RECT 153.4000 174.4000 153.8000 175.2000 ;
	    RECT 152.7000 173.4000 153.8000 173.7000 ;
	    RECT 142.2000 171.1000 142.6000 173.4000 ;
	    RECT 144.6000 171.1000 145.0000 173.4000 ;
	    RECT 147.0000 171.1000 147.4000 173.4000 ;
	    RECT 149.4000 171.1000 149.8000 173.4000 ;
	    RECT 153.4000 171.1000 153.8000 173.4000 ;
	    RECT 154.2000 173.6000 154.6000 175.3000 ;
	    RECT 155.9000 175.2000 156.3000 175.3000 ;
	    RECT 155.1000 174.9000 155.5000 175.0000 ;
	    RECT 155.1000 174.6000 157.0000 174.9000 ;
	    RECT 156.6000 174.5000 157.0000 174.6000 ;
	    RECT 157.5000 174.2000 157.8000 175.8000 ;
	    RECT 158.5000 175.9000 158.8000 176.5000 ;
	    RECT 159.1000 176.5000 159.5000 176.6000 ;
	    RECT 161.4000 176.5000 161.8000 176.6000 ;
	    RECT 159.1000 176.2000 161.8000 176.5000 ;
	    RECT 158.5000 175.7000 160.9000 175.9000 ;
	    RECT 163.0000 175.7000 163.4000 179.9000 ;
	    RECT 158.5000 175.6000 163.4000 175.7000 ;
	    RECT 160.5000 175.5000 163.4000 175.6000 ;
	    RECT 160.6000 175.4000 163.4000 175.5000 ;
	    RECT 159.8000 175.1000 160.2000 175.2000 ;
	    RECT 159.8000 174.8000 162.3000 175.1000 ;
	    RECT 160.6000 174.7000 161.0000 174.8000 ;
	    RECT 161.9000 174.7000 162.3000 174.8000 ;
	    RECT 161.1000 174.2000 161.5000 174.3000 ;
	    RECT 157.5000 174.1000 163.0000 174.2000 ;
	    RECT 164.6000 174.1000 165.0000 174.2000 ;
	    RECT 157.5000 173.9000 165.0000 174.1000 ;
	    RECT 157.7000 173.8000 158.1000 173.9000 ;
	    RECT 154.2000 173.3000 156.1000 173.6000 ;
	    RECT 154.2000 171.1000 154.6000 173.3000 ;
	    RECT 155.7000 173.2000 156.1000 173.3000 ;
	    RECT 160.6000 172.8000 160.9000 173.9000 ;
	    RECT 162.2000 173.8000 165.0000 173.9000 ;
	    RECT 159.7000 172.7000 160.1000 172.8000 ;
	    RECT 156.6000 172.1000 157.0000 172.5000 ;
	    RECT 158.7000 172.4000 160.1000 172.7000 ;
	    RECT 160.6000 172.4000 161.0000 172.8000 ;
	    RECT 158.7000 172.1000 159.0000 172.4000 ;
	    RECT 161.4000 172.1000 161.8000 172.5000 ;
	    RECT 156.3000 171.8000 157.0000 172.1000 ;
	    RECT 156.3000 171.1000 156.9000 171.8000 ;
	    RECT 158.6000 171.1000 159.0000 172.1000 ;
	    RECT 160.8000 171.8000 161.8000 172.1000 ;
	    RECT 160.8000 171.1000 161.2000 171.8000 ;
	    RECT 163.0000 171.1000 163.4000 173.5000 ;
	    RECT 165.4000 172.4000 165.8000 173.2000 ;
	    RECT 166.2000 171.1000 166.6000 179.9000 ;
	    RECT 167.0000 176.2000 167.4000 179.9000 ;
	    RECT 171.0000 176.2000 171.4000 179.9000 ;
	    RECT 167.0000 175.9000 168.1000 176.2000 ;
	    RECT 167.8000 175.6000 168.1000 175.9000 ;
	    RECT 170.3000 175.9000 171.4000 176.2000 ;
	    RECT 171.8000 176.2000 172.2000 179.9000 ;
	    RECT 171.8000 175.9000 172.9000 176.2000 ;
	    RECT 170.3000 175.6000 170.6000 175.9000 ;
	    RECT 167.8000 175.2000 168.4000 175.6000 ;
	    RECT 170.0000 175.2000 170.6000 175.6000 ;
	    RECT 172.6000 175.6000 172.9000 175.9000 ;
	    RECT 174.2000 175.7000 174.6000 179.9000 ;
	    RECT 176.4000 178.2000 176.8000 179.9000 ;
	    RECT 175.8000 177.9000 176.8000 178.2000 ;
	    RECT 178.6000 177.9000 179.0000 179.9000 ;
	    RECT 180.7000 177.9000 181.3000 179.9000 ;
	    RECT 175.8000 177.5000 176.2000 177.9000 ;
	    RECT 178.6000 177.6000 178.9000 177.9000 ;
	    RECT 177.5000 177.3000 179.3000 177.6000 ;
	    RECT 180.6000 177.5000 181.0000 177.9000 ;
	    RECT 177.5000 177.2000 177.9000 177.3000 ;
	    RECT 178.9000 177.2000 179.3000 177.3000 ;
	    RECT 175.8000 176.5000 176.2000 176.6000 ;
	    RECT 178.1000 176.5000 178.5000 176.6000 ;
	    RECT 175.8000 176.2000 178.5000 176.5000 ;
	    RECT 178.8000 176.5000 179.9000 176.8000 ;
	    RECT 178.8000 175.9000 179.1000 176.5000 ;
	    RECT 179.5000 176.4000 179.9000 176.5000 ;
	    RECT 180.7000 176.6000 181.4000 177.0000 ;
	    RECT 180.7000 176.1000 181.0000 176.6000 ;
	    RECT 176.7000 175.7000 179.1000 175.9000 ;
	    RECT 174.2000 175.6000 179.1000 175.7000 ;
	    RECT 179.8000 175.8000 181.0000 176.1000 ;
	    RECT 172.6000 175.2000 173.2000 175.6000 ;
	    RECT 174.2000 175.5000 177.1000 175.6000 ;
	    RECT 174.2000 175.4000 177.0000 175.5000 ;
	    RECT 167.0000 174.4000 167.4000 175.2000 ;
	    RECT 167.8000 173.7000 168.1000 175.2000 ;
	    RECT 167.0000 173.4000 168.1000 173.7000 ;
	    RECT 170.3000 173.7000 170.6000 175.2000 ;
	    RECT 171.0000 174.4000 171.4000 175.2000 ;
	    RECT 171.8000 174.4000 172.2000 175.2000 ;
	    RECT 172.6000 173.7000 172.9000 175.2000 ;
	    RECT 177.4000 175.1000 177.8000 175.2000 ;
	    RECT 175.3000 174.8000 177.8000 175.1000 ;
	    RECT 175.3000 174.7000 175.7000 174.8000 ;
	    RECT 176.1000 174.2000 176.5000 174.3000 ;
	    RECT 179.8000 174.2000 180.1000 175.8000 ;
	    RECT 183.0000 175.6000 183.4000 179.9000 ;
	    RECT 184.1000 176.3000 184.5000 179.9000 ;
	    RECT 184.1000 175.9000 185.0000 176.3000 ;
	    RECT 181.3000 175.3000 183.4000 175.6000 ;
	    RECT 181.3000 175.2000 181.7000 175.3000 ;
	    RECT 182.1000 174.9000 182.5000 175.0000 ;
	    RECT 180.6000 174.6000 182.5000 174.9000 ;
	    RECT 180.6000 174.5000 181.0000 174.6000 ;
	    RECT 174.6000 173.9000 180.1000 174.2000 ;
	    RECT 174.6000 173.8000 175.4000 173.9000 ;
	    RECT 170.3000 173.4000 171.4000 173.7000 ;
	    RECT 167.0000 171.1000 167.4000 173.4000 ;
	    RECT 171.0000 171.1000 171.4000 173.4000 ;
	    RECT 171.8000 173.4000 172.9000 173.7000 ;
	    RECT 171.8000 171.1000 172.2000 173.4000 ;
	    RECT 174.2000 171.1000 174.6000 173.5000 ;
	    RECT 176.7000 172.8000 177.0000 173.9000 ;
	    RECT 179.5000 173.8000 179.9000 173.9000 ;
	    RECT 183.0000 173.6000 183.4000 175.3000 ;
	    RECT 183.8000 174.8000 184.2000 175.6000 ;
	    RECT 184.6000 174.2000 184.9000 175.9000 ;
	    RECT 181.5000 173.3000 183.4000 173.6000 ;
	    RECT 181.5000 173.2000 181.9000 173.3000 ;
	    RECT 175.8000 172.1000 176.2000 172.5000 ;
	    RECT 176.6000 172.4000 177.0000 172.8000 ;
	    RECT 177.5000 172.7000 177.9000 172.8000 ;
	    RECT 177.5000 172.4000 178.9000 172.7000 ;
	    RECT 178.6000 172.1000 178.9000 172.4000 ;
	    RECT 180.6000 172.1000 181.0000 172.5000 ;
	    RECT 175.8000 171.8000 176.8000 172.1000 ;
	    RECT 176.4000 171.1000 176.8000 171.8000 ;
	    RECT 178.6000 171.1000 179.0000 172.1000 ;
	    RECT 180.6000 171.8000 181.3000 172.1000 ;
	    RECT 180.7000 171.1000 181.3000 171.8000 ;
	    RECT 183.0000 171.1000 183.4000 173.3000 ;
	    RECT 183.8000 173.8000 184.2000 174.2000 ;
	    RECT 184.6000 173.8000 185.0000 174.2000 ;
	    RECT 183.8000 173.1000 184.1000 173.8000 ;
	    RECT 184.6000 173.1000 184.9000 173.8000 ;
	    RECT 183.8000 172.8000 184.9000 173.1000 ;
	    RECT 184.6000 172.1000 184.9000 172.8000 ;
	    RECT 185.4000 173.1000 185.8000 173.2000 ;
	    RECT 186.2000 173.1000 186.6000 179.9000 ;
	    RECT 187.8000 176.2000 188.2000 179.9000 ;
	    RECT 187.8000 175.9000 188.9000 176.2000 ;
	    RECT 188.6000 175.6000 188.9000 175.9000 ;
	    RECT 190.2000 175.7000 190.6000 179.9000 ;
	    RECT 192.4000 178.2000 192.8000 179.9000 ;
	    RECT 191.8000 177.9000 192.8000 178.2000 ;
	    RECT 194.6000 177.9000 195.0000 179.9000 ;
	    RECT 196.7000 177.9000 197.3000 179.9000 ;
	    RECT 191.8000 177.5000 192.2000 177.9000 ;
	    RECT 194.6000 177.6000 194.9000 177.9000 ;
	    RECT 193.5000 177.3000 195.3000 177.6000 ;
	    RECT 196.6000 177.5000 197.0000 177.9000 ;
	    RECT 193.5000 177.2000 193.9000 177.3000 ;
	    RECT 194.9000 177.2000 195.3000 177.3000 ;
	    RECT 191.8000 176.5000 192.2000 176.6000 ;
	    RECT 194.1000 176.5000 194.5000 176.6000 ;
	    RECT 191.8000 176.2000 194.5000 176.5000 ;
	    RECT 194.8000 176.5000 195.9000 176.8000 ;
	    RECT 194.8000 175.9000 195.1000 176.5000 ;
	    RECT 195.5000 176.4000 195.9000 176.5000 ;
	    RECT 196.7000 176.6000 197.4000 177.0000 ;
	    RECT 196.7000 176.1000 197.0000 176.6000 ;
	    RECT 192.7000 175.7000 195.1000 175.9000 ;
	    RECT 190.2000 175.6000 195.1000 175.7000 ;
	    RECT 195.8000 175.8000 197.0000 176.1000 ;
	    RECT 188.6000 175.2000 189.2000 175.6000 ;
	    RECT 190.2000 175.5000 193.1000 175.6000 ;
	    RECT 190.2000 175.4000 193.0000 175.5000 ;
	    RECT 187.0000 175.1000 187.4000 175.2000 ;
	    RECT 187.8000 175.1000 188.2000 175.2000 ;
	    RECT 187.0000 174.8000 188.2000 175.1000 ;
	    RECT 187.8000 174.4000 188.2000 174.8000 ;
	    RECT 188.6000 173.7000 188.9000 175.2000 ;
	    RECT 193.4000 175.1000 193.8000 175.2000 ;
	    RECT 191.3000 174.8000 193.8000 175.1000 ;
	    RECT 191.3000 174.7000 191.7000 174.8000 ;
	    RECT 192.1000 174.2000 192.5000 174.3000 ;
	    RECT 195.8000 174.2000 196.1000 175.8000 ;
	    RECT 199.0000 175.6000 199.4000 179.9000 ;
	    RECT 201.1000 176.2000 201.5000 179.9000 ;
	    RECT 201.8000 176.8000 202.2000 177.2000 ;
	    RECT 201.9000 176.2000 202.2000 176.8000 ;
	    RECT 203.0000 176.2000 203.4000 179.9000 ;
	    RECT 204.6000 176.2000 205.0000 179.9000 ;
	    RECT 201.1000 175.9000 201.6000 176.2000 ;
	    RECT 201.9000 175.9000 202.6000 176.2000 ;
	    RECT 203.0000 175.9000 205.0000 176.2000 ;
	    RECT 197.3000 175.3000 199.4000 175.6000 ;
	    RECT 197.3000 175.2000 197.7000 175.3000 ;
	    RECT 198.1000 174.9000 198.5000 175.0000 ;
	    RECT 196.6000 174.6000 198.5000 174.9000 ;
	    RECT 196.6000 174.5000 197.0000 174.6000 ;
	    RECT 190.6000 173.9000 196.1000 174.2000 ;
	    RECT 190.6000 173.8000 191.4000 173.9000 ;
	    RECT 187.8000 173.4000 188.9000 173.7000 ;
	    RECT 185.4000 172.8000 186.6000 173.1000 ;
	    RECT 185.4000 172.4000 185.8000 172.8000 ;
	    RECT 184.6000 171.1000 185.0000 172.1000 ;
	    RECT 186.2000 171.1000 186.6000 172.8000 ;
	    RECT 187.0000 172.4000 187.4000 173.2000 ;
	    RECT 187.8000 171.1000 188.2000 173.4000 ;
	    RECT 190.2000 171.1000 190.6000 173.5000 ;
	    RECT 192.7000 172.8000 193.0000 173.9000 ;
	    RECT 195.5000 173.8000 195.9000 173.9000 ;
	    RECT 199.0000 173.6000 199.4000 175.3000 ;
	    RECT 200.6000 174.4000 201.0000 175.2000 ;
	    RECT 201.3000 175.1000 201.6000 175.9000 ;
	    RECT 202.2000 175.8000 202.6000 175.9000 ;
	    RECT 205.4000 175.8000 205.8000 179.9000 ;
	    RECT 203.4000 175.2000 203.8000 175.4000 ;
	    RECT 205.4000 175.2000 205.7000 175.8000 ;
	    RECT 206.2000 175.7000 206.6000 179.9000 ;
	    RECT 208.4000 178.2000 208.8000 179.9000 ;
	    RECT 207.8000 177.9000 208.8000 178.2000 ;
	    RECT 210.6000 177.9000 211.0000 179.9000 ;
	    RECT 212.7000 177.9000 213.3000 179.9000 ;
	    RECT 207.8000 177.5000 208.2000 177.9000 ;
	    RECT 210.6000 177.6000 210.9000 177.9000 ;
	    RECT 209.5000 177.3000 211.3000 177.6000 ;
	    RECT 212.6000 177.5000 213.0000 177.9000 ;
	    RECT 209.5000 177.2000 209.9000 177.3000 ;
	    RECT 210.9000 177.2000 211.3000 177.3000 ;
	    RECT 207.8000 176.5000 208.2000 176.6000 ;
	    RECT 210.1000 176.5000 210.5000 176.6000 ;
	    RECT 207.8000 176.2000 210.5000 176.5000 ;
	    RECT 210.8000 176.5000 211.9000 176.8000 ;
	    RECT 210.8000 175.9000 211.1000 176.5000 ;
	    RECT 211.5000 176.4000 211.9000 176.5000 ;
	    RECT 212.7000 176.6000 213.4000 177.0000 ;
	    RECT 212.7000 176.1000 213.0000 176.6000 ;
	    RECT 208.7000 175.7000 211.1000 175.9000 ;
	    RECT 206.2000 175.6000 211.1000 175.7000 ;
	    RECT 211.8000 175.8000 213.0000 176.1000 ;
	    RECT 206.2000 175.5000 209.1000 175.6000 ;
	    RECT 206.2000 175.4000 209.0000 175.5000 ;
	    RECT 203.0000 175.1000 203.8000 175.2000 ;
	    RECT 201.3000 174.9000 203.8000 175.1000 ;
	    RECT 204.6000 174.9000 205.8000 175.2000 ;
	    RECT 209.4000 175.1000 209.8000 175.2000 ;
	    RECT 201.3000 174.8000 203.4000 174.9000 ;
	    RECT 201.3000 174.2000 201.6000 174.8000 ;
	    RECT 199.8000 174.1000 200.2000 174.2000 ;
	    RECT 199.8000 173.8000 200.6000 174.1000 ;
	    RECT 201.3000 173.8000 202.6000 174.2000 ;
	    RECT 203.8000 173.8000 204.2000 174.6000 ;
	    RECT 200.2000 173.6000 200.6000 173.8000 ;
	    RECT 197.5000 173.3000 199.4000 173.6000 ;
	    RECT 197.5000 173.2000 197.9000 173.3000 ;
	    RECT 191.8000 172.1000 192.2000 172.5000 ;
	    RECT 192.6000 172.4000 193.0000 172.8000 ;
	    RECT 193.5000 172.7000 193.9000 172.8000 ;
	    RECT 193.5000 172.4000 194.9000 172.7000 ;
	    RECT 194.6000 172.1000 194.9000 172.4000 ;
	    RECT 196.6000 172.1000 197.0000 172.5000 ;
	    RECT 191.8000 171.8000 192.8000 172.1000 ;
	    RECT 192.4000 171.1000 192.8000 171.8000 ;
	    RECT 194.6000 171.1000 195.0000 172.1000 ;
	    RECT 196.6000 171.8000 197.3000 172.1000 ;
	    RECT 196.7000 171.1000 197.3000 171.8000 ;
	    RECT 199.0000 171.1000 199.4000 173.3000 ;
	    RECT 199.9000 173.1000 201.7000 173.3000 ;
	    RECT 202.2000 173.1000 202.5000 173.8000 ;
	    RECT 204.6000 173.1000 204.9000 174.9000 ;
	    RECT 205.4000 174.8000 205.8000 174.9000 ;
	    RECT 207.3000 174.8000 209.8000 175.1000 ;
	    RECT 207.3000 174.7000 207.7000 174.8000 ;
	    RECT 208.6000 174.7000 209.0000 174.8000 ;
	    RECT 208.1000 174.2000 208.5000 174.3000 ;
	    RECT 211.8000 174.2000 212.1000 175.8000 ;
	    RECT 215.0000 175.6000 215.4000 179.9000 ;
	    RECT 217.7000 176.3000 218.1000 179.9000 ;
	    RECT 217.7000 175.9000 218.6000 176.3000 ;
	    RECT 221.1000 176.2000 221.5000 179.9000 ;
	    RECT 221.8000 176.8000 222.2000 177.2000 ;
	    RECT 221.9000 176.2000 222.2000 176.8000 ;
	    RECT 221.1000 175.9000 221.6000 176.2000 ;
	    RECT 221.9000 175.9000 222.6000 176.2000 ;
	    RECT 213.3000 175.3000 215.4000 175.6000 ;
	    RECT 213.3000 175.2000 213.7000 175.3000 ;
	    RECT 214.1000 174.9000 214.5000 175.0000 ;
	    RECT 212.6000 174.6000 214.5000 174.9000 ;
	    RECT 212.6000 174.5000 213.0000 174.6000 ;
	    RECT 206.6000 173.9000 212.1000 174.2000 ;
	    RECT 206.6000 173.8000 207.4000 173.9000 ;
	    RECT 199.8000 173.0000 201.8000 173.1000 ;
	    RECT 199.8000 171.1000 200.2000 173.0000 ;
	    RECT 201.4000 171.1000 201.8000 173.0000 ;
	    RECT 202.2000 171.1000 202.6000 173.1000 ;
	    RECT 204.6000 171.1000 205.0000 173.1000 ;
	    RECT 205.4000 172.8000 205.8000 173.2000 ;
	    RECT 205.3000 172.4000 205.7000 172.8000 ;
	    RECT 206.2000 171.1000 206.6000 173.5000 ;
	    RECT 208.7000 172.8000 209.0000 173.9000 ;
	    RECT 211.5000 173.8000 211.9000 173.9000 ;
	    RECT 215.0000 173.6000 215.4000 175.3000 ;
	    RECT 217.4000 174.8000 217.8000 175.6000 ;
	    RECT 218.2000 175.1000 218.5000 175.9000 ;
	    RECT 219.0000 175.1000 219.4000 175.2000 ;
	    RECT 218.2000 174.8000 219.4000 175.1000 ;
	    RECT 213.5000 173.3000 215.4000 173.6000 ;
	    RECT 213.5000 173.2000 213.9000 173.3000 ;
	    RECT 207.8000 172.1000 208.2000 172.5000 ;
	    RECT 208.6000 172.4000 209.0000 172.8000 ;
	    RECT 209.5000 172.7000 209.9000 172.8000 ;
	    RECT 209.5000 172.4000 210.9000 172.7000 ;
	    RECT 210.6000 172.1000 210.9000 172.4000 ;
	    RECT 212.6000 172.1000 213.0000 172.5000 ;
	    RECT 207.8000 171.8000 208.8000 172.1000 ;
	    RECT 208.4000 171.1000 208.8000 171.8000 ;
	    RECT 210.6000 171.1000 211.0000 172.1000 ;
	    RECT 212.6000 171.8000 213.3000 172.1000 ;
	    RECT 212.7000 171.1000 213.3000 171.8000 ;
	    RECT 215.0000 171.1000 215.4000 173.3000 ;
	    RECT 218.2000 174.2000 218.5000 174.8000 ;
	    RECT 220.6000 174.4000 221.0000 175.2000 ;
	    RECT 221.3000 174.2000 221.6000 175.9000 ;
	    RECT 222.2000 175.8000 222.6000 175.9000 ;
	    RECT 223.0000 175.8000 223.4000 176.6000 ;
	    RECT 222.2000 174.8000 222.6000 175.2000 ;
	    RECT 222.2000 174.2000 222.5000 174.8000 ;
	    RECT 218.2000 173.8000 218.6000 174.2000 ;
	    RECT 219.8000 174.1000 220.2000 174.2000 ;
	    RECT 219.8000 173.8000 220.6000 174.1000 ;
	    RECT 221.3000 173.8000 222.6000 174.2000 ;
	    RECT 223.0000 174.1000 223.4000 174.2000 ;
	    RECT 223.8000 174.1000 224.2000 179.9000 ;
	    RECT 225.4000 176.2000 225.8000 179.9000 ;
	    RECT 227.0000 176.2000 227.4000 179.9000 ;
	    RECT 225.4000 175.9000 227.4000 176.2000 ;
	    RECT 227.8000 175.9000 228.2000 179.9000 ;
	    RECT 225.8000 175.2000 226.2000 175.4000 ;
	    RECT 227.8000 175.2000 228.1000 175.9000 ;
	    RECT 228.6000 175.7000 229.0000 179.9000 ;
	    RECT 230.8000 178.2000 231.2000 179.9000 ;
	    RECT 230.2000 177.9000 231.2000 178.2000 ;
	    RECT 233.0000 177.9000 233.4000 179.9000 ;
	    RECT 235.1000 177.9000 235.7000 179.9000 ;
	    RECT 230.2000 177.5000 230.6000 177.9000 ;
	    RECT 233.0000 177.6000 233.3000 177.9000 ;
	    RECT 231.9000 177.3000 233.7000 177.6000 ;
	    RECT 235.0000 177.5000 235.4000 177.9000 ;
	    RECT 231.9000 177.2000 232.3000 177.3000 ;
	    RECT 233.3000 177.2000 233.7000 177.3000 ;
	    RECT 237.4000 177.1000 237.8000 179.9000 ;
	    RECT 238.2000 177.1000 238.6000 177.2000 ;
	    RECT 230.2000 176.5000 230.6000 176.6000 ;
	    RECT 232.5000 176.5000 232.9000 176.6000 ;
	    RECT 230.2000 176.2000 232.9000 176.5000 ;
	    RECT 233.2000 176.5000 234.3000 176.8000 ;
	    RECT 233.2000 175.9000 233.5000 176.5000 ;
	    RECT 233.9000 176.4000 234.3000 176.5000 ;
	    RECT 235.1000 176.6000 235.8000 177.0000 ;
	    RECT 237.4000 176.8000 238.6000 177.1000 ;
	    RECT 235.1000 176.1000 235.4000 176.6000 ;
	    RECT 231.1000 175.7000 233.5000 175.9000 ;
	    RECT 228.6000 175.6000 233.5000 175.7000 ;
	    RECT 234.2000 175.8000 235.4000 176.1000 ;
	    RECT 228.6000 175.5000 231.5000 175.6000 ;
	    RECT 228.6000 175.4000 231.4000 175.5000 ;
	    RECT 225.4000 174.9000 226.2000 175.2000 ;
	    RECT 227.0000 174.9000 228.2000 175.2000 ;
	    RECT 231.8000 175.1000 232.2000 175.2000 ;
	    RECT 225.4000 174.8000 225.8000 174.9000 ;
	    RECT 223.0000 173.8000 224.2000 174.1000 ;
	    RECT 218.2000 172.1000 218.5000 173.8000 ;
	    RECT 220.2000 173.6000 220.6000 173.8000 ;
	    RECT 219.0000 172.4000 219.4000 173.2000 ;
	    RECT 219.9000 173.1000 221.7000 173.3000 ;
	    RECT 222.2000 173.1000 222.5000 173.8000 ;
	    RECT 223.8000 173.1000 224.2000 173.8000 ;
	    RECT 224.6000 173.4000 225.0000 174.2000 ;
	    RECT 226.2000 173.8000 226.6000 174.6000 ;
	    RECT 219.8000 173.0000 221.8000 173.1000 ;
	    RECT 218.2000 171.1000 218.6000 172.1000 ;
	    RECT 219.8000 171.1000 220.2000 173.0000 ;
	    RECT 221.4000 171.1000 221.8000 173.0000 ;
	    RECT 222.2000 171.1000 222.6000 173.1000 ;
	    RECT 223.3000 172.8000 224.2000 173.1000 ;
	    RECT 227.0000 173.1000 227.3000 174.9000 ;
	    RECT 227.8000 174.8000 228.2000 174.9000 ;
	    RECT 229.7000 174.8000 232.2000 175.1000 ;
	    RECT 227.8000 174.2000 228.1000 174.8000 ;
	    RECT 229.7000 174.7000 230.1000 174.8000 ;
	    RECT 231.0000 174.7000 231.4000 174.8000 ;
	    RECT 230.5000 174.2000 230.9000 174.3000 ;
	    RECT 234.2000 174.2000 234.5000 175.8000 ;
	    RECT 237.4000 175.6000 237.8000 176.8000 ;
	    RECT 235.7000 175.3000 237.8000 175.6000 ;
	    RECT 235.7000 175.2000 236.1000 175.3000 ;
	    RECT 236.5000 174.9000 236.9000 175.0000 ;
	    RECT 235.0000 174.6000 236.9000 174.9000 ;
	    RECT 235.0000 174.5000 235.4000 174.6000 ;
	    RECT 227.8000 173.8000 228.2000 174.2000 ;
	    RECT 229.0000 173.9000 234.5000 174.2000 ;
	    RECT 229.0000 173.8000 229.8000 173.9000 ;
	    RECT 223.3000 171.1000 223.7000 172.8000 ;
	    RECT 227.0000 171.1000 227.4000 173.1000 ;
	    RECT 227.8000 172.8000 228.2000 173.2000 ;
	    RECT 227.7000 172.4000 228.1000 172.8000 ;
	    RECT 228.6000 171.1000 229.0000 173.5000 ;
	    RECT 231.1000 172.8000 231.4000 173.9000 ;
	    RECT 233.9000 173.8000 234.3000 173.9000 ;
	    RECT 237.4000 173.6000 237.8000 175.3000 ;
	    RECT 235.9000 173.3000 237.8000 173.6000 ;
	    RECT 238.2000 173.4000 238.6000 174.2000 ;
	    RECT 235.9000 173.2000 236.3000 173.3000 ;
	    RECT 230.2000 172.1000 230.6000 172.5000 ;
	    RECT 231.0000 172.4000 231.4000 172.8000 ;
	    RECT 231.9000 172.7000 232.3000 172.8000 ;
	    RECT 231.9000 172.4000 233.3000 172.7000 ;
	    RECT 233.0000 172.1000 233.3000 172.4000 ;
	    RECT 235.0000 172.1000 235.4000 172.5000 ;
	    RECT 230.2000 171.8000 231.2000 172.1000 ;
	    RECT 230.8000 171.1000 231.2000 171.8000 ;
	    RECT 233.0000 171.1000 233.4000 172.1000 ;
	    RECT 235.0000 171.8000 235.7000 172.1000 ;
	    RECT 235.1000 171.1000 235.7000 171.8000 ;
	    RECT 237.4000 171.1000 237.8000 173.3000 ;
	    RECT 239.0000 173.1000 239.4000 179.9000 ;
	    RECT 239.8000 175.8000 240.2000 176.6000 ;
	    RECT 241.9000 176.3000 242.3000 179.9000 ;
	    RECT 241.4000 175.9000 242.3000 176.3000 ;
	    RECT 241.5000 174.2000 241.8000 175.9000 ;
	    RECT 242.2000 175.1000 242.6000 175.6000 ;
	    RECT 243.0000 175.1000 243.4000 175.2000 ;
	    RECT 242.2000 174.8000 243.4000 175.1000 ;
	    RECT 243.8000 175.1000 244.2000 179.9000 ;
	    RECT 244.9000 176.3000 245.3000 179.9000 ;
	    RECT 247.3000 176.3000 247.7000 179.9000 ;
	    RECT 250.2000 177.9000 250.6000 179.9000 ;
	    RECT 244.9000 175.9000 245.8000 176.3000 ;
	    RECT 247.3000 175.9000 248.2000 176.3000 ;
	    RECT 244.6000 175.1000 245.0000 175.6000 ;
	    RECT 243.8000 174.8000 245.0000 175.1000 ;
	    RECT 241.4000 173.8000 241.8000 174.2000 ;
	    RECT 239.0000 172.8000 239.9000 173.1000 ;
	    RECT 239.5000 172.2000 239.9000 172.8000 ;
	    RECT 240.6000 172.4000 241.0000 173.2000 ;
	    RECT 241.5000 173.1000 241.8000 173.8000 ;
	    RECT 242.2000 173.8000 242.6000 174.2000 ;
	    RECT 242.2000 173.1000 242.5000 173.8000 ;
	    RECT 241.4000 172.8000 242.5000 173.1000 ;
	    RECT 239.5000 171.8000 240.2000 172.2000 ;
	    RECT 241.5000 172.1000 241.8000 172.8000 ;
	    RECT 243.0000 172.4000 243.4000 173.2000 ;
	    RECT 239.5000 171.1000 239.9000 171.8000 ;
	    RECT 241.4000 171.1000 241.8000 172.1000 ;
	    RECT 243.8000 171.1000 244.2000 174.8000 ;
	    RECT 245.4000 174.2000 245.7000 175.9000 ;
	    RECT 247.0000 174.8000 247.4000 175.6000 ;
	    RECT 247.8000 174.2000 248.1000 175.9000 ;
	    RECT 250.3000 175.8000 250.6000 177.9000 ;
	    RECT 251.8000 175.9000 252.2000 179.9000 ;
	    RECT 252.9000 176.3000 253.3000 179.9000 ;
	    RECT 252.9000 175.9000 253.8000 176.3000 ;
	    RECT 250.3000 175.5000 251.5000 175.8000 ;
	    RECT 250.2000 174.8000 250.6000 175.2000 ;
	    RECT 245.4000 173.8000 245.8000 174.2000 ;
	    RECT 247.8000 173.8000 248.2000 174.2000 ;
	    RECT 249.4000 173.8000 249.8000 174.6000 ;
	    RECT 250.3000 174.4000 250.6000 174.8000 ;
	    RECT 250.2000 174.0000 250.8000 174.4000 ;
	    RECT 251.2000 173.8000 251.5000 175.5000 ;
	    RECT 251.9000 175.2000 252.2000 175.9000 ;
	    RECT 251.8000 174.8000 252.2000 175.2000 ;
	    RECT 252.6000 174.8000 253.0000 175.6000 ;
	    RECT 253.4000 175.1000 253.7000 175.9000 ;
	    RECT 253.4000 174.8000 255.3000 175.1000 ;
	    RECT 245.4000 172.2000 245.7000 173.8000 ;
	    RECT 246.2000 172.4000 246.6000 173.2000 ;
	    RECT 247.8000 172.2000 248.1000 173.8000 ;
	    RECT 251.2000 173.7000 251.6000 173.8000 ;
	    RECT 250.1000 173.5000 251.6000 173.7000 ;
	    RECT 249.5000 173.4000 251.6000 173.5000 ;
	    RECT 249.5000 173.2000 250.4000 173.4000 ;
	    RECT 248.6000 172.4000 249.0000 173.2000 ;
	    RECT 249.5000 173.1000 249.8000 173.2000 ;
	    RECT 251.9000 173.1000 252.2000 174.8000 ;
	    RECT 245.4000 171.1000 245.8000 172.2000 ;
	    RECT 247.8000 171.1000 248.2000 172.2000 ;
	    RECT 249.4000 171.1000 249.8000 173.1000 ;
	    RECT 251.5000 172.6000 252.2000 173.1000 ;
	    RECT 253.4000 174.2000 253.7000 174.8000 ;
	    RECT 255.0000 174.2000 255.3000 174.8000 ;
	    RECT 253.4000 173.8000 253.8000 174.2000 ;
	    RECT 255.0000 173.8000 255.4000 174.2000 ;
	    RECT 251.5000 172.2000 251.9000 172.6000 ;
	    RECT 251.5000 171.8000 252.2000 172.2000 ;
	    RECT 253.4000 172.1000 253.7000 173.8000 ;
	    RECT 254.2000 172.4000 254.6000 173.2000 ;
	    RECT 251.5000 171.1000 251.9000 171.8000 ;
	    RECT 253.4000 171.1000 253.8000 172.1000 ;
	    RECT 255.8000 171.1000 256.2000 179.9000 ;
	    RECT 256.6000 175.7000 257.0000 179.9000 ;
	    RECT 258.8000 178.2000 259.2000 179.9000 ;
	    RECT 258.2000 177.9000 259.2000 178.2000 ;
	    RECT 261.0000 177.9000 261.4000 179.9000 ;
	    RECT 263.1000 177.9000 263.7000 179.9000 ;
	    RECT 258.2000 177.5000 258.6000 177.9000 ;
	    RECT 261.0000 177.6000 261.3000 177.9000 ;
	    RECT 259.9000 177.3000 261.7000 177.6000 ;
	    RECT 263.0000 177.5000 263.4000 177.9000 ;
	    RECT 259.9000 177.2000 260.3000 177.3000 ;
	    RECT 261.3000 177.2000 261.7000 177.3000 ;
	    RECT 258.2000 176.5000 258.6000 176.6000 ;
	    RECT 260.5000 176.5000 260.9000 176.6000 ;
	    RECT 258.2000 176.2000 260.9000 176.5000 ;
	    RECT 261.2000 176.5000 262.3000 176.8000 ;
	    RECT 261.2000 175.9000 261.5000 176.5000 ;
	    RECT 261.9000 176.4000 262.3000 176.5000 ;
	    RECT 263.1000 176.6000 263.8000 177.0000 ;
	    RECT 263.1000 176.1000 263.4000 176.6000 ;
	    RECT 259.1000 175.7000 261.5000 175.9000 ;
	    RECT 256.6000 175.6000 261.5000 175.7000 ;
	    RECT 262.2000 175.8000 263.4000 176.1000 ;
	    RECT 256.6000 175.5000 259.5000 175.6000 ;
	    RECT 256.6000 175.4000 259.4000 175.5000 ;
	    RECT 259.8000 175.1000 260.2000 175.2000 ;
	    RECT 257.7000 174.8000 260.2000 175.1000 ;
	    RECT 257.7000 174.7000 258.1000 174.8000 ;
	    RECT 259.0000 174.7000 259.4000 174.8000 ;
	    RECT 258.5000 174.2000 258.9000 174.3000 ;
	    RECT 262.2000 174.2000 262.5000 175.8000 ;
	    RECT 265.4000 175.6000 265.8000 179.9000 ;
	    RECT 263.7000 175.3000 265.8000 175.6000 ;
	    RECT 263.7000 175.2000 264.1000 175.3000 ;
	    RECT 264.5000 174.9000 264.9000 175.0000 ;
	    RECT 263.0000 174.6000 264.9000 174.9000 ;
	    RECT 263.0000 174.5000 263.4000 174.6000 ;
	    RECT 257.0000 173.9000 262.5000 174.2000 ;
	    RECT 257.0000 173.8000 257.8000 173.9000 ;
	    RECT 256.6000 171.1000 257.0000 173.5000 ;
	    RECT 259.1000 172.8000 259.4000 173.9000 ;
	    RECT 261.9000 173.8000 262.3000 173.9000 ;
	    RECT 265.4000 173.6000 265.8000 175.3000 ;
	    RECT 263.9000 173.3000 265.8000 173.6000 ;
	    RECT 263.9000 173.2000 264.3000 173.3000 ;
	    RECT 258.2000 172.1000 258.6000 172.5000 ;
	    RECT 259.0000 172.4000 259.4000 172.8000 ;
	    RECT 259.9000 172.7000 260.3000 172.8000 ;
	    RECT 259.9000 172.4000 261.3000 172.7000 ;
	    RECT 261.0000 172.1000 261.3000 172.4000 ;
	    RECT 263.0000 172.1000 263.4000 172.5000 ;
	    RECT 258.2000 171.8000 259.2000 172.1000 ;
	    RECT 258.8000 171.1000 259.2000 171.8000 ;
	    RECT 261.0000 171.1000 261.4000 172.1000 ;
	    RECT 263.0000 171.8000 263.7000 172.1000 ;
	    RECT 263.1000 171.1000 263.7000 171.8000 ;
	    RECT 265.4000 171.1000 265.8000 173.3000 ;
	    RECT 266.2000 176.1000 266.6000 179.9000 ;
	    RECT 267.8000 176.2000 268.2000 179.9000 ;
	    RECT 267.0000 176.1000 267.4000 176.2000 ;
	    RECT 266.2000 175.8000 267.4000 176.1000 ;
	    RECT 267.8000 175.9000 268.9000 176.2000 ;
	    RECT 266.2000 171.1000 266.6000 175.8000 ;
	    RECT 268.6000 175.6000 268.9000 175.9000 ;
	    RECT 268.6000 175.2000 269.2000 175.6000 ;
	    RECT 267.0000 175.1000 267.4000 175.2000 ;
	    RECT 267.8000 175.1000 268.2000 175.2000 ;
	    RECT 267.0000 174.8000 268.2000 175.1000 ;
	    RECT 267.8000 174.4000 268.2000 174.8000 ;
	    RECT 268.6000 173.7000 268.9000 175.2000 ;
	    RECT 267.8000 173.4000 268.9000 173.7000 ;
	    RECT 267.0000 172.4000 267.4000 173.2000 ;
	    RECT 267.8000 171.1000 268.2000 173.4000 ;
	    RECT 0.6000 167.6000 1.0000 169.9000 ;
	    RECT 0.6000 167.3000 1.7000 167.6000 ;
	    RECT 1.4000 165.8000 1.7000 167.3000 ;
	    RECT 2.2000 166.2000 2.6000 169.9000 ;
	    RECT 3.0000 167.9000 3.4000 169.9000 ;
	    RECT 3.8000 168.0000 4.2000 169.9000 ;
	    RECT 5.4000 168.0000 5.8000 169.9000 ;
	    RECT 3.8000 167.9000 5.8000 168.0000 ;
	    RECT 3.1000 167.2000 3.4000 167.9000 ;
	    RECT 3.9000 167.7000 5.7000 167.9000 ;
	    RECT 5.0000 167.2000 5.4000 167.4000 ;
	    RECT 3.0000 166.8000 4.3000 167.2000 ;
	    RECT 5.0000 167.1000 5.8000 167.2000 ;
	    RECT 7.0000 167.1000 7.4000 169.9000 ;
	    RECT 5.0000 166.9000 7.4000 167.1000 ;
	    RECT 9.6000 167.1000 10.0000 169.9000 ;
	    RECT 12.5000 167.9000 13.3000 169.9000 ;
	    RECT 9.6000 166.9000 10.5000 167.1000 ;
	    RECT 5.4000 166.8000 7.4000 166.9000 ;
	    RECT 9.7000 166.8000 10.5000 166.9000 ;
	    RECT 1.4000 165.4000 2.0000 165.8000 ;
	    RECT 1.4000 165.1000 1.7000 165.4000 ;
	    RECT 2.3000 165.1000 2.6000 166.2000 ;
	    RECT 0.6000 164.8000 1.7000 165.1000 ;
	    RECT 0.6000 161.1000 1.0000 164.8000 ;
	    RECT 2.2000 161.1000 2.6000 165.1000 ;
	    RECT 3.0000 165.1000 3.4000 165.2000 ;
	    RECT 4.0000 165.1000 4.3000 166.8000 ;
	    RECT 3.0000 164.8000 3.7000 165.1000 ;
	    RECT 4.0000 164.8000 4.5000 165.1000 ;
	    RECT 3.4000 164.2000 3.7000 164.8000 ;
	    RECT 3.4000 163.8000 3.8000 164.2000 ;
	    RECT 4.1000 162.2000 4.5000 164.8000 ;
	    RECT 4.1000 161.8000 5.0000 162.2000 ;
	    RECT 4.1000 161.1000 4.5000 161.8000 ;
	    RECT 7.0000 161.1000 7.4000 166.8000 ;
	    RECT 8.6000 165.8000 9.4000 166.2000 ;
	    RECT 7.8000 164.8000 8.2000 165.6000 ;
	    RECT 10.2000 165.2000 10.5000 166.8000 ;
	    RECT 12.7000 166.2000 13.0000 167.9000 ;
	    RECT 13.4000 167.1000 13.8000 167.2000 ;
	    RECT 15.0000 167.1000 15.4000 169.9000 ;
	    RECT 13.4000 166.8000 15.4000 167.1000 ;
	    RECT 13.4000 166.6000 13.7000 166.8000 ;
	    RECT 13.3000 166.2000 13.7000 166.6000 ;
	    RECT 11.0000 166.1000 11.4000 166.2000 ;
	    RECT 11.0000 165.8000 11.8000 166.1000 ;
	    RECT 12.6000 165.8000 13.0000 166.2000 ;
	    RECT 11.4000 165.6000 11.8000 165.8000 ;
	    RECT 12.7000 165.7000 13.0000 165.8000 ;
	    RECT 12.7000 165.4000 13.7000 165.7000 ;
	    RECT 10.2000 164.8000 10.6000 165.2000 ;
	    RECT 13.4000 165.1000 13.7000 165.4000 ;
	    RECT 11.0000 164.8000 13.0000 165.1000 ;
	    RECT 9.4000 163.8000 9.8000 164.6000 ;
	    RECT 10.2000 163.5000 10.5000 164.8000 ;
	    RECT 8.7000 163.2000 10.5000 163.5000 ;
	    RECT 8.7000 163.1000 9.0000 163.2000 ;
	    RECT 8.6000 161.1000 9.0000 163.1000 ;
	    RECT 10.2000 163.1000 10.5000 163.2000 ;
	    RECT 10.2000 161.1000 10.6000 163.1000 ;
	    RECT 11.0000 161.1000 11.4000 164.8000 ;
	    RECT 12.6000 161.4000 13.0000 164.8000 ;
	    RECT 13.4000 161.7000 13.8000 165.1000 ;
	    RECT 14.2000 161.4000 14.6000 165.1000 ;
	    RECT 12.6000 161.1000 14.6000 161.4000 ;
	    RECT 15.0000 161.1000 15.4000 166.8000 ;
	    RECT 16.6000 161.1000 17.0000 169.9000 ;
	    RECT 19.0000 167.1000 19.4000 169.9000 ;
	    RECT 21.1000 167.9000 21.9000 169.9000 ;
	    RECT 24.6000 168.9000 25.0000 169.9000 ;
	    RECT 20.6000 167.1000 21.0000 167.2000 ;
	    RECT 19.0000 166.8000 21.0000 167.1000 ;
	    RECT 19.0000 161.1000 19.4000 166.8000 ;
	    RECT 20.7000 166.6000 21.0000 166.8000 ;
	    RECT 20.7000 166.2000 21.1000 166.6000 ;
	    RECT 21.4000 166.2000 21.7000 167.9000 ;
	    RECT 24.7000 167.2000 25.0000 168.9000 ;
	    RECT 24.6000 166.8000 25.0000 167.2000 ;
	    RECT 21.4000 165.8000 21.8000 166.2000 ;
	    RECT 23.0000 166.1000 23.4000 166.2000 ;
	    RECT 22.6000 165.8000 23.4000 166.1000 ;
	    RECT 21.4000 165.7000 21.7000 165.8000 ;
	    RECT 20.7000 165.4000 21.7000 165.7000 ;
	    RECT 22.6000 165.6000 23.0000 165.8000 ;
	    RECT 20.7000 165.1000 21.0000 165.4000 ;
	    RECT 24.7000 165.1000 25.0000 166.8000 ;
	    RECT 25.4000 166.8000 25.8000 167.2000 ;
	    RECT 25.4000 166.2000 25.7000 166.8000 ;
	    RECT 25.4000 166.1000 25.8000 166.2000 ;
	    RECT 26.2000 166.1000 26.6000 169.9000 ;
	    RECT 29.6000 167.1000 30.0000 169.9000 ;
	    RECT 29.6000 166.9000 30.5000 167.1000 ;
	    RECT 29.7000 166.8000 30.5000 166.9000 ;
	    RECT 25.4000 165.8000 26.6000 166.1000 ;
	    RECT 28.6000 165.8000 29.4000 166.2000 ;
	    RECT 25.4000 165.4000 25.8000 165.8000 ;
	    RECT 19.8000 161.4000 20.2000 165.1000 ;
	    RECT 20.6000 161.7000 21.0000 165.1000 ;
	    RECT 21.4000 164.8000 23.4000 165.1000 ;
	    RECT 21.4000 161.4000 21.8000 164.8000 ;
	    RECT 19.8000 161.1000 21.8000 161.4000 ;
	    RECT 23.0000 161.1000 23.4000 164.8000 ;
	    RECT 24.6000 164.7000 25.5000 165.1000 ;
	    RECT 25.1000 162.2000 25.5000 164.7000 ;
	    RECT 24.6000 161.8000 25.5000 162.2000 ;
	    RECT 25.1000 161.1000 25.5000 161.8000 ;
	    RECT 26.2000 161.1000 26.6000 165.8000 ;
	    RECT 27.8000 164.8000 28.2000 165.6000 ;
	    RECT 30.2000 165.2000 30.5000 166.8000 ;
	    RECT 30.2000 164.8000 30.6000 165.2000 ;
	    RECT 31.8000 165.1000 32.2000 169.9000 ;
	    RECT 32.9000 168.2000 33.3000 169.9000 ;
	    RECT 32.9000 167.9000 33.8000 168.2000 ;
	    RECT 35.0000 168.0000 35.4000 169.9000 ;
	    RECT 36.6000 168.0000 37.0000 169.9000 ;
	    RECT 35.0000 167.9000 37.0000 168.0000 ;
	    RECT 37.4000 167.9000 37.8000 169.9000 ;
	    RECT 32.6000 166.8000 33.0000 167.2000 ;
	    RECT 32.6000 166.1000 32.9000 166.8000 ;
	    RECT 33.4000 166.1000 33.8000 167.9000 ;
	    RECT 35.1000 167.7000 36.9000 167.9000 ;
	    RECT 35.4000 167.2000 35.8000 167.4000 ;
	    RECT 37.4000 167.2000 37.7000 167.9000 ;
	    RECT 35.0000 166.9000 35.8000 167.2000 ;
	    RECT 35.0000 166.8000 35.4000 166.9000 ;
	    RECT 36.5000 166.8000 37.8000 167.2000 ;
	    RECT 32.6000 165.8000 33.8000 166.1000 ;
	    RECT 34.2000 166.1000 34.6000 166.2000 ;
	    RECT 35.8000 166.1000 36.2000 166.6000 ;
	    RECT 34.2000 165.8000 36.2000 166.1000 ;
	    RECT 32.6000 165.1000 33.0000 165.2000 ;
	    RECT 31.8000 164.8000 33.0000 165.1000 ;
	    RECT 27.0000 164.1000 27.4000 164.2000 ;
	    RECT 29.4000 164.1000 29.8000 164.6000 ;
	    RECT 27.0000 163.8000 29.8000 164.1000 ;
	    RECT 30.2000 163.5000 30.5000 164.8000 ;
	    RECT 28.7000 163.2000 30.5000 163.5000 ;
	    RECT 28.7000 163.1000 29.0000 163.2000 ;
	    RECT 28.6000 161.1000 29.0000 163.1000 ;
	    RECT 30.2000 163.1000 30.5000 163.2000 ;
	    RECT 30.2000 161.1000 30.6000 163.1000 ;
	    RECT 31.8000 161.1000 32.2000 164.8000 ;
	    RECT 32.6000 164.4000 33.0000 164.8000 ;
	    RECT 33.4000 161.1000 33.8000 165.8000 ;
	    RECT 36.5000 165.1000 36.8000 166.8000 ;
	    RECT 37.4000 165.1000 37.8000 165.2000 ;
	    RECT 36.3000 164.8000 36.8000 165.1000 ;
	    RECT 37.1000 164.8000 37.8000 165.1000 ;
	    RECT 36.3000 162.2000 36.7000 164.8000 ;
	    RECT 37.1000 164.2000 37.4000 164.8000 ;
	    RECT 37.0000 163.8000 37.4000 164.2000 ;
	    RECT 35.8000 161.8000 36.7000 162.2000 ;
	    RECT 36.3000 161.1000 36.7000 161.8000 ;
	    RECT 39.0000 161.1000 39.4000 169.9000 ;
	    RECT 40.6000 161.1000 41.0000 169.9000 ;
	    RECT 42.0000 167.2000 42.4000 169.9000 ;
	    RECT 41.4000 166.9000 42.4000 167.2000 ;
	    RECT 41.4000 166.8000 42.3000 166.9000 ;
	    RECT 41.5000 165.2000 41.8000 166.8000 ;
	    RECT 42.6000 165.8000 43.4000 166.2000 ;
	    RECT 45.4000 166.1000 45.8000 169.9000 ;
	    RECT 47.5000 167.9000 48.3000 169.9000 ;
	    RECT 47.8000 166.2000 48.1000 167.9000 ;
	    RECT 46.2000 166.1000 46.6000 166.2000 ;
	    RECT 45.4000 165.8000 46.6000 166.1000 ;
	    RECT 41.4000 164.8000 41.8000 165.2000 ;
	    RECT 43.8000 164.8000 44.2000 165.6000 ;
	    RECT 41.5000 163.5000 41.8000 164.8000 ;
	    RECT 42.2000 163.8000 42.6000 164.6000 ;
	    RECT 41.5000 163.2000 43.3000 163.5000 ;
	    RECT 41.5000 163.1000 41.8000 163.2000 ;
	    RECT 41.4000 161.1000 41.8000 163.1000 ;
	    RECT 43.0000 163.1000 43.3000 163.2000 ;
	    RECT 43.0000 161.1000 43.4000 163.1000 ;
	    RECT 45.4000 161.1000 45.8000 165.8000 ;
	    RECT 46.2000 165.4000 46.6000 165.8000 ;
	    RECT 47.8000 165.8000 48.2000 166.2000 ;
	    RECT 49.4000 166.1000 49.8000 166.2000 ;
	    RECT 51.0000 166.1000 51.4000 169.9000 ;
	    RECT 51.9000 168.2000 52.3000 168.6000 ;
	    RECT 51.8000 167.8000 52.2000 168.2000 ;
	    RECT 52.6000 167.9000 53.0000 169.9000 ;
	    RECT 51.8000 167.1000 52.2000 167.2000 ;
	    RECT 52.7000 167.1000 53.0000 167.9000 ;
	    RECT 51.8000 166.8000 53.0000 167.1000 ;
	    RECT 49.0000 165.8000 51.4000 166.1000 ;
	    RECT 51.8000 166.1000 52.2000 166.2000 ;
	    RECT 52.7000 166.1000 53.0000 166.8000 ;
	    RECT 55.8000 168.9000 56.2000 169.9000 ;
	    RECT 55.8000 167.2000 56.1000 168.9000 ;
	    RECT 56.6000 167.8000 57.0000 168.6000 ;
	    RECT 59.0000 168.0000 59.4000 169.9000 ;
	    RECT 60.6000 168.0000 61.0000 169.9000 ;
	    RECT 59.0000 167.9000 61.0000 168.0000 ;
	    RECT 61.4000 167.9000 61.8000 169.9000 ;
	    RECT 59.1000 167.7000 60.9000 167.9000 ;
	    RECT 59.4000 167.2000 59.8000 167.4000 ;
	    RECT 61.4000 167.2000 61.7000 167.9000 ;
	    RECT 62.2000 167.8000 62.6000 168.6000 ;
	    RECT 55.8000 166.8000 56.2000 167.2000 ;
	    RECT 58.2000 167.1000 58.6000 167.2000 ;
	    RECT 59.0000 167.1000 59.8000 167.2000 ;
	    RECT 58.2000 166.9000 59.8000 167.1000 ;
	    RECT 58.2000 166.8000 59.4000 166.9000 ;
	    RECT 60.5000 166.8000 61.8000 167.2000 ;
	    RECT 54.2000 166.1000 54.6000 166.2000 ;
	    RECT 51.8000 165.8000 53.0000 166.1000 ;
	    RECT 53.8000 165.8000 54.6000 166.1000 ;
	    RECT 47.8000 165.7000 48.1000 165.8000 ;
	    RECT 47.1000 165.4000 48.1000 165.7000 ;
	    RECT 49.0000 165.6000 49.4000 165.8000 ;
	    RECT 47.1000 165.1000 47.4000 165.4000 ;
	    RECT 46.2000 161.4000 46.6000 165.1000 ;
	    RECT 47.0000 161.7000 47.4000 165.1000 ;
	    RECT 47.8000 164.8000 49.8000 165.1000 ;
	    RECT 47.8000 161.4000 48.2000 164.8000 ;
	    RECT 46.2000 161.1000 48.2000 161.4000 ;
	    RECT 49.4000 161.1000 49.8000 164.8000 ;
	    RECT 51.0000 161.1000 51.4000 165.8000 ;
	    RECT 51.9000 165.1000 52.2000 165.8000 ;
	    RECT 53.8000 165.6000 54.2000 165.8000 ;
	    RECT 55.0000 165.4000 55.4000 166.2000 ;
	    RECT 55.8000 165.1000 56.1000 166.8000 ;
	    RECT 60.5000 165.1000 60.8000 166.8000 ;
	    RECT 63.0000 166.1000 63.4000 169.9000 ;
	    RECT 65.4000 167.9000 65.8000 169.9000 ;
	    RECT 66.1000 168.2000 66.5000 168.6000 ;
	    RECT 67.1000 168.2000 67.5000 168.6000 ;
	    RECT 66.2000 168.1000 66.6000 168.2000 ;
	    RECT 67.0000 168.1000 67.4000 168.2000 ;
	    RECT 64.6000 166.4000 65.0000 167.2000 ;
	    RECT 63.8000 166.1000 64.2000 166.2000 ;
	    RECT 65.4000 166.1000 65.7000 167.9000 ;
	    RECT 66.2000 167.8000 67.4000 168.1000 ;
	    RECT 67.8000 167.9000 68.2000 169.9000 ;
	    RECT 66.2000 166.1000 66.6000 166.2000 ;
	    RECT 63.0000 165.8000 64.6000 166.1000 ;
	    RECT 65.4000 165.8000 66.6000 166.1000 ;
	    RECT 67.0000 166.1000 67.4000 166.2000 ;
	    RECT 67.9000 166.1000 68.2000 167.9000 ;
	    RECT 68.6000 166.4000 69.0000 167.2000 ;
	    RECT 69.4000 166.1000 69.8000 166.2000 ;
	    RECT 70.2000 166.1000 70.6000 169.9000 ;
	    RECT 71.0000 167.8000 71.4000 168.6000 ;
	    RECT 71.9000 168.2000 72.3000 168.6000 ;
	    RECT 71.8000 167.8000 72.2000 168.2000 ;
	    RECT 72.6000 167.9000 73.0000 169.9000 ;
	    RECT 72.7000 166.2000 73.0000 167.9000 ;
	    RECT 73.4000 166.4000 73.8000 167.2000 ;
	    RECT 67.0000 165.8000 68.2000 166.1000 ;
	    RECT 69.0000 165.8000 70.6000 166.1000 ;
	    RECT 71.8000 166.1000 72.2000 166.2000 ;
	    RECT 72.6000 166.1000 73.0000 166.2000 ;
	    RECT 74.2000 166.1000 74.6000 166.2000 ;
	    RECT 75.0000 166.1000 75.4000 169.9000 ;
	    RECT 75.8000 168.1000 76.2000 168.6000 ;
	    RECT 76.6000 168.1000 77.0000 169.9000 ;
	    RECT 78.7000 169.2000 79.3000 169.9000 ;
	    RECT 78.7000 168.9000 79.4000 169.2000 ;
	    RECT 81.0000 168.9000 81.4000 169.9000 ;
	    RECT 83.2000 169.2000 83.6000 169.9000 ;
	    RECT 83.2000 168.9000 84.2000 169.2000 ;
	    RECT 79.0000 168.5000 79.4000 168.9000 ;
	    RECT 81.1000 168.6000 81.4000 168.9000 ;
	    RECT 81.1000 168.3000 82.5000 168.6000 ;
	    RECT 82.1000 168.2000 82.5000 168.3000 ;
	    RECT 83.0000 168.2000 83.4000 168.6000 ;
	    RECT 83.8000 168.5000 84.2000 168.9000 ;
	    RECT 75.8000 167.8000 77.0000 168.1000 ;
	    RECT 71.8000 165.8000 73.0000 166.1000 ;
	    RECT 73.8000 165.8000 75.4000 166.1000 ;
	    RECT 61.4000 165.1000 61.8000 165.2000 ;
	    RECT 51.8000 161.1000 52.2000 165.1000 ;
	    RECT 52.6000 164.8000 54.6000 165.1000 ;
	    RECT 52.6000 161.1000 53.0000 164.8000 ;
	    RECT 54.2000 161.1000 54.6000 164.8000 ;
	    RECT 55.3000 164.7000 56.2000 165.1000 ;
	    RECT 60.3000 164.8000 60.8000 165.1000 ;
	    RECT 61.1000 164.8000 61.8000 165.1000 ;
	    RECT 55.3000 164.2000 55.7000 164.7000 ;
	    RECT 55.0000 163.8000 55.7000 164.2000 ;
	    RECT 55.3000 161.1000 55.7000 163.8000 ;
	    RECT 60.3000 161.1000 60.7000 164.8000 ;
	    RECT 61.1000 164.2000 61.4000 164.8000 ;
	    RECT 61.0000 163.8000 61.4000 164.2000 ;
	    RECT 63.0000 161.1000 63.4000 165.8000 ;
	    RECT 64.2000 165.6000 64.6000 165.8000 ;
	    RECT 66.2000 165.1000 66.5000 165.8000 ;
	    RECT 67.1000 165.1000 67.4000 165.8000 ;
	    RECT 69.0000 165.6000 69.4000 165.8000 ;
	    RECT 63.8000 164.8000 65.8000 165.1000 ;
	    RECT 63.8000 161.1000 64.2000 164.8000 ;
	    RECT 65.4000 161.1000 65.8000 164.8000 ;
	    RECT 66.2000 161.1000 66.6000 165.1000 ;
	    RECT 67.0000 161.1000 67.4000 165.1000 ;
	    RECT 67.8000 164.8000 69.8000 165.1000 ;
	    RECT 67.8000 161.1000 68.2000 164.8000 ;
	    RECT 69.4000 161.1000 69.8000 164.8000 ;
	    RECT 70.2000 161.1000 70.6000 165.8000 ;
	    RECT 71.9000 165.1000 72.2000 165.8000 ;
	    RECT 73.8000 165.6000 74.2000 165.8000 ;
	    RECT 71.8000 161.1000 72.2000 165.1000 ;
	    RECT 72.6000 164.8000 74.6000 165.1000 ;
	    RECT 72.6000 161.1000 73.0000 164.8000 ;
	    RECT 74.2000 161.1000 74.6000 164.8000 ;
	    RECT 75.0000 161.1000 75.4000 165.8000 ;
	    RECT 76.6000 167.7000 77.0000 167.8000 ;
	    RECT 78.1000 167.7000 78.5000 167.8000 ;
	    RECT 76.6000 167.4000 78.5000 167.7000 ;
	    RECT 76.6000 165.7000 77.0000 167.4000 ;
	    RECT 77.4000 166.8000 77.8000 167.4000 ;
	    RECT 80.1000 167.1000 80.5000 167.2000 ;
	    RECT 82.2000 167.1000 82.6000 167.2000 ;
	    RECT 83.0000 167.1000 83.3000 168.2000 ;
	    RECT 85.4000 167.5000 85.8000 169.9000 ;
	    RECT 86.2000 167.5000 86.6000 169.9000 ;
	    RECT 88.4000 169.2000 88.8000 169.9000 ;
	    RECT 87.8000 168.9000 88.8000 169.2000 ;
	    RECT 90.6000 168.9000 91.0000 169.9000 ;
	    RECT 92.7000 169.2000 93.3000 169.9000 ;
	    RECT 92.6000 168.9000 93.3000 169.2000 ;
	    RECT 87.8000 168.5000 88.2000 168.9000 ;
	    RECT 90.6000 168.6000 90.9000 168.9000 ;
	    RECT 88.6000 168.2000 89.0000 168.6000 ;
	    RECT 89.5000 168.3000 90.9000 168.6000 ;
	    RECT 92.6000 168.5000 93.0000 168.9000 ;
	    RECT 89.5000 168.2000 89.9000 168.3000 ;
	    RECT 84.6000 167.1000 85.4000 167.2000 ;
	    RECT 86.6000 167.1000 87.4000 167.2000 ;
	    RECT 88.7000 167.1000 89.0000 168.2000 ;
	    RECT 95.0000 168.1000 95.4000 169.9000 ;
	    RECT 95.8000 168.1000 96.2000 168.6000 ;
	    RECT 95.0000 167.8000 96.2000 168.1000 ;
	    RECT 96.6000 168.1000 97.0000 169.9000 ;
	    RECT 98.2000 168.9000 98.6000 169.9000 ;
	    RECT 97.4000 168.1000 97.8000 168.6000 ;
	    RECT 96.6000 167.8000 97.8000 168.1000 ;
	    RECT 93.5000 167.7000 93.9000 167.8000 ;
	    RECT 95.0000 167.7000 95.4000 167.8000 ;
	    RECT 93.5000 167.4000 95.4000 167.7000 ;
	    RECT 91.5000 167.1000 91.9000 167.2000 ;
	    RECT 79.9000 166.8000 92.1000 167.1000 ;
	    RECT 79.0000 166.4000 79.4000 166.5000 ;
	    RECT 77.5000 166.1000 79.4000 166.4000 ;
	    RECT 77.5000 166.0000 77.9000 166.1000 ;
	    RECT 78.3000 165.7000 78.7000 165.8000 ;
	    RECT 76.6000 165.4000 78.7000 165.7000 ;
	    RECT 76.6000 161.1000 77.0000 165.4000 ;
	    RECT 79.9000 165.2000 80.2000 166.8000 ;
	    RECT 83.5000 166.7000 83.9000 166.8000 ;
	    RECT 88.1000 166.7000 88.5000 166.8000 ;
	    RECT 84.3000 166.2000 84.7000 166.3000 ;
	    RECT 81.4000 166.1000 81.8000 166.2000 ;
	    RECT 82.2000 166.1000 84.7000 166.2000 ;
	    RECT 81.4000 165.9000 84.7000 166.1000 ;
	    RECT 87.3000 166.2000 87.7000 166.3000 ;
	    RECT 91.8000 166.2000 92.1000 166.8000 ;
	    RECT 92.6000 166.4000 93.0000 166.5000 ;
	    RECT 87.3000 165.9000 89.8000 166.2000 ;
	    RECT 81.4000 165.8000 82.6000 165.9000 ;
	    RECT 89.4000 165.8000 89.8000 165.9000 ;
	    RECT 91.8000 165.8000 92.2000 166.2000 ;
	    RECT 92.6000 166.1000 94.5000 166.4000 ;
	    RECT 94.1000 166.0000 94.5000 166.1000 ;
	    RECT 83.0000 165.5000 85.8000 165.6000 ;
	    RECT 82.9000 165.4000 85.8000 165.5000 ;
	    RECT 79.0000 164.9000 80.2000 165.2000 ;
	    RECT 80.9000 165.3000 85.8000 165.4000 ;
	    RECT 80.9000 165.1000 83.3000 165.3000 ;
	    RECT 79.0000 164.4000 79.3000 164.9000 ;
	    RECT 78.6000 164.0000 79.3000 164.4000 ;
	    RECT 80.1000 164.5000 80.5000 164.6000 ;
	    RECT 80.9000 164.5000 81.2000 165.1000 ;
	    RECT 80.1000 164.2000 81.2000 164.5000 ;
	    RECT 81.5000 164.5000 84.2000 164.8000 ;
	    RECT 81.5000 164.4000 81.9000 164.5000 ;
	    RECT 83.8000 164.4000 84.2000 164.5000 ;
	    RECT 80.7000 163.7000 81.1000 163.8000 ;
	    RECT 82.1000 163.7000 82.5000 163.8000 ;
	    RECT 79.0000 163.1000 79.4000 163.5000 ;
	    RECT 80.7000 163.4000 82.5000 163.7000 ;
	    RECT 81.1000 163.1000 81.4000 163.4000 ;
	    RECT 83.8000 163.1000 84.2000 163.5000 ;
	    RECT 78.7000 161.1000 79.3000 163.1000 ;
	    RECT 81.0000 161.1000 81.4000 163.1000 ;
	    RECT 83.2000 162.8000 84.2000 163.1000 ;
	    RECT 83.2000 161.1000 83.6000 162.8000 ;
	    RECT 85.4000 161.1000 85.8000 165.3000 ;
	    RECT 86.2000 165.5000 89.0000 165.6000 ;
	    RECT 86.2000 165.4000 89.1000 165.5000 ;
	    RECT 86.2000 165.3000 91.1000 165.4000 ;
	    RECT 86.2000 161.1000 86.6000 165.3000 ;
	    RECT 88.7000 165.1000 91.1000 165.3000 ;
	    RECT 87.8000 164.5000 90.5000 164.8000 ;
	    RECT 87.8000 164.4000 88.2000 164.5000 ;
	    RECT 90.1000 164.4000 90.5000 164.5000 ;
	    RECT 90.8000 164.5000 91.1000 165.1000 ;
	    RECT 91.8000 165.2000 92.1000 165.8000 ;
	    RECT 93.3000 165.7000 93.7000 165.8000 ;
	    RECT 95.0000 165.7000 95.4000 167.4000 ;
	    RECT 93.3000 165.4000 95.4000 165.7000 ;
	    RECT 91.8000 164.9000 93.0000 165.2000 ;
	    RECT 91.5000 164.5000 91.9000 164.6000 ;
	    RECT 90.8000 164.2000 91.9000 164.5000 ;
	    RECT 92.7000 164.4000 93.0000 164.9000 ;
	    RECT 92.7000 164.0000 93.4000 164.4000 ;
	    RECT 89.5000 163.7000 89.9000 163.8000 ;
	    RECT 90.9000 163.7000 91.3000 163.8000 ;
	    RECT 87.8000 163.1000 88.2000 163.5000 ;
	    RECT 89.5000 163.4000 91.3000 163.7000 ;
	    RECT 90.6000 163.1000 90.9000 163.4000 ;
	    RECT 92.6000 163.1000 93.0000 163.5000 ;
	    RECT 87.8000 162.8000 88.8000 163.1000 ;
	    RECT 88.4000 161.1000 88.8000 162.8000 ;
	    RECT 90.6000 161.1000 91.0000 163.1000 ;
	    RECT 92.7000 161.1000 93.3000 163.1000 ;
	    RECT 95.0000 161.1000 95.4000 165.4000 ;
	    RECT 96.6000 161.1000 97.0000 167.8000 ;
	    RECT 98.3000 167.2000 98.6000 168.9000 ;
	    RECT 101.1000 167.9000 101.9000 169.9000 ;
	    RECT 98.2000 167.1000 98.6000 167.2000 ;
	    RECT 97.4000 166.8000 98.6000 167.1000 ;
	    RECT 100.6000 166.8000 101.0000 167.2000 ;
	    RECT 97.4000 166.2000 97.7000 166.8000 ;
	    RECT 97.4000 165.8000 97.8000 166.2000 ;
	    RECT 98.3000 165.1000 98.6000 166.8000 ;
	    RECT 100.7000 166.6000 101.0000 166.8000 ;
	    RECT 100.7000 166.2000 101.1000 166.6000 ;
	    RECT 101.4000 166.2000 101.7000 167.9000 ;
	    RECT 102.2000 166.4000 102.6000 167.2000 ;
	    RECT 99.0000 165.4000 99.4000 166.2000 ;
	    RECT 99.8000 165.4000 100.2000 166.2000 ;
	    RECT 101.4000 165.8000 101.8000 166.2000 ;
	    RECT 103.0000 166.1000 103.4000 166.2000 ;
	    RECT 103.8000 166.1000 104.2000 169.9000 ;
	    RECT 104.6000 168.1000 105.0000 168.6000 ;
	    RECT 106.2000 168.1000 106.6000 168.2000 ;
	    RECT 104.6000 167.8000 106.6000 168.1000 ;
	    RECT 107.0000 167.5000 107.4000 169.9000 ;
	    RECT 109.2000 169.2000 109.6000 169.9000 ;
	    RECT 108.6000 168.9000 109.6000 169.2000 ;
	    RECT 111.4000 168.9000 111.8000 169.9000 ;
	    RECT 113.5000 169.2000 114.1000 169.9000 ;
	    RECT 113.4000 168.9000 114.1000 169.2000 ;
	    RECT 108.6000 168.5000 109.0000 168.9000 ;
	    RECT 111.4000 168.6000 111.7000 168.9000 ;
	    RECT 109.4000 168.2000 109.8000 168.6000 ;
	    RECT 110.3000 168.3000 111.7000 168.6000 ;
	    RECT 113.4000 168.5000 113.8000 168.9000 ;
	    RECT 110.3000 168.2000 110.7000 168.3000 ;
	    RECT 107.4000 167.1000 108.2000 167.2000 ;
	    RECT 109.5000 167.1000 109.8000 168.2000 ;
	    RECT 114.3000 167.7000 114.7000 167.8000 ;
	    RECT 115.8000 167.7000 116.2000 169.9000 ;
	    RECT 116.6000 167.8000 117.0000 168.6000 ;
	    RECT 114.3000 167.4000 116.2000 167.7000 ;
	    RECT 112.3000 167.1000 112.7000 167.2000 ;
	    RECT 107.4000 166.8000 112.9000 167.1000 ;
	    RECT 108.9000 166.7000 109.3000 166.8000 ;
	    RECT 102.6000 165.8000 104.2000 166.1000 ;
	    RECT 108.1000 166.2000 108.5000 166.3000 ;
	    RECT 109.4000 166.2000 109.8000 166.3000 ;
	    RECT 108.1000 165.9000 110.6000 166.2000 ;
	    RECT 110.2000 165.8000 110.6000 165.9000 ;
	    RECT 101.4000 165.7000 101.7000 165.8000 ;
	    RECT 100.7000 165.4000 101.7000 165.7000 ;
	    RECT 102.6000 165.6000 103.0000 165.8000 ;
	    RECT 100.7000 165.1000 101.0000 165.4000 ;
	    RECT 98.2000 164.7000 99.1000 165.1000 ;
	    RECT 98.7000 161.1000 99.1000 164.7000 ;
	    RECT 99.8000 161.4000 100.2000 165.1000 ;
	    RECT 100.6000 161.7000 101.0000 165.1000 ;
	    RECT 101.4000 164.8000 103.4000 165.1000 ;
	    RECT 101.4000 161.4000 101.8000 164.8000 ;
	    RECT 99.8000 161.1000 101.8000 161.4000 ;
	    RECT 103.0000 161.1000 103.4000 164.8000 ;
	    RECT 103.8000 161.1000 104.2000 165.8000 ;
	    RECT 107.0000 165.5000 109.8000 165.6000 ;
	    RECT 107.0000 165.4000 109.9000 165.5000 ;
	    RECT 107.0000 165.3000 111.9000 165.4000 ;
	    RECT 107.0000 161.1000 107.4000 165.3000 ;
	    RECT 109.5000 165.1000 111.9000 165.3000 ;
	    RECT 108.6000 164.5000 111.3000 164.8000 ;
	    RECT 108.6000 164.4000 109.0000 164.5000 ;
	    RECT 110.9000 164.4000 111.3000 164.5000 ;
	    RECT 111.6000 164.5000 111.9000 165.1000 ;
	    RECT 112.6000 165.2000 112.9000 166.8000 ;
	    RECT 113.4000 166.4000 113.8000 166.5000 ;
	    RECT 113.4000 166.1000 115.3000 166.4000 ;
	    RECT 114.9000 166.0000 115.3000 166.1000 ;
	    RECT 114.1000 165.7000 114.5000 165.8000 ;
	    RECT 115.8000 165.7000 116.2000 167.4000 ;
	    RECT 114.1000 165.4000 116.2000 165.7000 ;
	    RECT 112.6000 164.9000 113.8000 165.2000 ;
	    RECT 112.3000 164.5000 112.7000 164.6000 ;
	    RECT 111.6000 164.2000 112.7000 164.5000 ;
	    RECT 113.5000 164.4000 113.8000 164.9000 ;
	    RECT 113.5000 164.0000 114.2000 164.4000 ;
	    RECT 110.3000 163.7000 110.7000 163.8000 ;
	    RECT 111.7000 163.7000 112.1000 163.8000 ;
	    RECT 108.6000 163.1000 109.0000 163.5000 ;
	    RECT 110.3000 163.4000 112.1000 163.7000 ;
	    RECT 111.4000 163.1000 111.7000 163.4000 ;
	    RECT 113.4000 163.1000 113.8000 163.5000 ;
	    RECT 108.6000 162.8000 109.6000 163.1000 ;
	    RECT 109.2000 161.1000 109.6000 162.8000 ;
	    RECT 111.4000 161.1000 111.8000 163.1000 ;
	    RECT 113.5000 161.1000 114.1000 163.1000 ;
	    RECT 115.8000 161.1000 116.2000 165.4000 ;
	    RECT 117.4000 166.1000 117.8000 169.9000 ;
	    RECT 119.8000 167.9000 120.2000 169.9000 ;
	    RECT 120.5000 168.2000 120.9000 168.6000 ;
	    RECT 119.0000 166.4000 119.4000 167.2000 ;
	    RECT 118.2000 166.1000 118.6000 166.2000 ;
	    RECT 119.8000 166.1000 120.1000 167.9000 ;
	    RECT 120.6000 167.8000 121.0000 168.2000 ;
	    RECT 121.4000 167.7000 121.8000 169.9000 ;
	    RECT 123.5000 169.2000 124.1000 169.9000 ;
	    RECT 123.5000 168.9000 124.2000 169.2000 ;
	    RECT 125.8000 168.9000 126.2000 169.9000 ;
	    RECT 128.0000 169.2000 128.4000 169.9000 ;
	    RECT 128.0000 168.9000 129.0000 169.2000 ;
	    RECT 123.8000 168.5000 124.2000 168.9000 ;
	    RECT 125.9000 168.6000 126.2000 168.9000 ;
	    RECT 125.9000 168.3000 127.3000 168.6000 ;
	    RECT 126.9000 168.2000 127.3000 168.3000 ;
	    RECT 127.8000 168.2000 128.2000 168.6000 ;
	    RECT 128.6000 168.5000 129.0000 168.9000 ;
	    RECT 122.9000 167.7000 123.3000 167.8000 ;
	    RECT 121.4000 167.4000 123.3000 167.7000 ;
	    RECT 120.6000 166.1000 121.0000 166.2000 ;
	    RECT 117.4000 165.8000 119.0000 166.1000 ;
	    RECT 119.8000 165.8000 121.0000 166.1000 ;
	    RECT 117.4000 161.1000 117.8000 165.8000 ;
	    RECT 118.6000 165.6000 119.0000 165.8000 ;
	    RECT 120.6000 165.1000 120.9000 165.8000 ;
	    RECT 121.4000 165.7000 121.8000 167.4000 ;
	    RECT 124.9000 167.1000 125.3000 167.2000 ;
	    RECT 127.8000 167.1000 128.1000 168.2000 ;
	    RECT 130.2000 167.5000 130.6000 169.9000 ;
	    RECT 131.0000 167.8000 131.4000 168.6000 ;
	    RECT 131.8000 168.1000 132.2000 169.9000 ;
	    RECT 133.4000 168.9000 133.8000 169.9000 ;
	    RECT 132.6000 168.1000 133.0000 168.6000 ;
	    RECT 131.8000 167.8000 133.0000 168.1000 ;
	    RECT 129.4000 167.1000 130.2000 167.2000 ;
	    RECT 124.7000 166.8000 130.2000 167.1000 ;
	    RECT 123.8000 166.4000 124.2000 166.5000 ;
	    RECT 122.3000 166.1000 124.2000 166.4000 ;
	    RECT 122.3000 166.0000 122.7000 166.1000 ;
	    RECT 123.1000 165.7000 123.5000 165.8000 ;
	    RECT 121.4000 165.4000 123.5000 165.7000 ;
	    RECT 118.2000 164.8000 120.2000 165.1000 ;
	    RECT 118.2000 161.1000 118.6000 164.8000 ;
	    RECT 119.8000 161.1000 120.2000 164.8000 ;
	    RECT 120.6000 161.1000 121.0000 165.1000 ;
	    RECT 121.4000 161.1000 121.8000 165.4000 ;
	    RECT 124.7000 165.2000 125.0000 166.8000 ;
	    RECT 128.3000 166.7000 128.7000 166.8000 ;
	    RECT 127.8000 166.2000 128.2000 166.3000 ;
	    RECT 129.1000 166.2000 129.5000 166.3000 ;
	    RECT 127.0000 165.9000 129.5000 166.2000 ;
	    RECT 127.0000 165.8000 127.4000 165.9000 ;
	    RECT 127.8000 165.5000 130.6000 165.6000 ;
	    RECT 127.7000 165.4000 130.6000 165.5000 ;
	    RECT 123.8000 164.9000 125.0000 165.2000 ;
	    RECT 125.7000 165.3000 130.6000 165.4000 ;
	    RECT 125.7000 165.1000 128.1000 165.3000 ;
	    RECT 123.8000 164.4000 124.1000 164.9000 ;
	    RECT 123.4000 164.0000 124.1000 164.4000 ;
	    RECT 124.9000 164.5000 125.3000 164.6000 ;
	    RECT 125.7000 164.5000 126.0000 165.1000 ;
	    RECT 124.9000 164.2000 126.0000 164.5000 ;
	    RECT 126.3000 164.5000 129.0000 164.8000 ;
	    RECT 126.3000 164.4000 126.7000 164.5000 ;
	    RECT 128.6000 164.4000 129.0000 164.5000 ;
	    RECT 125.5000 163.7000 125.9000 163.8000 ;
	    RECT 126.9000 163.7000 127.3000 163.8000 ;
	    RECT 123.8000 163.1000 124.2000 163.5000 ;
	    RECT 125.5000 163.4000 127.3000 163.7000 ;
	    RECT 125.9000 163.1000 126.2000 163.4000 ;
	    RECT 128.6000 163.1000 129.0000 163.5000 ;
	    RECT 123.5000 161.1000 124.1000 163.1000 ;
	    RECT 125.8000 161.1000 126.2000 163.1000 ;
	    RECT 128.0000 162.8000 129.0000 163.1000 ;
	    RECT 128.0000 161.1000 128.4000 162.8000 ;
	    RECT 130.2000 161.1000 130.6000 165.3000 ;
	    RECT 131.8000 161.1000 132.2000 167.8000 ;
	    RECT 133.5000 167.2000 133.8000 168.9000 ;
	    RECT 135.1000 168.2000 135.5000 168.6000 ;
	    RECT 135.0000 167.8000 135.4000 168.2000 ;
	    RECT 135.8000 167.9000 136.2000 169.9000 ;
	    RECT 132.6000 166.8000 133.0000 167.2000 ;
	    RECT 133.4000 166.8000 133.8000 167.2000 ;
	    RECT 132.6000 166.1000 132.9000 166.8000 ;
	    RECT 133.5000 166.1000 133.8000 166.8000 ;
	    RECT 132.6000 165.8000 133.8000 166.1000 ;
	    RECT 133.5000 165.1000 133.8000 165.8000 ;
	    RECT 134.2000 165.4000 134.6000 166.2000 ;
	    RECT 135.0000 166.1000 135.4000 166.2000 ;
	    RECT 135.9000 166.1000 136.2000 167.9000 ;
	    RECT 136.6000 166.4000 137.0000 167.2000 ;
	    RECT 137.4000 166.1000 137.8000 166.2000 ;
	    RECT 138.2000 166.1000 138.6000 169.9000 ;
	    RECT 140.6000 168.9000 141.0000 169.9000 ;
	    RECT 139.0000 168.1000 139.4000 168.6000 ;
	    RECT 139.8000 168.1000 140.2000 168.2000 ;
	    RECT 139.0000 167.8000 140.2000 168.1000 ;
	    RECT 140.6000 167.2000 140.9000 168.9000 ;
	    RECT 141.4000 168.1000 141.8000 168.6000 ;
	    RECT 142.2000 168.1000 142.6000 169.9000 ;
	    RECT 141.4000 167.8000 142.6000 168.1000 ;
	    RECT 143.0000 168.1000 143.4000 168.6000 ;
	    RECT 143.8000 168.1000 144.2000 169.9000 ;
	    RECT 145.9000 169.2000 146.5000 169.9000 ;
	    RECT 145.9000 168.9000 146.6000 169.2000 ;
	    RECT 148.2000 168.9000 148.6000 169.9000 ;
	    RECT 150.4000 169.2000 150.8000 169.9000 ;
	    RECT 150.4000 168.9000 151.4000 169.2000 ;
	    RECT 146.2000 168.5000 146.6000 168.9000 ;
	    RECT 148.3000 168.6000 148.6000 168.9000 ;
	    RECT 148.3000 168.3000 149.7000 168.6000 ;
	    RECT 149.3000 168.2000 149.7000 168.3000 ;
	    RECT 150.2000 168.2000 150.6000 168.6000 ;
	    RECT 151.0000 168.5000 151.4000 168.9000 ;
	    RECT 143.0000 167.8000 144.2000 168.1000 ;
	    RECT 140.6000 166.8000 141.0000 167.2000 ;
	    RECT 141.4000 166.8000 141.8000 167.2000 ;
	    RECT 135.0000 165.8000 136.2000 166.1000 ;
	    RECT 137.0000 165.8000 138.6000 166.1000 ;
	    RECT 135.1000 165.1000 135.4000 165.8000 ;
	    RECT 137.0000 165.6000 137.4000 165.8000 ;
	    RECT 133.4000 164.7000 134.3000 165.1000 ;
	    RECT 133.9000 161.1000 134.3000 164.7000 ;
	    RECT 135.0000 161.1000 135.4000 165.1000 ;
	    RECT 135.8000 164.8000 137.8000 165.1000 ;
	    RECT 135.8000 161.1000 136.2000 164.8000 ;
	    RECT 137.4000 161.1000 137.8000 164.8000 ;
	    RECT 138.2000 161.1000 138.6000 165.8000 ;
	    RECT 139.8000 165.4000 140.2000 166.2000 ;
	    RECT 140.6000 166.1000 140.9000 166.8000 ;
	    RECT 141.4000 166.1000 141.7000 166.8000 ;
	    RECT 140.6000 165.8000 141.7000 166.1000 ;
	    RECT 140.6000 165.1000 140.9000 165.8000 ;
	    RECT 140.1000 164.7000 141.0000 165.1000 ;
	    RECT 140.1000 161.1000 140.5000 164.7000 ;
	    RECT 142.2000 161.1000 142.6000 167.8000 ;
	    RECT 143.8000 167.7000 144.2000 167.8000 ;
	    RECT 145.3000 167.7000 145.7000 167.8000 ;
	    RECT 143.8000 167.4000 145.7000 167.7000 ;
	    RECT 143.8000 165.7000 144.2000 167.4000 ;
	    RECT 144.6000 166.8000 145.0000 167.4000 ;
	    RECT 147.3000 167.1000 147.7000 167.2000 ;
	    RECT 150.2000 167.1000 150.5000 168.2000 ;
	    RECT 152.6000 167.5000 153.0000 169.9000 ;
	    RECT 153.4000 167.8000 153.8000 168.6000 ;
	    RECT 151.8000 167.1000 152.6000 167.2000 ;
	    RECT 147.1000 166.8000 153.7000 167.1000 ;
	    RECT 146.2000 166.4000 146.6000 166.5000 ;
	    RECT 144.7000 166.1000 146.6000 166.4000 ;
	    RECT 147.1000 166.2000 147.4000 166.8000 ;
	    RECT 150.7000 166.7000 151.1000 166.8000 ;
	    RECT 151.5000 166.2000 151.9000 166.3000 ;
	    RECT 144.7000 166.0000 145.1000 166.1000 ;
	    RECT 147.0000 165.8000 147.4000 166.2000 ;
	    RECT 148.6000 166.1000 149.0000 166.2000 ;
	    RECT 149.4000 166.1000 151.9000 166.2000 ;
	    RECT 148.6000 165.9000 151.9000 166.1000 ;
	    RECT 153.4000 166.2000 153.7000 166.8000 ;
	    RECT 148.6000 165.8000 149.8000 165.9000 ;
	    RECT 153.4000 165.8000 153.8000 166.2000 ;
	    RECT 145.5000 165.7000 145.9000 165.8000 ;
	    RECT 143.8000 165.4000 145.9000 165.7000 ;
	    RECT 143.8000 161.1000 144.2000 165.4000 ;
	    RECT 147.1000 165.2000 147.4000 165.8000 ;
	    RECT 150.2000 165.5000 153.0000 165.6000 ;
	    RECT 150.1000 165.4000 153.0000 165.5000 ;
	    RECT 146.2000 164.9000 147.4000 165.2000 ;
	    RECT 148.1000 165.3000 153.0000 165.4000 ;
	    RECT 148.1000 165.1000 150.5000 165.3000 ;
	    RECT 146.2000 164.4000 146.5000 164.9000 ;
	    RECT 145.8000 164.0000 146.5000 164.4000 ;
	    RECT 147.3000 164.5000 147.7000 164.6000 ;
	    RECT 148.1000 164.5000 148.4000 165.1000 ;
	    RECT 147.3000 164.2000 148.4000 164.5000 ;
	    RECT 148.7000 164.5000 151.4000 164.8000 ;
	    RECT 148.7000 164.4000 149.1000 164.5000 ;
	    RECT 151.0000 164.4000 151.4000 164.5000 ;
	    RECT 147.9000 163.7000 148.3000 163.8000 ;
	    RECT 149.3000 163.7000 149.7000 163.8000 ;
	    RECT 146.2000 163.1000 146.6000 163.5000 ;
	    RECT 147.9000 163.4000 149.7000 163.7000 ;
	    RECT 148.3000 163.1000 148.6000 163.4000 ;
	    RECT 151.0000 163.1000 151.4000 163.5000 ;
	    RECT 145.9000 161.1000 146.5000 163.1000 ;
	    RECT 148.2000 161.1000 148.6000 163.1000 ;
	    RECT 150.4000 162.8000 151.4000 163.1000 ;
	    RECT 150.4000 161.1000 150.8000 162.8000 ;
	    RECT 152.6000 161.1000 153.0000 165.3000 ;
	    RECT 154.2000 161.1000 154.6000 169.9000 ;
	    RECT 155.0000 167.7000 155.4000 169.9000 ;
	    RECT 157.1000 169.2000 157.7000 169.9000 ;
	    RECT 157.1000 168.9000 157.8000 169.2000 ;
	    RECT 159.4000 168.9000 159.8000 169.9000 ;
	    RECT 161.6000 169.2000 162.0000 169.9000 ;
	    RECT 161.6000 168.9000 162.6000 169.2000 ;
	    RECT 157.4000 168.5000 157.8000 168.9000 ;
	    RECT 159.5000 168.6000 159.8000 168.9000 ;
	    RECT 159.5000 168.3000 160.9000 168.6000 ;
	    RECT 160.5000 168.2000 160.9000 168.3000 ;
	    RECT 161.4000 168.2000 161.8000 168.6000 ;
	    RECT 162.2000 168.5000 162.6000 168.9000 ;
	    RECT 156.5000 167.7000 156.9000 167.8000 ;
	    RECT 155.0000 167.4000 156.9000 167.7000 ;
	    RECT 155.0000 165.7000 155.4000 167.4000 ;
	    RECT 158.5000 167.1000 158.9000 167.2000 ;
	    RECT 161.4000 167.1000 161.7000 168.2000 ;
	    RECT 163.8000 167.5000 164.2000 169.9000 ;
	    RECT 167.0000 168.8000 167.4000 169.9000 ;
	    RECT 166.2000 167.8000 166.6000 168.6000 ;
	    RECT 167.1000 167.2000 167.4000 168.8000 ;
	    RECT 163.0000 167.1000 163.8000 167.2000 ;
	    RECT 158.3000 166.8000 163.8000 167.1000 ;
	    RECT 167.0000 166.8000 167.4000 167.2000 ;
	    RECT 157.4000 166.4000 157.8000 166.5000 ;
	    RECT 155.9000 166.1000 157.8000 166.4000 ;
	    RECT 158.3000 166.2000 158.6000 166.8000 ;
	    RECT 161.9000 166.7000 162.3000 166.8000 ;
	    RECT 162.7000 166.2000 163.1000 166.3000 ;
	    RECT 155.9000 166.0000 156.3000 166.1000 ;
	    RECT 158.2000 165.8000 158.6000 166.2000 ;
	    RECT 160.6000 165.9000 163.1000 166.2000 ;
	    RECT 160.6000 165.8000 161.0000 165.9000 ;
	    RECT 156.7000 165.7000 157.1000 165.8000 ;
	    RECT 155.0000 165.4000 157.1000 165.7000 ;
	    RECT 155.0000 161.1000 155.4000 165.4000 ;
	    RECT 158.3000 165.2000 158.6000 165.8000 ;
	    RECT 161.4000 165.5000 164.2000 165.6000 ;
	    RECT 161.3000 165.4000 164.2000 165.5000 ;
	    RECT 157.4000 164.9000 158.6000 165.2000 ;
	    RECT 159.3000 165.3000 164.2000 165.4000 ;
	    RECT 159.3000 165.1000 161.7000 165.3000 ;
	    RECT 157.4000 164.4000 157.7000 164.9000 ;
	    RECT 157.0000 164.0000 157.7000 164.4000 ;
	    RECT 158.5000 164.5000 158.9000 164.6000 ;
	    RECT 159.3000 164.5000 159.6000 165.1000 ;
	    RECT 158.5000 164.2000 159.6000 164.5000 ;
	    RECT 159.9000 164.5000 162.6000 164.8000 ;
	    RECT 159.9000 164.4000 160.3000 164.5000 ;
	    RECT 162.2000 164.4000 162.6000 164.5000 ;
	    RECT 159.1000 163.7000 159.5000 163.8000 ;
	    RECT 160.5000 163.7000 160.9000 163.8000 ;
	    RECT 157.4000 163.1000 157.8000 163.5000 ;
	    RECT 159.1000 163.4000 160.9000 163.7000 ;
	    RECT 159.5000 163.1000 159.8000 163.4000 ;
	    RECT 162.2000 163.1000 162.6000 163.5000 ;
	    RECT 157.1000 161.1000 157.7000 163.1000 ;
	    RECT 159.4000 161.1000 159.8000 163.1000 ;
	    RECT 161.6000 162.8000 162.6000 163.1000 ;
	    RECT 161.6000 161.1000 162.0000 162.8000 ;
	    RECT 163.8000 161.1000 164.2000 165.3000 ;
	    RECT 167.1000 165.1000 167.4000 166.8000 ;
	    RECT 169.4000 168.9000 169.8000 169.9000 ;
	    RECT 169.4000 167.2000 169.7000 168.9000 ;
	    RECT 170.2000 168.1000 170.6000 168.6000 ;
	    RECT 171.0000 168.1000 171.4000 169.9000 ;
	    RECT 170.2000 167.8000 171.4000 168.1000 ;
	    RECT 171.8000 167.8000 172.2000 168.6000 ;
	    RECT 169.4000 166.8000 169.8000 167.2000 ;
	    RECT 170.2000 166.8000 170.6000 167.2000 ;
	    RECT 167.8000 166.1000 168.2000 166.2000 ;
	    RECT 168.6000 166.1000 169.0000 166.2000 ;
	    RECT 167.8000 165.8000 169.0000 166.1000 ;
	    RECT 167.8000 165.4000 168.2000 165.8000 ;
	    RECT 168.6000 165.4000 169.0000 165.8000 ;
	    RECT 169.4000 166.1000 169.7000 166.8000 ;
	    RECT 170.2000 166.1000 170.5000 166.8000 ;
	    RECT 169.4000 165.8000 170.5000 166.1000 ;
	    RECT 169.4000 165.1000 169.7000 165.8000 ;
	    RECT 167.0000 164.7000 167.9000 165.1000 ;
	    RECT 167.5000 161.1000 167.9000 164.7000 ;
	    RECT 168.9000 164.7000 169.8000 165.1000 ;
	    RECT 168.9000 161.1000 169.3000 164.7000 ;
	    RECT 171.0000 161.1000 171.4000 167.8000 ;
	    RECT 172.6000 167.5000 173.0000 169.9000 ;
	    RECT 174.8000 169.2000 175.2000 169.9000 ;
	    RECT 174.2000 168.9000 175.2000 169.2000 ;
	    RECT 177.0000 168.9000 177.4000 169.9000 ;
	    RECT 179.1000 169.2000 179.7000 169.9000 ;
	    RECT 179.0000 168.9000 179.7000 169.2000 ;
	    RECT 174.2000 168.5000 174.6000 168.9000 ;
	    RECT 177.0000 168.6000 177.3000 168.9000 ;
	    RECT 175.0000 168.2000 175.4000 168.6000 ;
	    RECT 175.9000 168.3000 177.3000 168.6000 ;
	    RECT 179.0000 168.5000 179.4000 168.9000 ;
	    RECT 175.9000 168.2000 176.3000 168.3000 ;
	    RECT 173.0000 167.1000 173.8000 167.2000 ;
	    RECT 175.1000 167.1000 175.4000 168.2000 ;
	    RECT 179.9000 167.7000 180.3000 167.8000 ;
	    RECT 181.4000 167.7000 181.8000 169.9000 ;
	    RECT 179.9000 167.4000 181.8000 167.7000 ;
	    RECT 177.9000 167.1000 178.3000 167.2000 ;
	    RECT 173.0000 166.8000 178.5000 167.1000 ;
	    RECT 174.5000 166.7000 174.9000 166.8000 ;
	    RECT 173.7000 166.2000 174.1000 166.3000 ;
	    RECT 175.0000 166.2000 175.4000 166.3000 ;
	    RECT 173.7000 165.9000 176.2000 166.2000 ;
	    RECT 175.8000 165.8000 176.2000 165.9000 ;
	    RECT 172.6000 165.5000 175.4000 165.6000 ;
	    RECT 172.6000 165.4000 175.5000 165.5000 ;
	    RECT 172.6000 165.3000 177.5000 165.4000 ;
	    RECT 172.6000 161.1000 173.0000 165.3000 ;
	    RECT 175.1000 165.1000 177.5000 165.3000 ;
	    RECT 174.2000 164.5000 176.9000 164.8000 ;
	    RECT 174.2000 164.4000 174.6000 164.5000 ;
	    RECT 176.5000 164.4000 176.9000 164.5000 ;
	    RECT 177.2000 164.5000 177.5000 165.1000 ;
	    RECT 178.2000 165.2000 178.5000 166.8000 ;
	    RECT 179.0000 166.4000 179.4000 166.5000 ;
	    RECT 179.0000 166.1000 180.9000 166.4000 ;
	    RECT 180.5000 166.0000 180.9000 166.1000 ;
	    RECT 179.7000 165.7000 180.1000 165.8000 ;
	    RECT 181.4000 165.7000 181.8000 167.4000 ;
	    RECT 183.0000 168.9000 183.4000 169.9000 ;
	    RECT 183.0000 167.2000 183.3000 168.9000 ;
	    RECT 183.8000 168.1000 184.2000 168.6000 ;
	    RECT 184.6000 168.1000 185.0000 169.9000 ;
	    RECT 183.8000 167.8000 185.0000 168.1000 ;
	    RECT 185.4000 168.1000 185.8000 168.6000 ;
	    RECT 186.2000 168.1000 186.6000 169.9000 ;
	    RECT 188.3000 169.2000 188.9000 169.9000 ;
	    RECT 188.3000 168.9000 189.0000 169.2000 ;
	    RECT 190.6000 168.9000 191.0000 169.9000 ;
	    RECT 192.8000 169.2000 193.2000 169.9000 ;
	    RECT 192.8000 168.9000 193.8000 169.2000 ;
	    RECT 188.6000 168.5000 189.0000 168.9000 ;
	    RECT 190.7000 168.6000 191.0000 168.9000 ;
	    RECT 190.7000 168.3000 192.1000 168.6000 ;
	    RECT 191.7000 168.2000 192.1000 168.3000 ;
	    RECT 192.6000 168.2000 193.0000 168.6000 ;
	    RECT 193.4000 168.5000 193.8000 168.9000 ;
	    RECT 185.4000 167.8000 186.6000 168.1000 ;
	    RECT 183.0000 166.8000 183.4000 167.2000 ;
	    RECT 183.8000 166.8000 184.2000 167.2000 ;
	    RECT 179.7000 165.4000 181.8000 165.7000 ;
	    RECT 182.2000 165.4000 182.6000 166.2000 ;
	    RECT 183.0000 166.1000 183.3000 166.8000 ;
	    RECT 183.8000 166.1000 184.1000 166.8000 ;
	    RECT 183.0000 165.8000 184.1000 166.1000 ;
	    RECT 178.2000 164.9000 179.4000 165.2000 ;
	    RECT 177.9000 164.5000 178.3000 164.6000 ;
	    RECT 177.2000 164.2000 178.3000 164.5000 ;
	    RECT 179.1000 164.4000 179.4000 164.9000 ;
	    RECT 179.1000 164.0000 179.8000 164.4000 ;
	    RECT 175.9000 163.7000 176.3000 163.8000 ;
	    RECT 177.3000 163.7000 177.7000 163.8000 ;
	    RECT 174.2000 163.1000 174.6000 163.5000 ;
	    RECT 175.9000 163.4000 177.7000 163.7000 ;
	    RECT 177.0000 163.1000 177.3000 163.4000 ;
	    RECT 179.0000 163.1000 179.4000 163.5000 ;
	    RECT 174.2000 162.8000 175.2000 163.1000 ;
	    RECT 174.8000 161.1000 175.2000 162.8000 ;
	    RECT 177.0000 161.1000 177.4000 163.1000 ;
	    RECT 179.1000 161.1000 179.7000 163.1000 ;
	    RECT 181.4000 161.1000 181.8000 165.4000 ;
	    RECT 183.0000 165.1000 183.3000 165.8000 ;
	    RECT 182.5000 164.7000 183.4000 165.1000 ;
	    RECT 182.5000 161.1000 182.9000 164.7000 ;
	    RECT 184.6000 161.1000 185.0000 167.8000 ;
	    RECT 186.2000 167.7000 186.6000 167.8000 ;
	    RECT 187.7000 167.7000 188.1000 167.8000 ;
	    RECT 186.2000 167.4000 188.1000 167.7000 ;
	    RECT 186.2000 165.7000 186.6000 167.4000 ;
	    RECT 189.7000 167.1000 190.1000 167.2000 ;
	    RECT 191.0000 167.1000 191.4000 167.2000 ;
	    RECT 192.6000 167.1000 192.9000 168.2000 ;
	    RECT 195.0000 167.5000 195.4000 169.9000 ;
	    RECT 195.8000 167.5000 196.2000 169.9000 ;
	    RECT 198.0000 169.2000 198.4000 169.9000 ;
	    RECT 197.4000 168.9000 198.4000 169.2000 ;
	    RECT 200.2000 168.9000 200.6000 169.9000 ;
	    RECT 202.3000 169.2000 202.9000 169.9000 ;
	    RECT 202.2000 168.9000 202.9000 169.2000 ;
	    RECT 197.4000 168.5000 197.8000 168.9000 ;
	    RECT 200.2000 168.6000 200.5000 168.9000 ;
	    RECT 198.2000 168.2000 198.6000 168.6000 ;
	    RECT 199.1000 168.3000 200.5000 168.6000 ;
	    RECT 202.2000 168.5000 202.6000 168.9000 ;
	    RECT 199.1000 168.2000 199.5000 168.3000 ;
	    RECT 194.2000 167.1000 195.0000 167.2000 ;
	    RECT 196.2000 167.1000 197.0000 167.2000 ;
	    RECT 198.3000 167.1000 198.6000 168.2000 ;
	    RECT 203.1000 167.7000 203.5000 167.8000 ;
	    RECT 204.6000 167.7000 205.0000 169.9000 ;
	    RECT 205.5000 168.2000 205.9000 168.6000 ;
	    RECT 205.4000 167.8000 205.8000 168.2000 ;
	    RECT 206.2000 167.9000 206.6000 169.9000 ;
	    RECT 209.4000 168.9000 209.8000 169.9000 ;
	    RECT 203.1000 167.4000 205.0000 167.7000 ;
	    RECT 201.1000 167.1000 201.5000 167.2000 ;
	    RECT 189.5000 166.8000 201.7000 167.1000 ;
	    RECT 188.6000 166.4000 189.0000 166.5000 ;
	    RECT 187.1000 166.1000 189.0000 166.4000 ;
	    RECT 187.1000 166.0000 187.5000 166.1000 ;
	    RECT 187.9000 165.7000 188.3000 165.8000 ;
	    RECT 186.2000 165.4000 188.3000 165.7000 ;
	    RECT 186.2000 161.1000 186.6000 165.4000 ;
	    RECT 189.5000 165.2000 189.8000 166.8000 ;
	    RECT 193.1000 166.7000 193.5000 166.8000 ;
	    RECT 197.7000 166.7000 198.1000 166.8000 ;
	    RECT 193.9000 166.2000 194.3000 166.3000 ;
	    RECT 191.8000 165.9000 194.3000 166.2000 ;
	    RECT 196.9000 166.2000 197.3000 166.3000 ;
	    RECT 198.2000 166.2000 198.6000 166.3000 ;
	    RECT 196.9000 165.9000 199.4000 166.2000 ;
	    RECT 191.8000 165.8000 192.2000 165.9000 ;
	    RECT 199.0000 165.8000 199.4000 165.9000 ;
	    RECT 192.6000 165.5000 195.4000 165.6000 ;
	    RECT 192.5000 165.4000 195.4000 165.5000 ;
	    RECT 188.6000 164.9000 189.8000 165.2000 ;
	    RECT 190.5000 165.3000 195.4000 165.4000 ;
	    RECT 190.5000 165.1000 192.9000 165.3000 ;
	    RECT 188.6000 164.4000 188.9000 164.9000 ;
	    RECT 188.2000 164.0000 188.9000 164.4000 ;
	    RECT 189.7000 164.5000 190.1000 164.6000 ;
	    RECT 190.5000 164.5000 190.8000 165.1000 ;
	    RECT 189.7000 164.2000 190.8000 164.5000 ;
	    RECT 191.1000 164.5000 193.8000 164.8000 ;
	    RECT 191.1000 164.4000 191.5000 164.5000 ;
	    RECT 193.4000 164.4000 193.8000 164.5000 ;
	    RECT 190.3000 163.7000 190.7000 163.8000 ;
	    RECT 191.7000 163.7000 192.1000 163.8000 ;
	    RECT 188.6000 163.1000 189.0000 163.5000 ;
	    RECT 190.3000 163.4000 192.1000 163.7000 ;
	    RECT 190.7000 163.1000 191.0000 163.4000 ;
	    RECT 193.4000 163.1000 193.8000 163.5000 ;
	    RECT 188.3000 161.1000 188.9000 163.1000 ;
	    RECT 190.6000 161.1000 191.0000 163.1000 ;
	    RECT 192.8000 162.8000 193.8000 163.1000 ;
	    RECT 192.8000 161.1000 193.2000 162.8000 ;
	    RECT 195.0000 161.1000 195.4000 165.3000 ;
	    RECT 195.8000 165.5000 198.6000 165.6000 ;
	    RECT 195.8000 165.4000 198.7000 165.5000 ;
	    RECT 195.8000 165.3000 200.7000 165.4000 ;
	    RECT 195.8000 161.1000 196.2000 165.3000 ;
	    RECT 198.3000 165.1000 200.7000 165.3000 ;
	    RECT 197.4000 164.5000 200.1000 164.8000 ;
	    RECT 197.4000 164.4000 197.8000 164.5000 ;
	    RECT 199.7000 164.4000 200.1000 164.5000 ;
	    RECT 200.4000 164.5000 200.7000 165.1000 ;
	    RECT 201.4000 165.2000 201.7000 166.8000 ;
	    RECT 202.2000 166.4000 202.6000 166.5000 ;
	    RECT 202.2000 166.1000 204.1000 166.4000 ;
	    RECT 203.7000 166.0000 204.1000 166.1000 ;
	    RECT 202.9000 165.7000 203.3000 165.8000 ;
	    RECT 204.6000 165.7000 205.0000 167.4000 ;
	    RECT 205.4000 166.1000 205.8000 166.2000 ;
	    RECT 206.3000 166.1000 206.6000 167.9000 ;
	    RECT 208.6000 167.8000 209.0000 168.6000 ;
	    RECT 209.5000 167.2000 209.8000 168.9000 ;
	    RECT 212.9000 168.2000 213.3000 169.9000 ;
	    RECT 210.2000 168.1000 210.6000 168.2000 ;
	    RECT 212.9000 168.1000 213.8000 168.2000 ;
	    RECT 210.2000 167.8000 213.8000 168.1000 ;
	    RECT 215.0000 167.9000 215.4000 169.9000 ;
	    RECT 215.8000 168.0000 216.2000 169.9000 ;
	    RECT 217.4000 168.0000 217.8000 169.9000 ;
	    RECT 219.0000 168.9000 219.4000 169.9000 ;
	    RECT 220.9000 169.2000 221.3000 169.9000 ;
	    RECT 215.8000 167.9000 217.8000 168.0000 ;
	    RECT 207.0000 167.1000 207.4000 167.2000 ;
	    RECT 208.6000 167.1000 209.0000 167.2000 ;
	    RECT 207.0000 166.8000 209.0000 167.1000 ;
	    RECT 209.4000 166.8000 209.8000 167.2000 ;
	    RECT 207.0000 166.4000 207.4000 166.8000 ;
	    RECT 207.8000 166.1000 208.2000 166.2000 ;
	    RECT 205.4000 165.8000 206.6000 166.1000 ;
	    RECT 207.4000 165.8000 208.2000 166.1000 ;
	    RECT 202.9000 165.4000 205.0000 165.7000 ;
	    RECT 201.4000 164.9000 202.6000 165.2000 ;
	    RECT 201.1000 164.5000 201.5000 164.6000 ;
	    RECT 200.4000 164.2000 201.5000 164.5000 ;
	    RECT 202.3000 164.4000 202.6000 164.9000 ;
	    RECT 202.3000 164.2000 203.0000 164.4000 ;
	    RECT 202.3000 164.0000 203.4000 164.2000 ;
	    RECT 202.7000 163.8000 203.4000 164.0000 ;
	    RECT 199.1000 163.7000 199.5000 163.8000 ;
	    RECT 200.5000 163.7000 200.9000 163.8000 ;
	    RECT 197.4000 163.1000 197.8000 163.5000 ;
	    RECT 199.1000 163.4000 200.9000 163.7000 ;
	    RECT 200.2000 163.1000 200.5000 163.4000 ;
	    RECT 202.2000 163.1000 202.6000 163.5000 ;
	    RECT 197.4000 162.8000 198.4000 163.1000 ;
	    RECT 198.0000 161.1000 198.4000 162.8000 ;
	    RECT 200.2000 161.1000 200.6000 163.1000 ;
	    RECT 202.3000 161.1000 202.9000 163.1000 ;
	    RECT 204.6000 161.1000 205.0000 165.4000 ;
	    RECT 205.5000 165.1000 205.8000 165.8000 ;
	    RECT 207.4000 165.6000 207.8000 165.8000 ;
	    RECT 209.5000 165.1000 209.8000 166.8000 ;
	    RECT 210.2000 165.4000 210.6000 166.2000 ;
	    RECT 212.6000 165.1000 213.0000 165.2000 ;
	    RECT 205.4000 161.1000 205.8000 165.1000 ;
	    RECT 206.2000 164.8000 208.2000 165.1000 ;
	    RECT 206.2000 161.1000 206.6000 164.8000 ;
	    RECT 207.8000 161.1000 208.2000 164.8000 ;
	    RECT 209.4000 164.7000 210.3000 165.1000 ;
	    RECT 209.9000 164.1000 210.3000 164.7000 ;
	    RECT 211.8000 164.8000 213.0000 165.1000 ;
	    RECT 211.8000 164.1000 212.1000 164.8000 ;
	    RECT 212.6000 164.4000 213.0000 164.8000 ;
	    RECT 209.9000 163.8000 212.1000 164.1000 ;
	    RECT 209.9000 161.1000 210.3000 163.8000 ;
	    RECT 213.4000 161.1000 213.8000 167.8000 ;
	    RECT 214.2000 166.8000 214.6000 167.6000 ;
	    RECT 215.1000 167.2000 215.4000 167.9000 ;
	    RECT 215.9000 167.7000 217.7000 167.9000 ;
	    RECT 218.2000 167.8000 218.6000 168.6000 ;
	    RECT 217.0000 167.2000 217.4000 167.4000 ;
	    RECT 219.1000 167.2000 219.4000 168.9000 ;
	    RECT 220.6000 168.8000 221.3000 169.2000 ;
	    RECT 220.9000 168.2000 221.3000 168.8000 ;
	    RECT 224.3000 168.2000 224.7000 169.9000 ;
	    RECT 220.9000 167.9000 221.8000 168.2000 ;
	    RECT 215.0000 166.8000 216.3000 167.2000 ;
	    RECT 217.0000 166.9000 217.8000 167.2000 ;
	    RECT 217.4000 166.8000 217.8000 166.9000 ;
	    RECT 219.0000 166.8000 219.4000 167.2000 ;
	    RECT 215.0000 166.1000 215.4000 166.2000 ;
	    RECT 216.0000 166.1000 216.3000 166.8000 ;
	    RECT 215.0000 165.8000 216.3000 166.1000 ;
	    RECT 216.6000 166.1000 217.0000 166.6000 ;
	    RECT 218.2000 166.1000 218.6000 166.2000 ;
	    RECT 216.6000 165.8000 218.6000 166.1000 ;
	    RECT 215.0000 165.1000 215.4000 165.2000 ;
	    RECT 216.0000 165.1000 216.3000 165.8000 ;
	    RECT 219.1000 165.1000 219.4000 166.8000 ;
	    RECT 219.8000 165.4000 220.2000 166.2000 ;
	    RECT 215.0000 164.8000 215.7000 165.1000 ;
	    RECT 216.0000 164.8000 216.5000 165.1000 ;
	    RECT 215.4000 164.2000 215.7000 164.8000 ;
	    RECT 215.4000 163.8000 215.8000 164.2000 ;
	    RECT 216.1000 161.1000 216.5000 164.8000 ;
	    RECT 219.0000 164.7000 219.9000 165.1000 ;
	    RECT 219.5000 164.1000 219.9000 164.7000 ;
	    RECT 220.6000 164.1000 221.0000 165.2000 ;
	    RECT 219.5000 163.8000 221.0000 164.1000 ;
	    RECT 219.5000 161.1000 219.9000 163.8000 ;
	    RECT 221.4000 161.1000 221.8000 167.9000 ;
	    RECT 223.8000 168.1000 224.7000 168.2000 ;
	    RECT 225.4000 168.1000 225.8000 168.6000 ;
	    RECT 223.8000 167.8000 225.8000 168.1000 ;
	    RECT 222.2000 166.8000 222.6000 167.6000 ;
	    RECT 223.0000 166.8000 223.4000 167.6000 ;
	    RECT 223.8000 161.1000 224.2000 167.8000 ;
	    RECT 226.2000 167.1000 226.6000 169.9000 ;
	    RECT 227.8000 168.9000 228.2000 169.9000 ;
	    RECT 227.0000 167.8000 227.4000 168.6000 ;
	    RECT 227.9000 167.2000 228.2000 168.9000 ;
	    RECT 229.4000 168.0000 229.8000 169.9000 ;
	    RECT 231.0000 168.0000 231.4000 169.9000 ;
	    RECT 229.4000 167.9000 231.4000 168.0000 ;
	    RECT 231.8000 167.9000 232.2000 169.9000 ;
	    RECT 232.6000 168.0000 233.0000 169.9000 ;
	    RECT 234.2000 168.0000 234.6000 169.9000 ;
	    RECT 232.6000 167.9000 234.6000 168.0000 ;
	    RECT 235.0000 167.9000 235.4000 169.9000 ;
	    RECT 235.8000 168.0000 236.2000 169.9000 ;
	    RECT 237.4000 168.0000 237.8000 169.9000 ;
	    RECT 235.8000 167.9000 237.8000 168.0000 ;
	    RECT 238.2000 167.9000 238.6000 169.9000 ;
	    RECT 239.0000 169.6000 241.0000 169.9000 ;
	    RECT 239.0000 167.9000 239.4000 169.6000 ;
	    RECT 239.8000 167.9000 240.2000 169.3000 ;
	    RECT 240.6000 168.0000 241.0000 169.6000 ;
	    RECT 242.2000 168.0000 242.6000 169.9000 ;
	    RECT 243.3000 168.4000 243.7000 169.9000 ;
	    RECT 240.6000 167.9000 242.6000 168.0000 ;
	    RECT 243.0000 167.9000 243.7000 168.4000 ;
	    RECT 245.4000 167.9000 245.8000 169.9000 ;
	    RECT 246.2000 168.0000 246.6000 169.9000 ;
	    RECT 247.8000 168.0000 248.2000 169.9000 ;
	    RECT 246.2000 167.9000 248.2000 168.0000 ;
	    RECT 248.6000 167.9000 249.0000 169.9000 ;
	    RECT 250.2000 168.2000 250.6000 169.9000 ;
	    RECT 250.1000 167.9000 250.6000 168.2000 ;
	    RECT 229.5000 167.7000 231.3000 167.9000 ;
	    RECT 229.8000 167.2000 230.2000 167.4000 ;
	    RECT 231.8000 167.2000 232.1000 167.9000 ;
	    RECT 232.7000 167.7000 234.5000 167.9000 ;
	    RECT 233.0000 167.2000 233.4000 167.4000 ;
	    RECT 235.0000 167.2000 235.3000 167.9000 ;
	    RECT 235.9000 167.7000 237.7000 167.9000 ;
	    RECT 236.2000 167.2000 236.6000 167.4000 ;
	    RECT 238.2000 167.2000 238.5000 167.9000 ;
	    RECT 239.8000 167.2000 240.1000 167.9000 ;
	    RECT 240.7000 167.7000 242.5000 167.9000 ;
	    RECT 241.8000 167.2000 242.2000 167.4000 ;
	    RECT 226.2000 166.8000 227.3000 167.1000 ;
	    RECT 227.8000 166.8000 228.2000 167.2000 ;
	    RECT 229.4000 166.9000 230.2000 167.2000 ;
	    RECT 229.4000 166.8000 229.8000 166.9000 ;
	    RECT 230.9000 166.8000 232.2000 167.2000 ;
	    RECT 232.6000 166.9000 233.4000 167.2000 ;
	    RECT 232.6000 166.8000 233.0000 166.9000 ;
	    RECT 234.1000 166.8000 235.4000 167.2000 ;
	    RECT 235.8000 166.9000 236.6000 167.2000 ;
	    RECT 235.8000 166.8000 236.2000 166.9000 ;
	    RECT 237.3000 166.8000 238.6000 167.2000 ;
	    RECT 224.6000 164.4000 225.0000 165.2000 ;
	    RECT 226.2000 161.1000 226.6000 166.8000 ;
	    RECT 227.0000 166.2000 227.3000 166.8000 ;
	    RECT 227.9000 166.2000 228.2000 166.8000 ;
	    RECT 227.0000 165.8000 227.4000 166.2000 ;
	    RECT 227.8000 165.8000 228.2000 166.2000 ;
	    RECT 227.9000 165.1000 228.2000 165.8000 ;
	    RECT 228.6000 166.1000 229.0000 166.2000 ;
	    RECT 229.4000 166.1000 229.8000 166.2000 ;
	    RECT 228.6000 165.8000 229.8000 166.1000 ;
	    RECT 230.2000 165.8000 230.6000 166.6000 ;
	    RECT 230.9000 166.2000 231.2000 166.8000 ;
	    RECT 230.9000 165.8000 231.4000 166.2000 ;
	    RECT 233.4000 166.1000 233.8000 166.6000 ;
	    RECT 231.8000 165.8000 233.8000 166.1000 ;
	    RECT 228.6000 165.4000 229.0000 165.8000 ;
	    RECT 230.9000 165.1000 231.2000 165.8000 ;
	    RECT 231.8000 165.2000 232.1000 165.8000 ;
	    RECT 231.8000 165.1000 232.2000 165.2000 ;
	    RECT 234.1000 165.1000 234.4000 166.8000 ;
	    RECT 236.6000 165.8000 237.0000 166.6000 ;
	    RECT 237.3000 165.2000 237.6000 166.8000 ;
	    RECT 239.0000 166.4000 239.4000 167.2000 ;
	    RECT 239.8000 166.9000 241.0000 167.2000 ;
	    RECT 241.8000 166.9000 242.6000 167.2000 ;
	    RECT 240.6000 166.8000 241.0000 166.9000 ;
	    RECT 239.8000 165.8000 240.2000 166.6000 ;
	    RECT 235.0000 165.1000 235.4000 165.2000 ;
	    RECT 227.8000 164.7000 228.7000 165.1000 ;
	    RECT 228.3000 161.1000 228.7000 164.7000 ;
	    RECT 230.7000 164.8000 231.2000 165.1000 ;
	    RECT 231.5000 164.8000 232.2000 165.1000 ;
	    RECT 233.9000 164.8000 234.4000 165.1000 ;
	    RECT 234.7000 164.8000 235.4000 165.1000 ;
	    RECT 236.6000 164.8000 237.6000 165.2000 ;
	    RECT 238.2000 165.1000 238.6000 165.2000 ;
	    RECT 240.7000 165.1000 241.0000 166.8000 ;
	    RECT 242.2000 166.8000 242.6000 166.9000 ;
	    RECT 241.4000 165.8000 241.8000 166.6000 ;
	    RECT 242.2000 166.1000 242.5000 166.8000 ;
	    RECT 243.0000 166.2000 243.3000 167.9000 ;
	    RECT 245.4000 167.8000 245.7000 167.9000 ;
	    RECT 244.8000 167.6000 245.7000 167.8000 ;
	    RECT 246.3000 167.7000 248.1000 167.9000 ;
	    RECT 243.6000 167.5000 245.7000 167.6000 ;
	    RECT 243.6000 167.3000 245.1000 167.5000 ;
	    RECT 243.6000 167.2000 244.0000 167.3000 ;
	    RECT 246.6000 167.2000 247.0000 167.4000 ;
	    RECT 248.6000 167.2000 248.9000 167.9000 ;
	    RECT 250.1000 167.2000 250.4000 167.9000 ;
	    RECT 251.8000 167.6000 252.2000 169.9000 ;
	    RECT 252.6000 168.0000 253.0000 169.9000 ;
	    RECT 254.2000 168.0000 254.6000 169.9000 ;
	    RECT 252.6000 167.9000 254.6000 168.0000 ;
	    RECT 255.0000 167.9000 255.4000 169.9000 ;
	    RECT 255.9000 168.2000 256.3000 168.6000 ;
	    RECT 252.7000 167.7000 254.5000 167.9000 ;
	    RECT 250.9000 167.3000 252.2000 167.6000 ;
	    RECT 243.0000 166.1000 243.4000 166.2000 ;
	    RECT 242.2000 165.8000 243.4000 166.1000 ;
	    RECT 243.0000 165.1000 243.3000 165.8000 ;
	    RECT 243.7000 165.5000 244.0000 167.2000 ;
	    RECT 244.4000 166.9000 244.8000 167.0000 ;
	    RECT 244.4000 166.6000 244.9000 166.9000 ;
	    RECT 244.6000 166.2000 244.9000 166.6000 ;
	    RECT 245.4000 166.4000 245.8000 167.2000 ;
	    RECT 246.2000 166.9000 247.0000 167.2000 ;
	    RECT 246.2000 166.8000 246.6000 166.9000 ;
	    RECT 247.7000 166.8000 249.0000 167.2000 ;
	    RECT 250.1000 167.1000 250.6000 167.2000 ;
	    RECT 249.4000 166.8000 250.6000 167.1000 ;
	    RECT 244.6000 165.8000 245.0000 166.2000 ;
	    RECT 246.2000 166.1000 246.6000 166.2000 ;
	    RECT 247.0000 166.1000 247.4000 166.6000 ;
	    RECT 246.2000 165.8000 247.4000 166.1000 ;
	    RECT 247.7000 166.1000 248.0000 166.8000 ;
	    RECT 249.4000 166.2000 249.7000 166.8000 ;
	    RECT 248.6000 166.1000 249.0000 166.2000 ;
	    RECT 247.7000 165.8000 249.0000 166.1000 ;
	    RECT 249.4000 165.8000 249.8000 166.2000 ;
	    RECT 243.7000 165.2000 244.9000 165.5000 ;
	    RECT 237.9000 164.8000 238.6000 165.1000 ;
	    RECT 230.7000 161.1000 231.1000 164.8000 ;
	    RECT 231.5000 164.2000 231.8000 164.8000 ;
	    RECT 231.4000 163.8000 231.8000 164.2000 ;
	    RECT 233.9000 161.1000 234.3000 164.8000 ;
	    RECT 234.7000 164.2000 235.0000 164.8000 ;
	    RECT 234.6000 163.8000 235.0000 164.2000 ;
	    RECT 237.1000 161.1000 237.5000 164.8000 ;
	    RECT 237.9000 164.2000 238.2000 164.8000 ;
	    RECT 237.8000 163.8000 238.2000 164.2000 ;
	    RECT 240.3000 161.1000 241.3000 165.1000 ;
	    RECT 243.0000 161.1000 243.4000 165.1000 ;
	    RECT 244.6000 163.1000 244.9000 165.2000 ;
	    RECT 247.7000 165.1000 248.0000 165.8000 ;
	    RECT 248.6000 165.1000 249.0000 165.2000 ;
	    RECT 247.5000 164.8000 248.0000 165.1000 ;
	    RECT 248.3000 164.8000 249.0000 165.1000 ;
	    RECT 250.1000 165.1000 250.4000 166.8000 ;
	    RECT 250.9000 166.5000 251.2000 167.3000 ;
	    RECT 253.0000 167.2000 253.4000 167.4000 ;
	    RECT 255.0000 167.2000 255.3000 167.9000 ;
	    RECT 255.8000 167.8000 256.2000 168.2000 ;
	    RECT 256.6000 167.9000 257.0000 169.9000 ;
	    RECT 259.1000 168.2000 259.5000 168.6000 ;
	    RECT 252.6000 166.9000 253.4000 167.2000 ;
	    RECT 252.6000 166.8000 253.0000 166.9000 ;
	    RECT 254.1000 166.8000 255.4000 167.2000 ;
	    RECT 250.7000 166.1000 251.2000 166.5000 ;
	    RECT 250.9000 165.1000 251.2000 166.1000 ;
	    RECT 251.7000 166.2000 252.1000 166.6000 ;
	    RECT 251.7000 165.8000 252.2000 166.2000 ;
	    RECT 253.4000 165.8000 253.8000 166.6000 ;
	    RECT 254.1000 166.2000 254.4000 166.8000 ;
	    RECT 254.1000 165.8000 254.6000 166.2000 ;
	    RECT 255.8000 166.1000 256.2000 166.2000 ;
	    RECT 256.7000 166.1000 257.0000 167.9000 ;
	    RECT 259.0000 167.8000 259.4000 168.2000 ;
	    RECT 259.8000 167.9000 260.2000 169.9000 ;
	    RECT 257.4000 166.4000 257.8000 167.2000 ;
	    RECT 258.2000 166.1000 258.6000 166.2000 ;
	    RECT 259.0000 166.1000 259.4000 166.2000 ;
	    RECT 259.9000 166.1000 260.2000 167.9000 ;
	    RECT 262.2000 167.9000 262.6000 169.9000 ;
	    RECT 264.4000 169.2000 265.2000 169.9000 ;
	    RECT 263.8000 168.8000 265.2000 169.2000 ;
	    RECT 264.4000 168.1000 265.2000 168.8000 ;
	    RECT 262.2000 167.6000 263.4000 167.9000 ;
	    RECT 263.0000 167.5000 263.4000 167.6000 ;
	    RECT 263.7000 167.4000 264.1000 167.8000 ;
	    RECT 263.7000 167.2000 264.0000 167.4000 ;
	    RECT 260.6000 166.4000 261.0000 167.2000 ;
	    RECT 262.2000 166.8000 263.0000 167.2000 ;
	    RECT 263.6000 166.8000 264.0000 167.2000 ;
	    RECT 264.4000 167.1000 264.7000 168.1000 ;
	    RECT 267.0000 167.9000 267.4000 169.9000 ;
	    RECT 265.0000 167.4000 265.8000 167.8000 ;
	    RECT 266.1000 167.6000 267.4000 167.9000 ;
	    RECT 267.8000 167.6000 268.2000 169.9000 ;
	    RECT 269.4000 168.2000 269.8000 169.9000 ;
	    RECT 269.4000 167.9000 269.9000 168.2000 ;
	    RECT 266.1000 167.5000 266.5000 167.6000 ;
	    RECT 267.8000 167.3000 269.1000 167.6000 ;
	    RECT 264.4000 166.8000 264.9000 167.1000 ;
	    RECT 264.6000 166.2000 264.9000 166.8000 ;
	    RECT 267.9000 166.2000 268.3000 166.6000 ;
	    RECT 261.4000 166.1000 261.8000 166.2000 ;
	    RECT 255.8000 165.8000 257.0000 166.1000 ;
	    RECT 257.8000 165.8000 260.2000 166.1000 ;
	    RECT 261.0000 165.8000 261.8000 166.1000 ;
	    RECT 264.6000 165.8000 265.0000 166.2000 ;
	    RECT 265.9000 166.1000 266.3000 166.2000 ;
	    RECT 265.5000 165.8000 266.3000 166.1000 ;
	    RECT 267.8000 165.8000 268.3000 166.2000 ;
	    RECT 268.8000 166.5000 269.1000 167.3000 ;
	    RECT 269.6000 167.2000 269.9000 167.9000 ;
	    RECT 269.4000 166.8000 269.9000 167.2000 ;
	    RECT 268.8000 166.1000 269.3000 166.5000 ;
	    RECT 254.1000 165.1000 254.4000 165.8000 ;
	    RECT 255.0000 165.1000 255.4000 165.2000 ;
	    RECT 255.9000 165.1000 256.2000 165.8000 ;
	    RECT 257.8000 165.6000 258.2000 165.8000 ;
	    RECT 259.1000 165.1000 259.4000 165.8000 ;
	    RECT 261.0000 165.6000 261.4000 165.8000 ;
	    RECT 264.6000 165.1000 264.9000 165.8000 ;
	    RECT 265.5000 165.7000 265.9000 165.8000 ;
	    RECT 268.8000 165.1000 269.1000 166.1000 ;
	    RECT 269.6000 165.1000 269.9000 166.8000 ;
	    RECT 244.6000 161.1000 245.0000 163.1000 ;
	    RECT 247.5000 161.1000 247.9000 164.8000 ;
	    RECT 248.3000 164.2000 248.6000 164.8000 ;
	    RECT 250.1000 164.6000 250.6000 165.1000 ;
	    RECT 250.9000 164.8000 252.2000 165.1000 ;
	    RECT 248.2000 163.8000 248.6000 164.2000 ;
	    RECT 250.2000 161.1000 250.6000 164.6000 ;
	    RECT 251.8000 161.1000 252.2000 164.8000 ;
	    RECT 253.9000 164.8000 254.4000 165.1000 ;
	    RECT 254.7000 164.8000 255.4000 165.1000 ;
	    RECT 253.9000 161.1000 254.3000 164.8000 ;
	    RECT 254.7000 164.2000 255.0000 164.8000 ;
	    RECT 254.6000 163.8000 255.0000 164.2000 ;
	    RECT 255.8000 161.1000 256.2000 165.1000 ;
	    RECT 256.6000 164.8000 258.6000 165.1000 ;
	    RECT 256.6000 161.1000 257.0000 164.8000 ;
	    RECT 258.2000 161.1000 258.6000 164.8000 ;
	    RECT 259.0000 161.1000 259.4000 165.1000 ;
	    RECT 259.8000 164.8000 261.8000 165.1000 ;
	    RECT 259.8000 161.1000 260.2000 164.8000 ;
	    RECT 261.4000 161.1000 261.8000 164.8000 ;
	    RECT 262.2000 164.8000 263.4000 165.1000 ;
	    RECT 262.2000 161.1000 262.6000 164.8000 ;
	    RECT 263.0000 164.7000 263.4000 164.8000 ;
	    RECT 264.4000 161.1000 265.2000 165.1000 ;
	    RECT 266.1000 164.8000 267.4000 165.1000 ;
	    RECT 266.1000 164.7000 266.5000 164.8000 ;
	    RECT 267.0000 161.1000 267.4000 164.8000 ;
	    RECT 267.8000 164.8000 269.1000 165.1000 ;
	    RECT 267.8000 161.1000 268.2000 164.8000 ;
	    RECT 269.4000 164.6000 269.9000 165.1000 ;
	    RECT 269.4000 161.1000 269.8000 164.6000 ;
	    RECT 1.4000 154.1000 1.8000 159.9000 ;
	    RECT 2.2000 159.6000 4.2000 159.9000 ;
	    RECT 2.2000 155.9000 2.6000 159.6000 ;
	    RECT 3.0000 155.9000 3.4000 159.3000 ;
	    RECT 3.8000 156.2000 4.2000 159.6000 ;
	    RECT 5.4000 156.2000 5.8000 159.9000 ;
	    RECT 3.8000 155.9000 5.8000 156.2000 ;
	    RECT 3.1000 155.6000 3.4000 155.9000 ;
	    RECT 3.1000 155.3000 4.1000 155.6000 ;
	    RECT 3.8000 155.2000 4.1000 155.3000 ;
	    RECT 5.0000 155.2000 5.4000 155.4000 ;
	    RECT 3.8000 154.8000 4.2000 155.2000 ;
	    RECT 5.0000 155.1000 5.8000 155.2000 ;
	    RECT 6.2000 155.1000 6.6000 159.9000 ;
	    RECT 5.0000 154.9000 6.6000 155.1000 ;
	    RECT 5.4000 154.8000 6.6000 154.9000 ;
	    RECT 3.1000 154.4000 3.5000 154.8000 ;
	    RECT 3.1000 154.2000 3.4000 154.4000 ;
	    RECT 3.0000 154.1000 3.4000 154.2000 ;
	    RECT 1.4000 153.8000 3.4000 154.1000 ;
	    RECT 1.4000 151.1000 1.8000 153.8000 ;
	    RECT 3.8000 153.1000 4.1000 154.8000 ;
	    RECT 3.5000 151.1000 4.3000 153.1000 ;
	    RECT 6.2000 151.1000 6.6000 154.8000 ;
	    RECT 8.6000 156.1000 9.0000 159.9000 ;
	    RECT 9.4000 156.1000 9.8000 156.6000 ;
	    RECT 8.6000 155.8000 9.8000 156.1000 ;
	    RECT 8.6000 154.1000 9.0000 155.8000 ;
	    RECT 9.4000 154.1000 9.8000 154.2000 ;
	    RECT 8.6000 153.8000 9.8000 154.1000 ;
	    RECT 8.6000 151.1000 9.0000 153.8000 ;
	    RECT 10.2000 153.1000 10.6000 159.9000 ;
	    RECT 9.7000 152.8000 10.6000 153.1000 ;
	    RECT 12.6000 155.1000 13.0000 159.9000 ;
	    RECT 15.0000 157.9000 15.4000 159.9000 ;
	    RECT 15.1000 157.8000 15.4000 157.9000 ;
	    RECT 16.6000 157.9000 17.0000 159.9000 ;
	    RECT 16.6000 157.8000 16.9000 157.9000 ;
	    RECT 15.1000 157.5000 16.9000 157.8000 ;
	    RECT 13.4000 155.8000 13.8000 156.6000 ;
	    RECT 15.8000 156.4000 16.2000 157.2000 ;
	    RECT 16.6000 156.2000 16.9000 157.5000 ;
	    RECT 17.7000 156.3000 18.1000 159.9000 ;
	    RECT 14.2000 155.4000 14.6000 156.2000 ;
	    RECT 16.6000 155.8000 17.0000 156.2000 ;
	    RECT 17.7000 155.9000 18.6000 156.3000 ;
	    RECT 12.6000 154.8000 13.7000 155.1000 ;
	    RECT 15.0000 154.8000 15.8000 155.2000 ;
	    RECT 16.6000 155.1000 16.9000 155.8000 ;
	    RECT 17.4000 155.1000 17.8000 155.6000 ;
	    RECT 16.6000 154.8000 17.8000 155.1000 ;
	    RECT 12.6000 153.1000 13.0000 154.8000 ;
	    RECT 13.4000 154.2000 13.7000 154.8000 ;
	    RECT 16.6000 154.2000 16.9000 154.8000 ;
	    RECT 13.4000 153.8000 13.8000 154.2000 ;
	    RECT 16.1000 154.1000 16.9000 154.2000 ;
	    RECT 16.0000 153.9000 16.9000 154.1000 ;
	    RECT 18.2000 154.2000 18.5000 155.9000 ;
	    RECT 19.8000 155.6000 20.2000 159.9000 ;
	    RECT 21.9000 156.2000 22.3000 159.9000 ;
	    RECT 24.3000 156.2000 24.7000 159.9000 ;
	    RECT 25.0000 156.8000 25.4000 157.2000 ;
	    RECT 25.1000 156.2000 25.4000 156.8000 ;
	    RECT 27.5000 156.3000 27.9000 159.9000 ;
	    RECT 28.6000 157.9000 29.0000 159.9000 ;
	    RECT 21.9000 155.9000 22.6000 156.2000 ;
	    RECT 24.3000 155.9000 24.8000 156.2000 ;
	    RECT 25.1000 155.9000 25.8000 156.2000 ;
	    RECT 27.0000 155.9000 27.9000 156.3000 ;
	    RECT 28.7000 157.8000 29.0000 157.9000 ;
	    RECT 30.2000 157.9000 30.6000 159.9000 ;
	    RECT 30.2000 157.8000 30.5000 157.9000 ;
	    RECT 28.7000 157.5000 30.5000 157.8000 ;
	    RECT 28.7000 156.2000 29.0000 157.5000 ;
	    RECT 29.4000 156.4000 29.8000 157.2000 ;
	    RECT 31.8000 156.2000 32.2000 159.9000 ;
	    RECT 33.4000 159.6000 35.4000 159.9000 ;
	    RECT 33.4000 156.2000 33.8000 159.6000 ;
	    RECT 19.8000 155.4000 21.8000 155.6000 ;
	    RECT 19.8000 155.3000 21.9000 155.4000 ;
	    RECT 21.5000 155.0000 21.9000 155.3000 ;
	    RECT 22.3000 155.2000 22.6000 155.9000 ;
	    RECT 20.8000 154.2000 21.2000 154.6000 ;
	    RECT 12.6000 152.8000 13.5000 153.1000 ;
	    RECT 9.7000 152.2000 10.1000 152.8000 ;
	    RECT 9.7000 151.8000 10.6000 152.2000 ;
	    RECT 9.7000 151.1000 10.1000 151.8000 ;
	    RECT 13.1000 151.1000 13.5000 152.8000 ;
	    RECT 16.0000 151.1000 16.4000 153.9000 ;
	    RECT 18.2000 153.8000 18.6000 154.2000 ;
	    RECT 20.6000 153.8000 21.1000 154.2000 ;
	    RECT 18.2000 152.2000 18.5000 153.8000 ;
	    RECT 21.6000 153.5000 21.9000 155.0000 ;
	    RECT 22.2000 155.1000 22.6000 155.2000 ;
	    RECT 23.8000 155.1000 24.2000 155.2000 ;
	    RECT 22.2000 154.8000 24.2000 155.1000 ;
	    RECT 20.7000 153.2000 21.9000 153.5000 ;
	    RECT 19.0000 152.4000 19.4000 153.2000 ;
	    RECT 19.8000 152.4000 20.2000 153.2000 ;
	    RECT 18.2000 151.1000 18.6000 152.2000 ;
	    RECT 20.7000 152.1000 21.0000 153.2000 ;
	    RECT 22.3000 153.1000 22.6000 154.8000 ;
	    RECT 23.8000 154.4000 24.2000 154.8000 ;
	    RECT 24.5000 154.2000 24.8000 155.9000 ;
	    RECT 25.4000 155.8000 25.8000 155.9000 ;
	    RECT 27.1000 154.2000 27.4000 155.9000 ;
	    RECT 28.6000 155.8000 29.0000 156.2000 ;
	    RECT 27.8000 154.8000 28.2000 155.6000 ;
	    RECT 23.0000 154.1000 23.4000 154.2000 ;
	    RECT 23.0000 153.8000 23.8000 154.1000 ;
	    RECT 24.5000 153.8000 25.8000 154.2000 ;
	    RECT 27.0000 153.8000 27.4000 154.2000 ;
	    RECT 28.7000 154.2000 29.0000 155.8000 ;
	    RECT 31.0000 155.4000 31.4000 156.2000 ;
	    RECT 31.8000 155.9000 33.8000 156.2000 ;
	    RECT 34.2000 155.9000 34.6000 159.3000 ;
	    RECT 35.0000 155.9000 35.4000 159.6000 ;
	    RECT 35.8000 156.2000 36.2000 159.9000 ;
	    RECT 37.4000 156.2000 37.8000 159.9000 ;
	    RECT 35.8000 155.9000 37.8000 156.2000 ;
	    RECT 38.2000 155.9000 38.6000 159.9000 ;
	    RECT 39.3000 156.3000 39.7000 159.9000 ;
	    RECT 39.3000 155.9000 40.2000 156.3000 ;
	    RECT 42.7000 156.2000 43.1000 159.9000 ;
	    RECT 43.4000 156.8000 43.8000 157.2000 ;
	    RECT 43.5000 156.2000 43.8000 156.8000 ;
	    RECT 46.2000 156.2000 46.6000 159.9000 ;
	    RECT 42.7000 155.9000 43.2000 156.2000 ;
	    RECT 43.5000 155.9000 44.2000 156.2000 ;
	    RECT 34.2000 155.6000 34.5000 155.9000 ;
	    RECT 32.2000 155.2000 32.6000 155.4000 ;
	    RECT 33.5000 155.3000 34.5000 155.6000 ;
	    RECT 33.5000 155.2000 33.8000 155.3000 ;
	    RECT 29.8000 154.8000 30.6000 155.2000 ;
	    RECT 31.8000 154.9000 32.6000 155.2000 ;
	    RECT 31.8000 154.8000 32.2000 154.9000 ;
	    RECT 33.4000 154.8000 33.8000 155.2000 ;
	    RECT 35.0000 154.8000 35.4000 155.6000 ;
	    RECT 36.2000 155.2000 36.6000 155.4000 ;
	    RECT 38.2000 155.2000 38.5000 155.9000 ;
	    RECT 35.8000 154.9000 36.6000 155.2000 ;
	    RECT 37.4000 155.1000 38.6000 155.2000 ;
	    RECT 39.0000 155.1000 39.4000 155.6000 ;
	    RECT 37.4000 154.9000 39.4000 155.1000 ;
	    RECT 35.8000 154.8000 36.2000 154.9000 ;
	    RECT 28.7000 154.1000 29.5000 154.2000 ;
	    RECT 23.4000 153.6000 23.8000 153.8000 ;
	    RECT 23.1000 153.1000 24.9000 153.3000 ;
	    RECT 25.4000 153.1000 25.7000 153.8000 ;
	    RECT 20.6000 151.1000 21.0000 152.1000 ;
	    RECT 22.2000 151.1000 22.6000 153.1000 ;
	    RECT 23.0000 153.0000 25.0000 153.1000 ;
	    RECT 23.0000 151.1000 23.4000 153.0000 ;
	    RECT 24.6000 151.1000 25.0000 153.0000 ;
	    RECT 25.4000 151.1000 25.8000 153.1000 ;
	    RECT 26.2000 152.4000 26.6000 153.2000 ;
	    RECT 27.1000 152.2000 27.4000 153.8000 ;
	    RECT 27.8000 153.8000 29.6000 154.1000 ;
	    RECT 27.8000 153.2000 28.1000 153.8000 ;
	    RECT 27.8000 152.8000 28.2000 153.2000 ;
	    RECT 27.0000 151.1000 27.4000 152.2000 ;
	    RECT 29.2000 151.1000 29.6000 153.8000 ;
	    RECT 33.5000 153.1000 33.8000 154.8000 ;
	    RECT 37.4000 153.1000 37.7000 154.9000 ;
	    RECT 38.2000 154.8000 39.4000 154.9000 ;
	    RECT 39.8000 154.2000 40.1000 155.9000 ;
	    RECT 42.9000 154.2000 43.2000 155.9000 ;
	    RECT 43.8000 155.8000 44.2000 155.9000 ;
	    RECT 45.5000 155.9000 46.6000 156.2000 ;
	    RECT 45.5000 155.6000 45.8000 155.9000 ;
	    RECT 45.2000 155.2000 45.8000 155.6000 ;
	    RECT 39.0000 153.8000 39.4000 154.2000 ;
	    RECT 39.8000 153.8000 40.2000 154.2000 ;
	    RECT 40.6000 154.1000 41.0000 154.2000 ;
	    RECT 41.4000 154.1000 41.8000 154.2000 ;
	    RECT 40.6000 153.8000 42.2000 154.1000 ;
	    RECT 42.9000 153.8000 44.2000 154.2000 ;
	    RECT 33.3000 151.1000 34.1000 153.1000 ;
	    RECT 37.4000 151.1000 37.8000 153.1000 ;
	    RECT 38.2000 152.8000 38.6000 153.2000 ;
	    RECT 39.0000 153.1000 39.3000 153.8000 ;
	    RECT 39.8000 153.1000 40.1000 153.8000 ;
	    RECT 41.8000 153.6000 42.2000 153.8000 ;
	    RECT 39.0000 152.8000 40.1000 153.1000 ;
	    RECT 38.1000 152.4000 38.5000 152.8000 ;
	    RECT 39.8000 152.1000 40.1000 152.8000 ;
	    RECT 40.6000 152.4000 41.0000 153.2000 ;
	    RECT 41.5000 153.1000 43.3000 153.3000 ;
	    RECT 43.8000 153.1000 44.1000 153.8000 ;
	    RECT 45.5000 153.7000 45.8000 155.2000 ;
	    RECT 46.2000 155.1000 46.6000 155.2000 ;
	    RECT 47.0000 155.1000 47.4000 155.2000 ;
	    RECT 46.2000 154.8000 47.4000 155.1000 ;
	    RECT 46.2000 154.4000 46.6000 154.8000 ;
	    RECT 45.5000 153.4000 46.6000 153.7000 ;
	    RECT 41.4000 153.0000 43.4000 153.1000 ;
	    RECT 39.8000 151.1000 40.2000 152.1000 ;
	    RECT 41.4000 151.1000 41.8000 153.0000 ;
	    RECT 43.0000 151.1000 43.4000 153.0000 ;
	    RECT 43.8000 151.1000 44.2000 153.1000 ;
	    RECT 46.2000 151.1000 46.6000 153.4000 ;
	    RECT 47.0000 152.4000 47.4000 153.2000 ;
	    RECT 47.8000 153.1000 48.2000 159.9000 ;
	    RECT 49.9000 156.3000 50.3000 159.9000 ;
	    RECT 49.4000 155.9000 50.3000 156.3000 ;
	    RECT 49.4000 155.8000 49.8000 155.9000 ;
	    RECT 49.5000 154.2000 49.8000 155.8000 ;
	    RECT 51.0000 155.6000 51.4000 159.9000 ;
	    RECT 53.1000 157.9000 53.7000 159.9000 ;
	    RECT 55.4000 157.9000 55.8000 159.9000 ;
	    RECT 57.6000 158.2000 58.0000 159.9000 ;
	    RECT 57.6000 157.9000 58.6000 158.2000 ;
	    RECT 53.4000 157.5000 53.8000 157.9000 ;
	    RECT 55.5000 157.6000 55.8000 157.9000 ;
	    RECT 55.1000 157.3000 56.9000 157.6000 ;
	    RECT 58.2000 157.5000 58.6000 157.9000 ;
	    RECT 55.1000 157.2000 55.5000 157.3000 ;
	    RECT 56.5000 157.2000 56.9000 157.3000 ;
	    RECT 53.0000 156.6000 53.7000 157.0000 ;
	    RECT 53.4000 156.1000 53.7000 156.6000 ;
	    RECT 54.5000 156.5000 55.6000 156.8000 ;
	    RECT 54.5000 156.4000 54.9000 156.5000 ;
	    RECT 53.4000 155.8000 54.6000 156.1000 ;
	    RECT 50.2000 154.8000 50.6000 155.6000 ;
	    RECT 51.0000 155.3000 53.1000 155.6000 ;
	    RECT 49.4000 153.8000 49.8000 154.2000 ;
	    RECT 48.6000 153.1000 49.0000 153.2000 ;
	    RECT 47.8000 152.8000 49.0000 153.1000 ;
	    RECT 47.8000 151.1000 48.2000 152.8000 ;
	    RECT 48.6000 152.4000 49.0000 152.8000 ;
	    RECT 49.5000 152.1000 49.8000 153.8000 ;
	    RECT 49.4000 151.1000 49.8000 152.1000 ;
	    RECT 51.0000 153.6000 51.4000 155.3000 ;
	    RECT 52.7000 155.2000 53.1000 155.3000 ;
	    RECT 51.9000 154.9000 52.3000 155.0000 ;
	    RECT 51.9000 154.6000 53.8000 154.9000 ;
	    RECT 53.4000 154.5000 53.8000 154.6000 ;
	    RECT 54.3000 154.2000 54.6000 155.8000 ;
	    RECT 55.3000 155.9000 55.6000 156.5000 ;
	    RECT 55.9000 156.5000 56.3000 156.6000 ;
	    RECT 58.2000 156.5000 58.6000 156.6000 ;
	    RECT 55.9000 156.2000 58.6000 156.5000 ;
	    RECT 55.3000 155.7000 57.7000 155.9000 ;
	    RECT 59.8000 155.7000 60.2000 159.9000 ;
	    RECT 55.3000 155.6000 60.2000 155.7000 ;
	    RECT 57.3000 155.5000 60.2000 155.6000 ;
	    RECT 57.4000 155.4000 60.2000 155.5000 ;
	    RECT 62.2000 155.7000 62.6000 159.9000 ;
	    RECT 64.4000 158.2000 64.8000 159.9000 ;
	    RECT 63.8000 157.9000 64.8000 158.2000 ;
	    RECT 66.6000 157.9000 67.0000 159.9000 ;
	    RECT 68.7000 157.9000 69.3000 159.9000 ;
	    RECT 63.8000 157.5000 64.2000 157.9000 ;
	    RECT 66.6000 157.6000 66.9000 157.9000 ;
	    RECT 65.5000 157.3000 67.3000 157.6000 ;
	    RECT 68.6000 157.5000 69.0000 157.9000 ;
	    RECT 65.5000 157.2000 65.9000 157.3000 ;
	    RECT 66.9000 157.2000 67.3000 157.3000 ;
	    RECT 63.8000 156.5000 64.2000 156.6000 ;
	    RECT 66.1000 156.5000 66.5000 156.6000 ;
	    RECT 63.8000 156.2000 66.5000 156.5000 ;
	    RECT 66.8000 156.5000 67.9000 156.8000 ;
	    RECT 66.8000 155.9000 67.1000 156.5000 ;
	    RECT 67.5000 156.4000 67.9000 156.5000 ;
	    RECT 68.7000 156.6000 69.4000 157.0000 ;
	    RECT 68.7000 156.1000 69.0000 156.6000 ;
	    RECT 64.7000 155.7000 67.1000 155.9000 ;
	    RECT 62.2000 155.6000 67.1000 155.7000 ;
	    RECT 67.8000 155.8000 69.0000 156.1000 ;
	    RECT 62.2000 155.5000 65.1000 155.6000 ;
	    RECT 62.2000 155.4000 65.0000 155.5000 ;
	    RECT 56.6000 155.1000 57.0000 155.2000 ;
	    RECT 65.4000 155.1000 65.8000 155.2000 ;
	    RECT 56.6000 154.8000 59.1000 155.1000 ;
	    RECT 58.7000 154.7000 59.1000 154.8000 ;
	    RECT 63.3000 154.8000 65.8000 155.1000 ;
	    RECT 63.3000 154.7000 63.7000 154.8000 ;
	    RECT 64.6000 154.7000 65.0000 154.8000 ;
	    RECT 57.9000 154.2000 58.3000 154.3000 ;
	    RECT 64.1000 154.2000 64.5000 154.3000 ;
	    RECT 67.8000 154.2000 68.1000 155.8000 ;
	    RECT 71.0000 155.6000 71.4000 159.9000 ;
	    RECT 72.6000 156.4000 73.0000 159.9000 ;
	    RECT 69.3000 155.3000 71.4000 155.6000 ;
	    RECT 69.3000 155.2000 69.7000 155.3000 ;
	    RECT 70.1000 154.9000 70.5000 155.0000 ;
	    RECT 68.6000 154.6000 70.5000 154.9000 ;
	    RECT 68.6000 154.5000 69.0000 154.6000 ;
	    RECT 54.3000 154.1000 59.8000 154.2000 ;
	    RECT 62.6000 154.1000 68.1000 154.2000 ;
	    RECT 54.3000 153.9000 68.1000 154.1000 ;
	    RECT 54.5000 153.8000 54.9000 153.9000 ;
	    RECT 51.0000 153.3000 52.9000 153.6000 ;
	    RECT 51.0000 151.1000 51.4000 153.3000 ;
	    RECT 52.5000 153.2000 52.9000 153.3000 ;
	    RECT 57.4000 152.8000 57.7000 153.9000 ;
	    RECT 59.0000 153.8000 63.4000 153.9000 ;
	    RECT 56.5000 152.7000 56.9000 152.8000 ;
	    RECT 53.4000 152.1000 53.8000 152.5000 ;
	    RECT 55.5000 152.4000 56.9000 152.7000 ;
	    RECT 57.4000 152.4000 57.8000 152.8000 ;
	    RECT 55.5000 152.1000 55.8000 152.4000 ;
	    RECT 58.2000 152.1000 58.6000 152.5000 ;
	    RECT 53.1000 151.8000 53.8000 152.1000 ;
	    RECT 53.1000 151.1000 53.7000 151.8000 ;
	    RECT 55.4000 151.1000 55.8000 152.1000 ;
	    RECT 57.6000 151.8000 58.6000 152.1000 ;
	    RECT 57.6000 151.1000 58.0000 151.8000 ;
	    RECT 59.8000 151.1000 60.2000 153.5000 ;
	    RECT 62.2000 151.1000 62.6000 153.5000 ;
	    RECT 64.7000 152.8000 65.0000 153.9000 ;
	    RECT 65.4000 153.8000 65.8000 153.9000 ;
	    RECT 66.2000 153.8000 66.6000 153.9000 ;
	    RECT 67.5000 153.8000 67.9000 153.9000 ;
	    RECT 71.0000 153.6000 71.4000 155.3000 ;
	    RECT 69.5000 153.3000 71.4000 153.6000 ;
	    RECT 69.5000 153.2000 69.9000 153.3000 ;
	    RECT 63.8000 152.1000 64.2000 152.5000 ;
	    RECT 64.6000 152.4000 65.0000 152.8000 ;
	    RECT 65.5000 152.7000 65.9000 152.8000 ;
	    RECT 65.5000 152.4000 66.9000 152.7000 ;
	    RECT 66.6000 152.1000 66.9000 152.4000 ;
	    RECT 68.6000 152.1000 69.0000 152.5000 ;
	    RECT 63.8000 151.8000 64.8000 152.1000 ;
	    RECT 64.4000 151.1000 64.8000 151.8000 ;
	    RECT 66.6000 151.1000 67.0000 152.1000 ;
	    RECT 68.6000 151.8000 69.3000 152.1000 ;
	    RECT 68.7000 151.1000 69.3000 151.8000 ;
	    RECT 71.0000 151.1000 71.4000 153.3000 ;
	    RECT 72.5000 155.9000 73.0000 156.4000 ;
	    RECT 74.2000 156.2000 74.6000 159.9000 ;
	    RECT 73.3000 155.9000 74.6000 156.2000 ;
	    RECT 75.0000 156.2000 75.4000 159.9000 ;
	    RECT 75.0000 155.9000 76.1000 156.2000 ;
	    RECT 72.5000 154.2000 72.8000 155.9000 ;
	    RECT 73.3000 154.9000 73.6000 155.9000 ;
	    RECT 75.8000 155.6000 76.1000 155.9000 ;
	    RECT 75.8000 155.2000 76.4000 155.6000 ;
	    RECT 73.1000 154.5000 73.6000 154.9000 ;
	    RECT 72.5000 153.8000 73.0000 154.2000 ;
	    RECT 72.5000 153.1000 72.8000 153.8000 ;
	    RECT 73.3000 153.7000 73.6000 154.5000 ;
	    RECT 75.0000 154.4000 75.4000 155.2000 ;
	    RECT 75.8000 153.7000 76.1000 155.2000 ;
	    RECT 73.3000 153.4000 74.6000 153.7000 ;
	    RECT 72.5000 152.8000 73.0000 153.1000 ;
	    RECT 72.6000 151.1000 73.0000 152.8000 ;
	    RECT 74.2000 151.1000 74.6000 153.4000 ;
	    RECT 75.0000 153.4000 76.1000 153.7000 ;
	    RECT 77.4000 153.8000 77.8000 154.2000 ;
	    RECT 75.0000 151.1000 75.4000 153.4000 ;
	    RECT 77.4000 153.2000 77.7000 153.8000 ;
	    RECT 77.4000 152.4000 77.8000 153.2000 ;
	    RECT 78.2000 153.1000 78.6000 159.9000 ;
	    RECT 80.3000 156.3000 80.7000 159.9000 ;
	    RECT 82.2000 156.4000 82.6000 159.9000 ;
	    RECT 79.8000 155.9000 80.7000 156.3000 ;
	    RECT 82.1000 155.9000 82.6000 156.4000 ;
	    RECT 83.8000 156.2000 84.2000 159.9000 ;
	    RECT 85.0000 156.8000 85.4000 157.2000 ;
	    RECT 85.0000 156.2000 85.3000 156.8000 ;
	    RECT 85.7000 156.2000 86.1000 159.9000 ;
	    RECT 82.9000 155.9000 84.2000 156.2000 ;
	    RECT 84.6000 155.9000 85.3000 156.2000 ;
	    RECT 85.6000 155.9000 86.1000 156.2000 ;
	    RECT 88.1000 159.2000 88.5000 159.9000 ;
	    RECT 91.5000 159.2000 91.9000 159.9000 ;
	    RECT 88.1000 158.8000 89.0000 159.2000 ;
	    RECT 91.0000 158.8000 91.9000 159.2000 ;
	    RECT 88.1000 156.3000 88.5000 158.8000 ;
	    RECT 88.1000 155.9000 89.0000 156.3000 ;
	    RECT 91.5000 156.2000 91.9000 158.8000 ;
	    RECT 91.5000 155.9000 92.0000 156.2000 ;
	    RECT 79.9000 154.2000 80.2000 155.9000 ;
	    RECT 79.8000 153.8000 80.2000 154.2000 ;
	    RECT 80.6000 154.8000 81.0000 155.6000 ;
	    RECT 80.6000 154.1000 80.9000 154.8000 ;
	    RECT 82.1000 154.2000 82.4000 155.9000 ;
	    RECT 82.9000 154.9000 83.2000 155.9000 ;
	    RECT 84.6000 155.8000 85.0000 155.9000 ;
	    RECT 82.7000 154.5000 83.2000 154.9000 ;
	    RECT 82.1000 154.1000 82.6000 154.2000 ;
	    RECT 80.6000 153.8000 82.6000 154.1000 ;
	    RECT 79.0000 153.1000 79.4000 153.2000 ;
	    RECT 78.2000 152.8000 79.4000 153.1000 ;
	    RECT 78.2000 151.1000 78.6000 152.8000 ;
	    RECT 79.0000 152.4000 79.4000 152.8000 ;
	    RECT 79.9000 152.2000 80.2000 153.8000 ;
	    RECT 82.1000 153.1000 82.4000 153.8000 ;
	    RECT 82.9000 153.7000 83.2000 154.5000 ;
	    RECT 83.7000 155.1000 84.2000 155.2000 ;
	    RECT 85.6000 155.1000 85.9000 155.9000 ;
	    RECT 83.7000 154.8000 85.9000 155.1000 ;
	    RECT 83.7000 154.4000 84.1000 154.8000 ;
	    RECT 85.6000 154.2000 85.9000 154.8000 ;
	    RECT 87.8000 154.8000 88.2000 155.6000 ;
	    RECT 84.6000 153.8000 85.9000 154.2000 ;
	    RECT 87.0000 154.1000 87.4000 154.2000 ;
	    RECT 87.8000 154.1000 88.1000 154.8000 ;
	    RECT 86.6000 153.8000 88.1000 154.1000 ;
	    RECT 88.6000 154.2000 88.9000 155.9000 ;
	    RECT 91.0000 154.4000 91.4000 155.2000 ;
	    RECT 91.7000 154.2000 92.0000 155.9000 ;
	    RECT 94.2000 155.1000 94.6000 159.9000 ;
	    RECT 95.0000 155.8000 95.4000 156.6000 ;
	    RECT 96.1000 156.3000 96.5000 159.9000 ;
	    RECT 96.1000 155.9000 97.0000 156.3000 ;
	    RECT 99.0000 156.1000 99.4000 159.9000 ;
	    RECT 99.8000 156.8000 100.2000 157.2000 ;
	    RECT 99.8000 156.1000 100.1000 156.8000 ;
	    RECT 95.8000 155.1000 96.2000 155.6000 ;
	    RECT 94.2000 154.8000 96.2000 155.1000 ;
	    RECT 88.6000 153.8000 89.0000 154.2000 ;
	    RECT 90.2000 154.1000 90.6000 154.2000 ;
	    RECT 90.2000 153.8000 91.0000 154.1000 ;
	    RECT 91.7000 153.8000 93.0000 154.2000 ;
	    RECT 82.9000 153.4000 84.2000 153.7000 ;
	    RECT 82.1000 152.8000 82.6000 153.1000 ;
	    RECT 79.8000 151.1000 80.2000 152.2000 ;
	    RECT 82.2000 151.1000 82.6000 152.8000 ;
	    RECT 83.8000 151.1000 84.2000 153.4000 ;
	    RECT 84.7000 153.1000 85.0000 153.8000 ;
	    RECT 86.6000 153.6000 87.0000 153.8000 ;
	    RECT 85.5000 153.1000 87.3000 153.3000 ;
	    RECT 84.6000 151.1000 85.0000 153.1000 ;
	    RECT 85.4000 153.0000 87.4000 153.1000 ;
	    RECT 85.4000 151.1000 85.8000 153.0000 ;
	    RECT 87.0000 151.1000 87.4000 153.0000 ;
	    RECT 88.6000 152.1000 88.9000 153.8000 ;
	    RECT 90.6000 153.6000 91.0000 153.8000 ;
	    RECT 90.3000 153.1000 92.1000 153.3000 ;
	    RECT 92.6000 153.1000 92.9000 153.8000 ;
	    RECT 93.4000 153.4000 93.8000 154.2000 ;
	    RECT 94.2000 153.1000 94.6000 154.8000 ;
	    RECT 96.6000 154.2000 96.9000 155.9000 ;
	    RECT 99.0000 155.8000 100.1000 156.1000 ;
	    RECT 96.6000 153.8000 97.0000 154.2000 ;
	    RECT 95.8000 153.1000 96.2000 153.2000 ;
	    RECT 96.6000 153.1000 96.9000 153.8000 ;
	    RECT 90.2000 153.0000 92.2000 153.1000 ;
	    RECT 88.6000 151.1000 89.0000 152.1000 ;
	    RECT 90.2000 151.1000 90.6000 153.0000 ;
	    RECT 91.8000 151.1000 92.2000 153.0000 ;
	    RECT 92.6000 151.1000 93.0000 153.1000 ;
	    RECT 94.2000 152.8000 95.1000 153.1000 ;
	    RECT 95.8000 152.8000 96.9000 153.1000 ;
	    RECT 94.7000 151.1000 95.1000 152.8000 ;
	    RECT 96.6000 152.2000 96.9000 152.8000 ;
	    RECT 97.4000 153.1000 97.8000 153.2000 ;
	    RECT 98.2000 153.1000 98.6000 153.2000 ;
	    RECT 97.4000 152.8000 98.6000 153.1000 ;
	    RECT 97.4000 152.4000 97.8000 152.8000 ;
	    RECT 98.2000 152.4000 98.6000 152.8000 ;
	    RECT 96.6000 151.1000 97.0000 152.2000 ;
	    RECT 99.0000 151.1000 99.4000 155.8000 ;
	    RECT 99.8000 153.4000 100.2000 154.2000 ;
	    RECT 100.6000 153.1000 101.0000 159.9000 ;
	    RECT 101.4000 155.8000 101.8000 156.6000 ;
	    RECT 102.5000 156.3000 102.9000 159.9000 ;
	    RECT 105.0000 156.8000 105.4000 157.2000 ;
	    RECT 102.5000 155.9000 103.4000 156.3000 ;
	    RECT 105.0000 156.2000 105.3000 156.8000 ;
	    RECT 105.7000 156.2000 106.1000 159.9000 ;
	    RECT 103.0000 155.8000 103.4000 155.9000 ;
	    RECT 104.6000 155.9000 105.3000 156.2000 ;
	    RECT 105.6000 155.9000 106.1000 156.2000 ;
	    RECT 104.6000 155.8000 105.0000 155.9000 ;
	    RECT 101.4000 155.1000 101.7000 155.8000 ;
	    RECT 102.2000 155.1000 102.6000 155.6000 ;
	    RECT 101.4000 154.8000 102.6000 155.1000 ;
	    RECT 103.0000 154.2000 103.3000 155.8000 ;
	    RECT 105.6000 154.2000 105.9000 155.9000 ;
	    RECT 107.8000 155.8000 108.2000 156.6000 ;
	    RECT 106.2000 155.1000 106.6000 155.2000 ;
	    RECT 107.8000 155.1000 108.2000 155.2000 ;
	    RECT 106.2000 154.8000 108.2000 155.1000 ;
	    RECT 106.2000 154.4000 106.6000 154.8000 ;
	    RECT 103.0000 153.8000 103.4000 154.2000 ;
	    RECT 104.6000 153.8000 105.9000 154.2000 ;
	    RECT 102.2000 153.1000 102.6000 153.2000 ;
	    RECT 100.6000 152.8000 102.6000 153.1000 ;
	    RECT 101.1000 151.1000 101.5000 152.8000 ;
	    RECT 103.0000 152.1000 103.3000 153.8000 ;
	    RECT 103.8000 153.1000 104.2000 153.2000 ;
	    RECT 104.7000 153.1000 105.0000 153.8000 ;
	    RECT 105.5000 153.1000 107.3000 153.3000 ;
	    RECT 108.6000 153.1000 109.0000 159.9000 ;
	    RECT 103.8000 152.8000 105.0000 153.1000 ;
	    RECT 103.8000 152.4000 104.2000 152.8000 ;
	    RECT 103.0000 151.1000 103.4000 152.1000 ;
	    RECT 104.6000 151.1000 105.0000 152.8000 ;
	    RECT 105.4000 153.0000 107.4000 153.1000 ;
	    RECT 105.4000 151.1000 105.8000 153.0000 ;
	    RECT 107.0000 151.1000 107.4000 153.0000 ;
	    RECT 108.1000 152.8000 109.0000 153.1000 ;
	    RECT 111.8000 155.6000 112.2000 159.9000 ;
	    RECT 113.9000 157.9000 114.5000 159.9000 ;
	    RECT 116.2000 157.9000 116.6000 159.9000 ;
	    RECT 118.4000 158.2000 118.8000 159.9000 ;
	    RECT 118.4000 157.9000 119.4000 158.2000 ;
	    RECT 114.2000 157.5000 114.6000 157.9000 ;
	    RECT 116.3000 157.6000 116.6000 157.9000 ;
	    RECT 115.9000 157.3000 117.7000 157.6000 ;
	    RECT 119.0000 157.5000 119.4000 157.9000 ;
	    RECT 115.9000 157.2000 116.3000 157.3000 ;
	    RECT 117.3000 157.2000 117.7000 157.3000 ;
	    RECT 113.8000 156.6000 114.5000 157.0000 ;
	    RECT 114.2000 156.1000 114.5000 156.6000 ;
	    RECT 115.3000 156.5000 116.4000 156.8000 ;
	    RECT 115.3000 156.4000 115.7000 156.5000 ;
	    RECT 114.2000 155.8000 115.4000 156.1000 ;
	    RECT 111.8000 155.3000 113.9000 155.6000 ;
	    RECT 111.8000 153.6000 112.2000 155.3000 ;
	    RECT 113.5000 155.2000 113.9000 155.3000 ;
	    RECT 112.7000 154.9000 113.1000 155.0000 ;
	    RECT 112.7000 154.6000 114.6000 154.9000 ;
	    RECT 114.2000 154.5000 114.6000 154.6000 ;
	    RECT 115.1000 154.2000 115.4000 155.8000 ;
	    RECT 116.1000 155.9000 116.4000 156.5000 ;
	    RECT 116.7000 156.5000 117.1000 156.6000 ;
	    RECT 119.0000 156.5000 119.4000 156.6000 ;
	    RECT 116.7000 156.2000 119.4000 156.5000 ;
	    RECT 116.1000 155.7000 118.5000 155.9000 ;
	    RECT 120.6000 155.7000 121.0000 159.9000 ;
	    RECT 123.0000 156.2000 123.4000 159.9000 ;
	    RECT 116.1000 155.6000 121.0000 155.7000 ;
	    RECT 122.3000 155.9000 123.4000 156.2000 ;
	    RECT 122.3000 155.6000 122.6000 155.9000 ;
	    RECT 118.1000 155.5000 121.0000 155.6000 ;
	    RECT 118.2000 155.4000 121.0000 155.5000 ;
	    RECT 122.0000 155.2000 122.6000 155.6000 ;
	    RECT 123.8000 155.7000 124.2000 159.9000 ;
	    RECT 126.0000 158.2000 126.4000 159.9000 ;
	    RECT 125.4000 157.9000 126.4000 158.2000 ;
	    RECT 128.2000 157.9000 128.6000 159.9000 ;
	    RECT 130.3000 157.9000 130.9000 159.9000 ;
	    RECT 125.4000 157.5000 125.8000 157.9000 ;
	    RECT 128.2000 157.6000 128.5000 157.9000 ;
	    RECT 127.1000 157.3000 128.9000 157.6000 ;
	    RECT 130.2000 157.5000 130.6000 157.9000 ;
	    RECT 127.1000 157.2000 127.5000 157.3000 ;
	    RECT 128.5000 157.2000 128.9000 157.3000 ;
	    RECT 125.4000 156.5000 125.8000 156.6000 ;
	    RECT 127.7000 156.5000 128.1000 156.6000 ;
	    RECT 125.4000 156.2000 128.1000 156.5000 ;
	    RECT 128.4000 156.5000 129.5000 156.8000 ;
	    RECT 128.4000 155.9000 128.7000 156.5000 ;
	    RECT 129.1000 156.4000 129.5000 156.5000 ;
	    RECT 130.3000 156.6000 131.0000 157.0000 ;
	    RECT 130.3000 156.1000 130.6000 156.6000 ;
	    RECT 126.3000 155.7000 128.7000 155.9000 ;
	    RECT 123.8000 155.6000 128.7000 155.7000 ;
	    RECT 129.4000 155.8000 130.6000 156.1000 ;
	    RECT 123.8000 155.5000 126.7000 155.6000 ;
	    RECT 123.8000 155.4000 126.6000 155.5000 ;
	    RECT 129.4000 155.2000 129.7000 155.8000 ;
	    RECT 132.6000 155.6000 133.0000 159.9000 ;
	    RECT 130.9000 155.3000 133.0000 155.6000 ;
	    RECT 133.4000 155.6000 133.8000 159.9000 ;
	    RECT 135.5000 157.2000 135.9000 159.9000 ;
	    RECT 135.5000 156.8000 136.2000 157.2000 ;
	    RECT 135.5000 156.2000 135.9000 156.8000 ;
	    RECT 135.5000 155.9000 136.2000 156.2000 ;
	    RECT 136.6000 155.9000 137.0000 159.9000 ;
	    RECT 137.4000 156.2000 137.8000 159.9000 ;
	    RECT 139.0000 156.2000 139.4000 159.9000 ;
	    RECT 137.4000 155.9000 139.4000 156.2000 ;
	    RECT 133.4000 155.4000 135.4000 155.6000 ;
	    RECT 133.4000 155.3000 135.5000 155.4000 ;
	    RECT 130.9000 155.2000 131.3000 155.3000 ;
	    RECT 117.4000 155.1000 117.8000 155.2000 ;
	    RECT 117.4000 154.8000 119.9000 155.1000 ;
	    RECT 119.5000 154.7000 119.9000 154.8000 ;
	    RECT 118.7000 154.2000 119.1000 154.3000 ;
	    RECT 115.1000 153.9000 120.6000 154.2000 ;
	    RECT 115.3000 153.8000 115.7000 153.9000 ;
	    RECT 111.8000 153.3000 113.7000 153.6000 ;
	    RECT 108.1000 152.2000 108.5000 152.8000 ;
	    RECT 107.8000 151.8000 108.5000 152.2000 ;
	    RECT 108.1000 151.1000 108.5000 151.8000 ;
	    RECT 111.8000 151.1000 112.2000 153.3000 ;
	    RECT 113.3000 153.2000 113.7000 153.3000 ;
	    RECT 118.2000 152.8000 118.5000 153.9000 ;
	    RECT 119.8000 153.8000 120.6000 153.9000 ;
	    RECT 122.3000 153.7000 122.6000 155.2000 ;
	    RECT 123.0000 154.4000 123.4000 155.2000 ;
	    RECT 127.0000 155.1000 127.4000 155.2000 ;
	    RECT 124.9000 154.8000 127.4000 155.1000 ;
	    RECT 129.4000 154.8000 129.8000 155.2000 ;
	    RECT 131.7000 154.9000 132.1000 155.0000 ;
	    RECT 124.9000 154.7000 125.3000 154.8000 ;
	    RECT 125.7000 154.2000 126.1000 154.3000 ;
	    RECT 129.4000 154.2000 129.7000 154.8000 ;
	    RECT 130.2000 154.6000 132.1000 154.9000 ;
	    RECT 130.2000 154.5000 130.6000 154.6000 ;
	    RECT 124.2000 153.9000 129.7000 154.2000 ;
	    RECT 124.2000 153.8000 125.0000 153.9000 ;
	    RECT 117.3000 152.7000 117.7000 152.8000 ;
	    RECT 114.2000 152.1000 114.6000 152.5000 ;
	    RECT 116.3000 152.4000 117.7000 152.7000 ;
	    RECT 118.2000 152.4000 118.6000 152.8000 ;
	    RECT 116.3000 152.1000 116.6000 152.4000 ;
	    RECT 119.0000 152.1000 119.4000 152.5000 ;
	    RECT 113.9000 151.8000 114.6000 152.1000 ;
	    RECT 113.9000 151.1000 114.5000 151.8000 ;
	    RECT 116.2000 151.1000 116.6000 152.1000 ;
	    RECT 118.4000 151.8000 119.4000 152.1000 ;
	    RECT 118.4000 151.1000 118.8000 151.8000 ;
	    RECT 120.6000 151.1000 121.0000 153.5000 ;
	    RECT 122.3000 153.4000 123.4000 153.7000 ;
	    RECT 123.0000 151.1000 123.4000 153.4000 ;
	    RECT 123.8000 151.1000 124.2000 153.5000 ;
	    RECT 126.3000 152.8000 126.6000 153.9000 ;
	    RECT 129.1000 153.8000 129.5000 153.9000 ;
	    RECT 132.6000 153.6000 133.0000 155.3000 ;
	    RECT 135.1000 155.0000 135.5000 155.3000 ;
	    RECT 135.9000 155.2000 136.2000 155.9000 ;
	    RECT 136.7000 155.2000 137.0000 155.9000 ;
	    RECT 138.6000 155.2000 139.0000 155.4000 ;
	    RECT 134.4000 154.2000 134.8000 154.6000 ;
	    RECT 134.2000 153.8000 134.7000 154.2000 ;
	    RECT 131.1000 153.3000 133.0000 153.6000 ;
	    RECT 135.2000 153.5000 135.5000 155.0000 ;
	    RECT 135.8000 154.8000 136.2000 155.2000 ;
	    RECT 136.6000 154.9000 137.8000 155.2000 ;
	    RECT 138.6000 155.1000 139.4000 155.2000 ;
	    RECT 139.8000 155.1000 140.2000 159.9000 ;
	    RECT 141.4000 155.7000 141.8000 159.9000 ;
	    RECT 143.6000 158.2000 144.0000 159.9000 ;
	    RECT 143.0000 157.9000 144.0000 158.2000 ;
	    RECT 145.8000 157.9000 146.2000 159.9000 ;
	    RECT 147.9000 157.9000 148.5000 159.9000 ;
	    RECT 143.0000 157.5000 143.4000 157.9000 ;
	    RECT 145.8000 157.6000 146.1000 157.9000 ;
	    RECT 144.7000 157.3000 146.5000 157.6000 ;
	    RECT 147.8000 157.5000 148.2000 157.9000 ;
	    RECT 144.7000 157.2000 145.1000 157.3000 ;
	    RECT 146.1000 157.2000 146.5000 157.3000 ;
	    RECT 143.0000 156.5000 143.4000 156.6000 ;
	    RECT 145.3000 156.5000 145.7000 156.6000 ;
	    RECT 143.0000 156.2000 145.7000 156.5000 ;
	    RECT 146.0000 156.5000 147.1000 156.8000 ;
	    RECT 146.0000 155.9000 146.3000 156.5000 ;
	    RECT 146.7000 156.4000 147.1000 156.5000 ;
	    RECT 147.9000 156.6000 148.6000 157.0000 ;
	    RECT 147.9000 156.1000 148.2000 156.6000 ;
	    RECT 143.9000 155.7000 146.3000 155.9000 ;
	    RECT 141.4000 155.6000 146.3000 155.7000 ;
	    RECT 147.0000 155.8000 148.2000 156.1000 ;
	    RECT 141.4000 155.5000 144.3000 155.6000 ;
	    RECT 141.4000 155.4000 144.2000 155.5000 ;
	    RECT 147.0000 155.2000 147.3000 155.8000 ;
	    RECT 150.2000 155.6000 150.6000 159.9000 ;
	    RECT 151.0000 159.6000 153.0000 159.9000 ;
	    RECT 151.0000 155.9000 151.4000 159.6000 ;
	    RECT 151.8000 155.9000 152.2000 159.3000 ;
	    RECT 152.6000 156.2000 153.0000 159.6000 ;
	    RECT 154.2000 156.2000 154.6000 159.9000 ;
	    RECT 152.6000 155.9000 154.6000 156.2000 ;
	    RECT 155.0000 156.2000 155.4000 159.9000 ;
	    RECT 155.0000 155.9000 156.1000 156.2000 ;
	    RECT 151.9000 155.6000 152.2000 155.9000 ;
	    RECT 155.8000 155.6000 156.1000 155.9000 ;
	    RECT 159.0000 155.6000 159.4000 159.9000 ;
	    RECT 161.1000 157.9000 161.7000 159.9000 ;
	    RECT 163.4000 157.9000 163.8000 159.9000 ;
	    RECT 165.6000 158.2000 166.0000 159.9000 ;
	    RECT 165.6000 157.9000 166.6000 158.2000 ;
	    RECT 161.4000 157.5000 161.8000 157.9000 ;
	    RECT 163.5000 157.6000 163.8000 157.9000 ;
	    RECT 163.1000 157.3000 164.9000 157.6000 ;
	    RECT 166.2000 157.5000 166.6000 157.9000 ;
	    RECT 163.1000 157.2000 163.5000 157.3000 ;
	    RECT 164.5000 157.2000 164.9000 157.3000 ;
	    RECT 161.0000 156.6000 161.7000 157.0000 ;
	    RECT 161.4000 156.1000 161.7000 156.6000 ;
	    RECT 162.5000 156.5000 163.6000 156.8000 ;
	    RECT 162.5000 156.4000 162.9000 156.5000 ;
	    RECT 161.4000 155.8000 162.6000 156.1000 ;
	    RECT 148.5000 155.3000 150.6000 155.6000 ;
	    RECT 148.5000 155.2000 148.9000 155.3000 ;
	    RECT 144.6000 155.1000 145.0000 155.2000 ;
	    RECT 138.6000 154.9000 140.2000 155.1000 ;
	    RECT 136.6000 154.8000 137.0000 154.9000 ;
	    RECT 137.4000 154.8000 137.8000 154.9000 ;
	    RECT 139.0000 154.8000 140.2000 154.9000 ;
	    RECT 131.1000 153.2000 131.5000 153.3000 ;
	    RECT 125.4000 152.1000 125.8000 152.5000 ;
	    RECT 126.2000 152.4000 126.6000 152.8000 ;
	    RECT 127.1000 152.7000 127.5000 152.8000 ;
	    RECT 127.1000 152.4000 128.5000 152.7000 ;
	    RECT 128.2000 152.1000 128.5000 152.4000 ;
	    RECT 130.2000 152.1000 130.6000 152.5000 ;
	    RECT 125.4000 151.8000 126.4000 152.1000 ;
	    RECT 126.0000 151.1000 126.4000 151.8000 ;
	    RECT 128.2000 151.1000 128.6000 152.1000 ;
	    RECT 130.2000 151.8000 130.9000 152.1000 ;
	    RECT 130.3000 151.1000 130.9000 151.8000 ;
	    RECT 132.6000 151.1000 133.0000 153.3000 ;
	    RECT 134.3000 153.2000 135.5000 153.5000 ;
	    RECT 133.4000 152.4000 133.8000 153.2000 ;
	    RECT 134.3000 152.1000 134.6000 153.2000 ;
	    RECT 135.9000 153.1000 136.2000 154.8000 ;
	    RECT 134.2000 151.1000 134.6000 152.1000 ;
	    RECT 135.8000 151.1000 136.2000 153.1000 ;
	    RECT 136.6000 152.8000 137.0000 153.2000 ;
	    RECT 137.5000 153.1000 137.8000 154.8000 ;
	    RECT 138.2000 153.8000 138.6000 154.6000 ;
	    RECT 136.7000 152.4000 137.1000 152.8000 ;
	    RECT 137.4000 151.1000 137.8000 153.1000 ;
	    RECT 139.8000 151.1000 140.2000 154.8000 ;
	    RECT 142.5000 154.8000 145.0000 155.1000 ;
	    RECT 147.0000 154.8000 147.4000 155.2000 ;
	    RECT 149.3000 154.9000 149.7000 155.0000 ;
	    RECT 142.5000 154.7000 142.9000 154.8000 ;
	    RECT 143.8000 154.7000 144.2000 154.8000 ;
	    RECT 143.3000 154.2000 143.7000 154.3000 ;
	    RECT 147.0000 154.2000 147.3000 154.8000 ;
	    RECT 147.8000 154.6000 149.7000 154.9000 ;
	    RECT 147.8000 154.5000 148.2000 154.6000 ;
	    RECT 141.8000 153.9000 147.3000 154.2000 ;
	    RECT 141.8000 153.8000 142.6000 153.9000 ;
	    RECT 140.6000 152.4000 141.0000 153.2000 ;
	    RECT 141.4000 151.1000 141.8000 153.5000 ;
	    RECT 143.9000 152.8000 144.2000 153.9000 ;
	    RECT 146.7000 153.8000 147.1000 153.9000 ;
	    RECT 150.2000 153.6000 150.6000 155.3000 ;
	    RECT 151.0000 154.8000 151.4000 155.6000 ;
	    RECT 151.9000 155.3000 152.9000 155.6000 ;
	    RECT 152.6000 155.2000 152.9000 155.3000 ;
	    RECT 153.8000 155.2000 154.2000 155.4000 ;
	    RECT 155.8000 155.2000 156.4000 155.6000 ;
	    RECT 159.0000 155.3000 161.1000 155.6000 ;
	    RECT 152.6000 154.8000 153.0000 155.2000 ;
	    RECT 153.8000 154.9000 154.6000 155.2000 ;
	    RECT 154.2000 154.8000 154.6000 154.9000 ;
	    RECT 151.9000 154.4000 152.3000 154.8000 ;
	    RECT 151.9000 154.2000 152.2000 154.4000 ;
	    RECT 151.8000 153.8000 152.2000 154.2000 ;
	    RECT 148.7000 153.3000 150.6000 153.6000 ;
	    RECT 148.7000 153.2000 149.1000 153.3000 ;
	    RECT 143.0000 152.1000 143.4000 152.5000 ;
	    RECT 143.8000 152.4000 144.2000 152.8000 ;
	    RECT 144.7000 152.7000 145.1000 152.8000 ;
	    RECT 144.7000 152.4000 146.1000 152.7000 ;
	    RECT 145.8000 152.1000 146.1000 152.4000 ;
	    RECT 147.8000 152.1000 148.2000 152.5000 ;
	    RECT 143.0000 151.8000 144.0000 152.1000 ;
	    RECT 143.6000 151.1000 144.0000 151.8000 ;
	    RECT 145.8000 151.1000 146.2000 152.1000 ;
	    RECT 147.8000 151.8000 148.5000 152.1000 ;
	    RECT 147.9000 151.1000 148.5000 151.8000 ;
	    RECT 150.2000 151.1000 150.6000 153.3000 ;
	    RECT 152.6000 153.1000 152.9000 154.8000 ;
	    RECT 153.4000 153.8000 153.8000 154.6000 ;
	    RECT 155.0000 154.4000 155.4000 155.2000 ;
	    RECT 155.8000 153.7000 156.1000 155.2000 ;
	    RECT 155.0000 153.4000 156.1000 153.7000 ;
	    RECT 159.0000 153.6000 159.4000 155.3000 ;
	    RECT 160.7000 155.2000 161.1000 155.3000 ;
	    RECT 159.9000 154.9000 160.3000 155.0000 ;
	    RECT 159.9000 154.6000 161.8000 154.9000 ;
	    RECT 161.4000 154.5000 161.8000 154.6000 ;
	    RECT 162.3000 154.2000 162.6000 155.8000 ;
	    RECT 163.3000 155.9000 163.6000 156.5000 ;
	    RECT 163.9000 156.5000 164.3000 156.6000 ;
	    RECT 166.2000 156.5000 166.6000 156.6000 ;
	    RECT 163.9000 156.2000 166.6000 156.5000 ;
	    RECT 163.3000 155.7000 165.7000 155.9000 ;
	    RECT 167.8000 155.7000 168.2000 159.9000 ;
	    RECT 168.6000 155.9000 169.0000 159.9000 ;
	    RECT 169.4000 156.2000 169.8000 159.9000 ;
	    RECT 171.0000 156.2000 171.4000 159.9000 ;
	    RECT 172.2000 156.8000 172.6000 157.2000 ;
	    RECT 172.2000 156.2000 172.5000 156.8000 ;
	    RECT 172.9000 156.2000 173.3000 159.9000 ;
	    RECT 169.4000 155.9000 171.4000 156.2000 ;
	    RECT 171.8000 155.9000 172.5000 156.2000 ;
	    RECT 172.8000 155.9000 173.3000 156.2000 ;
	    RECT 175.3000 156.3000 175.7000 159.9000 ;
	    RECT 175.3000 155.9000 176.2000 156.3000 ;
	    RECT 163.3000 155.6000 168.2000 155.7000 ;
	    RECT 165.3000 155.5000 168.2000 155.6000 ;
	    RECT 165.4000 155.4000 168.2000 155.5000 ;
	    RECT 168.7000 155.2000 169.0000 155.9000 ;
	    RECT 171.8000 155.8000 172.2000 155.9000 ;
	    RECT 170.6000 155.2000 171.0000 155.4000 ;
	    RECT 164.6000 155.1000 165.0000 155.2000 ;
	    RECT 164.6000 154.8000 167.1000 155.1000 ;
	    RECT 165.4000 154.7000 165.8000 154.8000 ;
	    RECT 166.7000 154.7000 167.1000 154.8000 ;
	    RECT 168.6000 154.9000 169.8000 155.2000 ;
	    RECT 170.6000 155.1000 171.4000 155.2000 ;
	    RECT 172.8000 155.1000 173.1000 155.9000 ;
	    RECT 170.6000 154.9000 173.1000 155.1000 ;
	    RECT 168.6000 154.8000 169.0000 154.9000 ;
	    RECT 165.9000 154.2000 166.3000 154.3000 ;
	    RECT 168.6000 154.2000 168.9000 154.8000 ;
	    RECT 162.3000 153.9000 167.8000 154.2000 ;
	    RECT 162.5000 153.8000 162.9000 153.9000 ;
	    RECT 164.6000 153.8000 165.0000 153.9000 ;
	    RECT 152.3000 151.1000 153.1000 153.1000 ;
	    RECT 155.0000 151.1000 155.4000 153.4000 ;
	    RECT 159.0000 153.3000 160.9000 153.6000 ;
	    RECT 159.0000 151.1000 159.4000 153.3000 ;
	    RECT 160.5000 153.2000 160.9000 153.3000 ;
	    RECT 165.4000 152.8000 165.7000 153.9000 ;
	    RECT 167.0000 153.8000 167.8000 153.9000 ;
	    RECT 168.6000 153.8000 169.0000 154.2000 ;
	    RECT 164.5000 152.7000 164.9000 152.8000 ;
	    RECT 161.4000 152.1000 161.8000 152.5000 ;
	    RECT 163.5000 152.4000 164.9000 152.7000 ;
	    RECT 165.4000 152.4000 165.8000 152.8000 ;
	    RECT 163.5000 152.1000 163.8000 152.4000 ;
	    RECT 166.2000 152.1000 166.6000 152.5000 ;
	    RECT 161.1000 151.8000 161.8000 152.1000 ;
	    RECT 161.1000 151.1000 161.7000 151.8000 ;
	    RECT 163.4000 151.1000 163.8000 152.1000 ;
	    RECT 165.6000 151.8000 166.6000 152.1000 ;
	    RECT 165.6000 151.1000 166.0000 151.8000 ;
	    RECT 167.8000 151.1000 168.2000 153.5000 ;
	    RECT 168.6000 152.8000 169.0000 153.2000 ;
	    RECT 169.5000 153.1000 169.8000 154.9000 ;
	    RECT 171.0000 154.8000 173.1000 154.9000 ;
	    RECT 170.2000 153.8000 170.6000 154.6000 ;
	    RECT 172.8000 154.2000 173.1000 154.8000 ;
	    RECT 173.4000 154.4000 173.8000 155.2000 ;
	    RECT 175.0000 154.8000 175.4000 155.6000 ;
	    RECT 175.8000 155.1000 176.1000 155.9000 ;
	    RECT 177.4000 155.8000 177.8000 156.6000 ;
	    RECT 177.4000 155.1000 177.7000 155.8000 ;
	    RECT 175.8000 154.8000 177.7000 155.1000 ;
	    RECT 175.8000 154.2000 176.1000 154.8000 ;
	    RECT 171.8000 153.8000 173.1000 154.2000 ;
	    RECT 174.2000 154.1000 174.6000 154.2000 ;
	    RECT 175.0000 154.1000 175.4000 154.2000 ;
	    RECT 173.8000 153.8000 175.4000 154.1000 ;
	    RECT 175.8000 153.8000 176.2000 154.2000 ;
	    RECT 177.4000 154.1000 177.8000 154.2000 ;
	    RECT 178.2000 154.1000 178.6000 159.9000 ;
	    RECT 177.4000 153.8000 178.6000 154.1000 ;
	    RECT 171.9000 153.1000 172.2000 153.8000 ;
	    RECT 173.8000 153.6000 174.2000 153.8000 ;
	    RECT 172.7000 153.1000 174.5000 153.3000 ;
	    RECT 168.7000 152.4000 169.1000 152.8000 ;
	    RECT 169.4000 151.1000 169.8000 153.1000 ;
	    RECT 171.8000 151.1000 172.2000 153.1000 ;
	    RECT 172.6000 153.0000 174.6000 153.1000 ;
	    RECT 172.6000 151.1000 173.0000 153.0000 ;
	    RECT 174.2000 151.1000 174.6000 153.0000 ;
	    RECT 175.8000 152.1000 176.1000 153.8000 ;
	    RECT 176.6000 152.4000 177.0000 153.2000 ;
	    RECT 178.2000 153.1000 178.6000 153.8000 ;
	    RECT 179.0000 153.4000 179.4000 154.2000 ;
	    RECT 179.8000 153.4000 180.2000 154.2000 ;
	    RECT 177.7000 152.8000 178.6000 153.1000 ;
	    RECT 180.6000 153.1000 181.0000 159.9000 ;
	    RECT 181.4000 155.8000 181.8000 156.6000 ;
	    RECT 183.5000 156.3000 183.9000 159.9000 ;
	    RECT 183.0000 155.9000 183.9000 156.3000 ;
	    RECT 184.6000 155.9000 185.0000 159.9000 ;
	    RECT 185.4000 156.2000 185.8000 159.9000 ;
	    RECT 187.0000 156.2000 187.4000 159.9000 ;
	    RECT 188.2000 156.8000 188.6000 157.2000 ;
	    RECT 188.2000 156.2000 188.5000 156.8000 ;
	    RECT 188.9000 156.2000 189.3000 159.9000 ;
	    RECT 185.4000 155.9000 187.4000 156.2000 ;
	    RECT 187.8000 155.9000 188.5000 156.2000 ;
	    RECT 188.8000 155.9000 189.3000 156.2000 ;
	    RECT 191.3000 157.2000 191.7000 159.9000 ;
	    RECT 191.3000 156.8000 192.2000 157.2000 ;
	    RECT 191.3000 156.3000 191.7000 156.8000 ;
	    RECT 191.3000 155.9000 192.2000 156.3000 ;
	    RECT 194.7000 156.2000 195.1000 159.9000 ;
	    RECT 195.4000 156.8000 195.8000 157.2000 ;
	    RECT 195.5000 156.2000 195.8000 156.8000 ;
	    RECT 196.6000 156.2000 197.0000 159.9000 ;
	    RECT 198.2000 156.2000 198.6000 159.9000 ;
	    RECT 194.7000 155.9000 195.2000 156.2000 ;
	    RECT 195.5000 155.9000 196.2000 156.2000 ;
	    RECT 196.6000 155.9000 198.6000 156.2000 ;
	    RECT 199.0000 155.9000 199.4000 159.9000 ;
	    RECT 183.1000 154.2000 183.4000 155.9000 ;
	    RECT 183.8000 154.8000 184.2000 155.6000 ;
	    RECT 184.7000 155.2000 185.0000 155.9000 ;
	    RECT 187.8000 155.8000 188.2000 155.9000 ;
	    RECT 186.6000 155.2000 187.0000 155.4000 ;
	    RECT 184.6000 154.9000 185.8000 155.2000 ;
	    RECT 186.6000 155.1000 187.4000 155.2000 ;
	    RECT 188.8000 155.1000 189.1000 155.9000 ;
	    RECT 186.6000 154.9000 189.1000 155.1000 ;
	    RECT 184.6000 154.8000 185.0000 154.9000 ;
	    RECT 183.0000 153.8000 183.4000 154.2000 ;
	    RECT 180.6000 152.8000 181.5000 153.1000 ;
	    RECT 175.8000 151.1000 176.2000 152.1000 ;
	    RECT 177.7000 151.1000 178.1000 152.8000 ;
	    RECT 181.1000 152.2000 181.5000 152.8000 ;
	    RECT 182.2000 152.4000 182.6000 153.2000 ;
	    RECT 183.1000 153.1000 183.4000 153.8000 ;
	    RECT 183.8000 153.1000 184.2000 153.2000 ;
	    RECT 183.0000 152.8000 184.2000 153.1000 ;
	    RECT 184.6000 152.8000 185.0000 153.2000 ;
	    RECT 185.5000 153.1000 185.8000 154.9000 ;
	    RECT 187.0000 154.8000 189.1000 154.9000 ;
	    RECT 186.2000 154.1000 186.6000 154.6000 ;
	    RECT 188.8000 154.2000 189.1000 154.8000 ;
	    RECT 189.4000 154.4000 189.8000 155.2000 ;
	    RECT 191.0000 155.1000 191.4000 155.6000 ;
	    RECT 190.2000 154.8000 191.4000 155.1000 ;
	    RECT 187.0000 154.1000 187.4000 154.2000 ;
	    RECT 186.2000 153.8000 187.4000 154.1000 ;
	    RECT 187.8000 153.8000 189.1000 154.2000 ;
	    RECT 190.2000 154.2000 190.5000 154.8000 ;
	    RECT 191.8000 154.2000 192.1000 155.9000 ;
	    RECT 192.6000 155.1000 193.0000 155.2000 ;
	    RECT 194.2000 155.1000 194.6000 155.2000 ;
	    RECT 192.6000 154.8000 194.6000 155.1000 ;
	    RECT 194.2000 154.4000 194.6000 154.8000 ;
	    RECT 194.9000 155.1000 195.2000 155.9000 ;
	    RECT 195.8000 155.8000 196.2000 155.9000 ;
	    RECT 197.0000 155.2000 197.4000 155.4000 ;
	    RECT 199.0000 155.2000 199.3000 155.9000 ;
	    RECT 199.8000 155.8000 200.2000 156.6000 ;
	    RECT 196.6000 155.1000 197.4000 155.2000 ;
	    RECT 194.9000 154.9000 197.4000 155.1000 ;
	    RECT 198.2000 155.1000 199.4000 155.2000 ;
	    RECT 199.8000 155.1000 200.2000 155.2000 ;
	    RECT 198.2000 154.9000 200.2000 155.1000 ;
	    RECT 194.9000 154.8000 197.0000 154.9000 ;
	    RECT 194.9000 154.2000 195.2000 154.8000 ;
	    RECT 190.2000 154.1000 190.6000 154.2000 ;
	    RECT 189.8000 153.8000 190.6000 154.1000 ;
	    RECT 191.8000 153.8000 192.2000 154.2000 ;
	    RECT 193.4000 154.1000 193.8000 154.2000 ;
	    RECT 193.4000 153.8000 194.2000 154.1000 ;
	    RECT 194.9000 153.8000 196.2000 154.2000 ;
	    RECT 197.4000 153.8000 197.8000 154.6000 ;
	    RECT 187.9000 153.1000 188.2000 153.8000 ;
	    RECT 189.8000 153.6000 190.2000 153.8000 ;
	    RECT 188.7000 153.1000 190.5000 153.3000 ;
	    RECT 180.6000 151.8000 181.5000 152.2000 ;
	    RECT 183.1000 152.1000 183.4000 152.8000 ;
	    RECT 184.7000 152.4000 185.1000 152.8000 ;
	    RECT 181.1000 151.1000 181.5000 151.8000 ;
	    RECT 183.0000 151.1000 183.4000 152.1000 ;
	    RECT 185.4000 151.1000 185.8000 153.1000 ;
	    RECT 187.8000 151.1000 188.2000 153.1000 ;
	    RECT 188.6000 153.0000 190.6000 153.1000 ;
	    RECT 188.6000 151.1000 189.0000 153.0000 ;
	    RECT 190.2000 151.1000 190.6000 153.0000 ;
	    RECT 191.8000 152.1000 192.1000 153.8000 ;
	    RECT 193.8000 153.6000 194.2000 153.8000 ;
	    RECT 192.6000 152.4000 193.0000 153.2000 ;
	    RECT 193.5000 153.1000 195.3000 153.3000 ;
	    RECT 195.8000 153.1000 196.1000 153.8000 ;
	    RECT 198.2000 153.1000 198.5000 154.9000 ;
	    RECT 199.0000 154.8000 200.2000 154.9000 ;
	    RECT 199.8000 154.1000 200.2000 154.2000 ;
	    RECT 200.6000 154.1000 201.0000 159.9000 ;
	    RECT 202.2000 155.7000 202.6000 159.9000 ;
	    RECT 204.4000 158.2000 204.8000 159.9000 ;
	    RECT 203.8000 157.9000 204.8000 158.2000 ;
	    RECT 206.6000 157.9000 207.0000 159.9000 ;
	    RECT 208.7000 157.9000 209.3000 159.9000 ;
	    RECT 203.8000 157.5000 204.2000 157.9000 ;
	    RECT 206.6000 157.6000 206.9000 157.9000 ;
	    RECT 205.5000 157.3000 207.3000 157.6000 ;
	    RECT 208.6000 157.5000 209.0000 157.9000 ;
	    RECT 205.5000 157.2000 205.9000 157.3000 ;
	    RECT 206.9000 157.2000 207.3000 157.3000 ;
	    RECT 203.8000 156.5000 204.2000 156.6000 ;
	    RECT 206.1000 156.5000 206.5000 156.6000 ;
	    RECT 203.8000 156.2000 206.5000 156.5000 ;
	    RECT 206.8000 156.5000 207.9000 156.8000 ;
	    RECT 206.8000 155.9000 207.1000 156.5000 ;
	    RECT 207.5000 156.4000 207.9000 156.5000 ;
	    RECT 208.7000 156.6000 209.4000 157.0000 ;
	    RECT 208.7000 156.1000 209.0000 156.6000 ;
	    RECT 204.7000 155.7000 207.1000 155.9000 ;
	    RECT 202.2000 155.6000 207.1000 155.7000 ;
	    RECT 207.8000 155.8000 209.0000 156.1000 ;
	    RECT 202.2000 155.5000 205.1000 155.6000 ;
	    RECT 202.2000 155.4000 205.0000 155.5000 ;
	    RECT 205.4000 155.1000 205.8000 155.2000 ;
	    RECT 203.3000 154.8000 205.8000 155.1000 ;
	    RECT 203.3000 154.7000 203.7000 154.8000 ;
	    RECT 204.6000 154.7000 205.0000 154.8000 ;
	    RECT 204.1000 154.2000 204.5000 154.3000 ;
	    RECT 207.8000 154.2000 208.1000 155.8000 ;
	    RECT 211.0000 155.6000 211.4000 159.9000 ;
	    RECT 209.3000 155.3000 211.4000 155.6000 ;
	    RECT 209.3000 155.2000 209.7000 155.3000 ;
	    RECT 210.1000 154.9000 210.5000 155.0000 ;
	    RECT 208.6000 154.6000 210.5000 154.9000 ;
	    RECT 208.6000 154.5000 209.0000 154.6000 ;
	    RECT 199.8000 153.8000 201.0000 154.1000 ;
	    RECT 193.4000 153.0000 195.4000 153.1000 ;
	    RECT 191.8000 151.1000 192.2000 152.1000 ;
	    RECT 193.4000 151.1000 193.8000 153.0000 ;
	    RECT 195.0000 151.1000 195.4000 153.0000 ;
	    RECT 195.8000 151.1000 196.2000 153.1000 ;
	    RECT 198.2000 151.1000 198.6000 153.1000 ;
	    RECT 199.0000 152.8000 199.4000 153.2000 ;
	    RECT 200.6000 153.1000 201.0000 153.8000 ;
	    RECT 201.4000 153.4000 201.8000 154.2000 ;
	    RECT 202.6000 153.9000 208.1000 154.2000 ;
	    RECT 202.6000 153.8000 203.4000 153.9000 ;
	    RECT 200.1000 152.8000 201.0000 153.1000 ;
	    RECT 198.9000 152.4000 199.3000 152.8000 ;
	    RECT 200.1000 151.1000 200.5000 152.8000 ;
	    RECT 202.2000 151.1000 202.6000 153.5000 ;
	    RECT 204.7000 152.8000 205.0000 153.9000 ;
	    RECT 207.5000 153.8000 207.9000 153.9000 ;
	    RECT 211.0000 153.6000 211.4000 155.3000 ;
	    RECT 209.5000 153.3000 211.4000 153.6000 ;
	    RECT 209.5000 153.2000 209.9000 153.3000 ;
	    RECT 203.8000 152.1000 204.2000 152.5000 ;
	    RECT 204.6000 152.4000 205.0000 152.8000 ;
	    RECT 205.5000 152.7000 205.9000 152.8000 ;
	    RECT 205.5000 152.4000 206.9000 152.7000 ;
	    RECT 206.6000 152.1000 206.9000 152.4000 ;
	    RECT 208.6000 152.1000 209.0000 152.5000 ;
	    RECT 203.8000 151.8000 204.8000 152.1000 ;
	    RECT 204.4000 151.1000 204.8000 151.8000 ;
	    RECT 206.6000 151.1000 207.0000 152.1000 ;
	    RECT 208.6000 151.8000 209.3000 152.1000 ;
	    RECT 208.7000 151.1000 209.3000 151.8000 ;
	    RECT 211.0000 151.1000 211.4000 153.3000 ;
	    RECT 213.4000 155.9000 213.8000 159.9000 ;
	    RECT 215.0000 157.9000 215.4000 159.9000 ;
	    RECT 213.4000 155.2000 213.7000 155.9000 ;
	    RECT 215.0000 155.8000 215.3000 157.9000 ;
	    RECT 217.9000 157.2000 218.3000 159.9000 ;
	    RECT 217.9000 156.8000 218.6000 157.2000 ;
	    RECT 217.9000 156.3000 218.3000 156.8000 ;
	    RECT 217.4000 155.9000 218.3000 156.3000 ;
	    RECT 220.3000 156.2000 220.7000 159.9000 ;
	    RECT 221.0000 156.8000 221.4000 157.2000 ;
	    RECT 221.1000 156.2000 221.4000 156.8000 ;
	    RECT 223.5000 156.2000 223.9000 159.9000 ;
	    RECT 224.2000 156.8000 224.6000 157.2000 ;
	    RECT 224.3000 156.2000 224.6000 156.8000 ;
	    RECT 220.3000 155.9000 220.8000 156.2000 ;
	    RECT 221.1000 155.9000 221.8000 156.2000 ;
	    RECT 223.5000 155.9000 224.0000 156.2000 ;
	    RECT 224.3000 156.1000 225.0000 156.2000 ;
	    RECT 225.4000 156.1000 225.8000 159.9000 ;
	    RECT 224.3000 155.9000 225.8000 156.1000 ;
	    RECT 227.3000 156.3000 227.7000 159.9000 ;
	    RECT 227.3000 155.9000 228.2000 156.3000 ;
	    RECT 229.4000 156.2000 229.8000 159.9000 ;
	    RECT 231.0000 156.4000 231.4000 159.9000 ;
	    RECT 233.9000 159.2000 234.3000 159.9000 ;
	    RECT 233.4000 158.8000 234.3000 159.2000 ;
	    RECT 229.4000 155.9000 230.7000 156.2000 ;
	    RECT 231.0000 155.9000 231.5000 156.4000 ;
	    RECT 233.9000 156.3000 234.3000 158.8000 ;
	    RECT 233.4000 155.9000 234.3000 156.3000 ;
	    RECT 235.0000 156.2000 235.4000 159.9000 ;
	    RECT 235.8000 156.2000 236.2000 156.3000 ;
	    RECT 237.2000 156.2000 238.0000 159.9000 ;
	    RECT 235.0000 155.9000 236.2000 156.2000 ;
	    RECT 237.0000 155.9000 238.0000 156.2000 ;
	    RECT 239.1000 156.2000 239.5000 156.3000 ;
	    RECT 239.8000 156.2000 240.2000 159.9000 ;
	    RECT 239.1000 155.9000 240.2000 156.2000 ;
	    RECT 240.9000 159.2000 241.3000 159.9000 ;
	    RECT 243.3000 159.2000 243.7000 159.9000 ;
	    RECT 240.9000 158.8000 241.8000 159.2000 ;
	    RECT 243.3000 158.8000 244.2000 159.2000 ;
	    RECT 240.9000 156.3000 241.3000 158.8000 ;
	    RECT 243.3000 156.3000 243.7000 158.8000 ;
	    RECT 240.9000 155.9000 241.8000 156.3000 ;
	    RECT 243.3000 155.9000 244.2000 156.3000 ;
	    RECT 245.4000 156.2000 245.8000 159.9000 ;
	    RECT 247.0000 156.2000 247.4000 159.9000 ;
	    RECT 245.4000 155.9000 247.4000 156.2000 ;
	    RECT 247.8000 155.9000 248.2000 159.9000 ;
	    RECT 249.9000 156.3000 250.3000 159.9000 ;
	    RECT 249.4000 155.9000 250.3000 156.3000 ;
	    RECT 251.0000 155.9000 251.4000 159.9000 ;
	    RECT 251.8000 156.2000 252.2000 159.9000 ;
	    RECT 253.4000 156.2000 253.8000 159.9000 ;
	    RECT 255.5000 159.2000 255.9000 159.9000 ;
	    RECT 255.0000 158.8000 255.9000 159.2000 ;
	    RECT 251.8000 155.9000 253.8000 156.2000 ;
	    RECT 255.5000 156.2000 255.9000 158.8000 ;
	    RECT 256.2000 156.8000 256.6000 157.2000 ;
	    RECT 256.3000 156.2000 256.6000 156.8000 ;
	    RECT 257.7000 156.3000 258.1000 159.9000 ;
	    RECT 261.1000 156.3000 261.5000 159.9000 ;
	    RECT 255.5000 155.9000 256.0000 156.2000 ;
	    RECT 256.3000 155.9000 257.0000 156.2000 ;
	    RECT 257.7000 155.9000 258.6000 156.3000 ;
	    RECT 260.6000 155.9000 261.5000 156.3000 ;
	    RECT 214.1000 155.5000 215.3000 155.8000 ;
	    RECT 213.4000 154.8000 213.8000 155.2000 ;
	    RECT 213.4000 153.1000 213.7000 154.8000 ;
	    RECT 214.1000 153.8000 214.4000 155.5000 ;
	    RECT 215.0000 154.8000 215.4000 155.2000 ;
	    RECT 215.0000 154.4000 215.3000 154.8000 ;
	    RECT 214.8000 154.1000 215.3000 154.4000 ;
	    RECT 214.8000 154.0000 215.2000 154.1000 ;
	    RECT 215.8000 153.8000 216.2000 154.6000 ;
	    RECT 217.5000 154.2000 217.8000 155.9000 ;
	    RECT 218.2000 154.8000 218.6000 155.6000 ;
	    RECT 219.8000 154.4000 220.2000 155.2000 ;
	    RECT 220.5000 154.2000 220.8000 155.9000 ;
	    RECT 221.4000 155.8000 221.8000 155.9000 ;
	    RECT 222.2000 155.1000 222.6000 155.2000 ;
	    RECT 223.0000 155.1000 223.4000 155.2000 ;
	    RECT 222.2000 154.8000 223.4000 155.1000 ;
	    RECT 223.0000 154.4000 223.4000 154.8000 ;
	    RECT 223.7000 154.2000 224.0000 155.9000 ;
	    RECT 224.6000 155.8000 225.8000 155.9000 ;
	    RECT 217.4000 153.8000 217.8000 154.2000 ;
	    RECT 219.0000 154.1000 219.4000 154.2000 ;
	    RECT 219.0000 153.8000 219.8000 154.1000 ;
	    RECT 220.5000 153.8000 221.8000 154.2000 ;
	    RECT 222.2000 154.1000 222.6000 154.2000 ;
	    RECT 222.2000 153.8000 223.0000 154.1000 ;
	    RECT 223.7000 153.8000 225.0000 154.2000 ;
	    RECT 214.0000 153.7000 214.4000 153.8000 ;
	    RECT 214.0000 153.5000 215.5000 153.7000 ;
	    RECT 214.0000 153.4000 216.1000 153.5000 ;
	    RECT 215.2000 153.2000 216.1000 153.4000 ;
	    RECT 215.8000 153.1000 216.1000 153.2000 ;
	    RECT 213.4000 152.6000 214.1000 153.1000 ;
	    RECT 213.7000 152.2000 214.1000 152.6000 ;
	    RECT 213.4000 151.8000 214.1000 152.2000 ;
	    RECT 213.7000 151.1000 214.1000 151.8000 ;
	    RECT 215.8000 151.1000 216.2000 153.1000 ;
	    RECT 216.6000 152.4000 217.0000 153.2000 ;
	    RECT 217.5000 152.1000 217.8000 153.8000 ;
	    RECT 219.4000 153.6000 219.8000 153.8000 ;
	    RECT 219.1000 153.1000 220.9000 153.3000 ;
	    RECT 221.4000 153.1000 221.7000 153.8000 ;
	    RECT 222.6000 153.6000 223.0000 153.8000 ;
	    RECT 222.3000 153.1000 224.1000 153.3000 ;
	    RECT 224.6000 153.1000 224.9000 153.8000 ;
	    RECT 217.4000 151.1000 217.8000 152.1000 ;
	    RECT 219.0000 153.0000 221.0000 153.1000 ;
	    RECT 219.0000 151.1000 219.4000 153.0000 ;
	    RECT 220.6000 151.1000 221.0000 153.0000 ;
	    RECT 221.4000 151.1000 221.8000 153.1000 ;
	    RECT 222.2000 153.0000 224.2000 153.1000 ;
	    RECT 222.2000 151.1000 222.6000 153.0000 ;
	    RECT 223.8000 151.1000 224.2000 153.0000 ;
	    RECT 224.6000 151.1000 225.0000 153.1000 ;
	    RECT 225.4000 151.1000 225.8000 155.8000 ;
	    RECT 227.8000 155.8000 228.2000 155.9000 ;
	    RECT 227.0000 154.8000 227.4000 155.6000 ;
	    RECT 227.8000 154.2000 228.1000 155.8000 ;
	    RECT 229.4000 154.8000 229.9000 155.2000 ;
	    RECT 229.5000 154.4000 229.9000 154.8000 ;
	    RECT 230.4000 154.9000 230.7000 155.9000 ;
	    RECT 230.4000 154.5000 230.9000 154.9000 ;
	    RECT 227.8000 153.8000 228.2000 154.2000 ;
	    RECT 226.2000 152.4000 226.6000 153.2000 ;
	    RECT 227.8000 152.1000 228.1000 153.8000 ;
	    RECT 230.4000 153.7000 230.7000 154.5000 ;
	    RECT 231.2000 154.2000 231.5000 155.9000 ;
	    RECT 233.5000 154.2000 233.8000 155.9000 ;
	    RECT 234.2000 154.8000 234.6000 155.6000 ;
	    RECT 237.0000 155.2000 237.3000 155.9000 ;
	    RECT 239.1000 155.6000 239.4000 155.9000 ;
	    RECT 237.7000 155.3000 239.4000 155.6000 ;
	    RECT 237.7000 155.2000 238.1000 155.3000 ;
	    RECT 236.6000 154.9000 237.3000 155.2000 ;
	    RECT 238.8000 154.9000 239.2000 155.0000 ;
	    RECT 236.6000 154.8000 237.5000 154.9000 ;
	    RECT 237.0000 154.6000 237.5000 154.8000 ;
	    RECT 231.0000 153.8000 231.5000 154.2000 ;
	    RECT 233.4000 153.8000 233.8000 154.2000 ;
	    RECT 235.0000 153.8000 235.8000 154.2000 ;
	    RECT 236.4000 153.8000 236.8000 154.2000 ;
	    RECT 229.4000 153.4000 230.7000 153.7000 ;
	    RECT 228.6000 152.4000 229.0000 153.2000 ;
	    RECT 227.8000 151.1000 228.2000 152.1000 ;
	    RECT 229.4000 151.1000 229.8000 153.4000 ;
	    RECT 231.2000 153.1000 231.5000 153.8000 ;
	    RECT 231.0000 152.8000 231.5000 153.1000 ;
	    RECT 231.0000 151.1000 231.4000 152.8000 ;
	    RECT 232.6000 152.4000 233.0000 153.2000 ;
	    RECT 233.5000 152.1000 233.8000 153.8000 ;
	    RECT 236.5000 153.6000 236.8000 153.8000 ;
	    RECT 235.8000 153.4000 236.2000 153.5000 ;
	    RECT 233.4000 151.1000 233.8000 152.1000 ;
	    RECT 235.0000 153.1000 236.2000 153.4000 ;
	    RECT 236.5000 153.2000 236.9000 153.6000 ;
	    RECT 235.0000 151.1000 235.4000 153.1000 ;
	    RECT 237.2000 152.9000 237.5000 154.6000 ;
	    RECT 237.9000 154.6000 239.2000 154.9000 ;
	    RECT 240.6000 154.8000 241.0000 155.6000 ;
	    RECT 237.9000 154.3000 238.2000 154.6000 ;
	    RECT 237.8000 153.9000 238.2000 154.3000 ;
	    RECT 241.4000 154.2000 241.7000 155.9000 ;
	    RECT 243.0000 154.8000 243.4000 155.6000 ;
	    RECT 243.8000 155.1000 244.1000 155.9000 ;
	    RECT 245.8000 155.2000 246.2000 155.4000 ;
	    RECT 247.8000 155.2000 248.1000 155.9000 ;
	    RECT 249.4000 155.8000 249.8000 155.9000 ;
	    RECT 245.4000 155.1000 246.2000 155.2000 ;
	    RECT 243.8000 154.9000 246.2000 155.1000 ;
	    RECT 247.0000 154.9000 248.2000 155.2000 ;
	    RECT 243.8000 154.8000 245.8000 154.9000 ;
	    RECT 243.8000 154.2000 244.1000 154.8000 ;
	    RECT 239.4000 154.1000 240.2000 154.2000 ;
	    RECT 238.5000 153.8000 240.2000 154.1000 ;
	    RECT 241.4000 153.8000 241.8000 154.2000 ;
	    RECT 243.8000 153.8000 244.2000 154.2000 ;
	    RECT 246.2000 153.8000 246.6000 154.6000 ;
	    RECT 238.5000 153.6000 238.8000 153.8000 ;
	    RECT 237.8000 153.3000 238.8000 153.6000 ;
	    RECT 239.1000 153.4000 239.5000 153.5000 ;
	    RECT 237.8000 153.2000 238.6000 153.3000 ;
	    RECT 239.1000 153.1000 240.2000 153.4000 ;
	    RECT 237.2000 151.1000 238.0000 152.9000 ;
	    RECT 239.8000 151.1000 240.2000 153.1000 ;
	    RECT 241.4000 152.1000 241.7000 153.8000 ;
	    RECT 242.2000 152.4000 242.6000 153.2000 ;
	    RECT 243.8000 152.1000 244.1000 153.8000 ;
	    RECT 244.6000 152.4000 245.0000 153.2000 ;
	    RECT 247.0000 153.1000 247.3000 154.9000 ;
	    RECT 247.8000 154.8000 248.2000 154.9000 ;
	    RECT 249.5000 154.2000 249.8000 155.8000 ;
	    RECT 250.2000 154.8000 250.6000 155.6000 ;
	    RECT 251.1000 155.2000 251.4000 155.9000 ;
	    RECT 253.0000 155.2000 253.4000 155.4000 ;
	    RECT 251.0000 154.9000 252.2000 155.2000 ;
	    RECT 253.0000 154.9000 253.8000 155.2000 ;
	    RECT 251.0000 154.8000 251.4000 154.9000 ;
	    RECT 249.4000 153.8000 249.8000 154.2000 ;
	    RECT 241.4000 151.1000 241.8000 152.1000 ;
	    RECT 243.8000 151.1000 244.2000 152.1000 ;
	    RECT 247.0000 151.1000 247.4000 153.1000 ;
	    RECT 247.8000 152.8000 248.2000 153.2000 ;
	    RECT 247.7000 152.4000 248.1000 152.8000 ;
	    RECT 248.6000 152.4000 249.0000 153.2000 ;
	    RECT 249.5000 152.1000 249.8000 153.8000 ;
	    RECT 251.0000 152.8000 251.4000 153.2000 ;
	    RECT 251.9000 153.1000 252.2000 154.9000 ;
	    RECT 253.4000 154.8000 253.8000 154.9000 ;
	    RECT 252.6000 153.8000 253.0000 154.6000 ;
	    RECT 255.0000 154.4000 255.4000 155.2000 ;
	    RECT 255.7000 154.2000 256.0000 155.9000 ;
	    RECT 256.6000 155.8000 257.0000 155.9000 ;
	    RECT 257.4000 154.8000 257.8000 155.6000 ;
	    RECT 258.2000 154.2000 258.5000 155.9000 ;
	    RECT 260.7000 154.2000 261.0000 155.9000 ;
	    RECT 261.4000 155.1000 261.8000 155.6000 ;
	    RECT 262.2000 155.1000 262.6000 159.9000 ;
	    RECT 263.8000 155.8000 264.2000 156.6000 ;
	    RECT 261.4000 154.8000 262.6000 155.1000 ;
	    RECT 254.2000 154.1000 254.6000 154.2000 ;
	    RECT 254.2000 153.8000 255.0000 154.1000 ;
	    RECT 255.7000 153.8000 257.0000 154.2000 ;
	    RECT 258.2000 154.1000 258.6000 154.2000 ;
	    RECT 258.2000 153.8000 260.1000 154.1000 ;
	    RECT 260.6000 153.8000 261.0000 154.2000 ;
	    RECT 254.6000 153.6000 255.0000 153.8000 ;
	    RECT 254.3000 153.1000 256.1000 153.3000 ;
	    RECT 256.6000 153.1000 256.9000 153.8000 ;
	    RECT 251.1000 152.4000 251.5000 152.8000 ;
	    RECT 249.4000 151.1000 249.8000 152.1000 ;
	    RECT 251.8000 151.1000 252.2000 153.1000 ;
	    RECT 254.2000 153.0000 256.2000 153.1000 ;
	    RECT 254.2000 151.1000 254.6000 153.0000 ;
	    RECT 255.8000 151.1000 256.2000 153.0000 ;
	    RECT 256.6000 151.1000 257.0000 153.1000 ;
	    RECT 258.2000 152.1000 258.5000 153.8000 ;
	    RECT 259.8000 153.2000 260.1000 153.8000 ;
	    RECT 259.0000 152.4000 259.4000 153.2000 ;
	    RECT 259.8000 152.4000 260.2000 153.2000 ;
	    RECT 260.7000 153.1000 261.0000 153.8000 ;
	    RECT 261.4000 153.1000 261.8000 153.2000 ;
	    RECT 260.6000 152.8000 261.8000 153.1000 ;
	    RECT 260.7000 152.1000 261.0000 152.8000 ;
	    RECT 258.2000 151.1000 258.6000 152.1000 ;
	    RECT 260.6000 151.1000 261.0000 152.1000 ;
	    RECT 262.2000 151.1000 262.6000 154.8000 ;
	    RECT 263.0000 153.1000 263.4000 153.2000 ;
	    RECT 264.6000 153.1000 265.0000 159.9000 ;
	    RECT 266.5000 156.2000 266.9000 159.9000 ;
	    RECT 266.2000 155.9000 266.9000 156.2000 ;
	    RECT 266.2000 155.2000 266.5000 155.9000 ;
	    RECT 268.6000 155.6000 269.0000 159.9000 ;
	    RECT 267.0000 155.4000 269.0000 155.6000 ;
	    RECT 266.9000 155.3000 269.0000 155.4000 ;
	    RECT 266.2000 154.8000 266.6000 155.2000 ;
	    RECT 266.9000 155.0000 267.3000 155.3000 ;
	    RECT 265.4000 153.4000 265.8000 154.2000 ;
	    RECT 263.0000 152.8000 265.0000 153.1000 ;
	    RECT 266.2000 153.1000 266.5000 154.8000 ;
	    RECT 266.9000 153.5000 267.2000 155.0000 ;
	    RECT 266.9000 153.2000 268.1000 153.5000 ;
	    RECT 263.0000 152.4000 263.4000 152.8000 ;
	    RECT 264.1000 151.1000 264.5000 152.8000 ;
	    RECT 266.2000 151.1000 266.6000 153.1000 ;
	    RECT 267.8000 152.1000 268.1000 153.2000 ;
	    RECT 268.6000 152.4000 269.0000 153.2000 ;
	    RECT 267.8000 151.1000 268.2000 152.1000 ;
	    RECT 1.4000 148.9000 1.8000 149.9000 ;
	    RECT 0.6000 147.8000 1.0000 148.6000 ;
	    RECT 1.5000 147.2000 1.8000 148.9000 ;
	    RECT 3.0000 148.0000 3.4000 149.9000 ;
	    RECT 4.6000 148.0000 5.0000 149.9000 ;
	    RECT 3.0000 147.9000 5.0000 148.0000 ;
	    RECT 5.4000 147.9000 5.8000 149.9000 ;
	    RECT 6.2000 148.0000 6.6000 149.9000 ;
	    RECT 7.8000 148.0000 8.2000 149.9000 ;
	    RECT 6.2000 147.9000 8.2000 148.0000 ;
	    RECT 8.6000 147.9000 9.0000 149.9000 ;
	    RECT 9.4000 149.6000 11.4000 149.9000 ;
	    RECT 9.4000 147.9000 9.8000 149.6000 ;
	    RECT 10.2000 147.9000 10.6000 149.3000 ;
	    RECT 11.0000 148.0000 11.4000 149.6000 ;
	    RECT 12.6000 148.0000 13.0000 149.9000 ;
	    RECT 11.0000 147.9000 13.0000 148.0000 ;
	    RECT 3.1000 147.7000 4.9000 147.9000 ;
	    RECT 3.4000 147.2000 3.8000 147.4000 ;
	    RECT 5.4000 147.2000 5.7000 147.9000 ;
	    RECT 6.3000 147.7000 8.1000 147.9000 ;
	    RECT 6.6000 147.2000 7.0000 147.4000 ;
	    RECT 8.6000 147.2000 8.9000 147.9000 ;
	    RECT 10.2000 147.2000 10.5000 147.9000 ;
	    RECT 11.1000 147.7000 12.9000 147.9000 ;
	    RECT 12.2000 147.2000 12.6000 147.4000 ;
	    RECT 1.4000 146.8000 1.8000 147.2000 ;
	    RECT 3.0000 147.1000 3.8000 147.2000 ;
	    RECT 1.5000 145.1000 1.8000 146.8000 ;
	    RECT 2.2000 146.9000 3.8000 147.1000 ;
	    RECT 2.2000 146.8000 3.4000 146.9000 ;
	    RECT 4.5000 146.8000 5.8000 147.2000 ;
	    RECT 6.2000 146.9000 7.0000 147.2000 ;
	    RECT 6.2000 146.8000 6.6000 146.9000 ;
	    RECT 7.7000 146.8000 9.0000 147.2000 ;
	    RECT 2.2000 146.2000 2.5000 146.8000 ;
	    RECT 2.2000 145.4000 2.6000 146.2000 ;
	    RECT 3.8000 145.8000 4.2000 146.6000 ;
	    RECT 4.5000 145.1000 4.8000 146.8000 ;
	    RECT 7.7000 146.1000 8.0000 146.8000 ;
	    RECT 9.4000 146.4000 9.8000 147.2000 ;
	    RECT 10.2000 146.9000 11.4000 147.2000 ;
	    RECT 12.2000 147.1000 13.0000 147.2000 ;
	    RECT 14.2000 147.1000 14.6000 149.9000 ;
	    RECT 15.6000 147.1000 16.0000 149.9000 ;
	    RECT 18.5000 148.2000 18.9000 149.9000 ;
	    RECT 18.5000 147.9000 19.4000 148.2000 ;
	    RECT 20.6000 148.0000 21.0000 149.9000 ;
	    RECT 22.2000 148.0000 22.6000 149.9000 ;
	    RECT 20.6000 147.9000 22.6000 148.0000 ;
	    RECT 23.0000 147.9000 23.4000 149.9000 ;
	    RECT 25.4000 147.9000 25.8000 149.9000 ;
	    RECT 26.1000 148.2000 26.5000 148.6000 ;
	    RECT 12.2000 146.9000 14.6000 147.1000 ;
	    RECT 11.0000 146.8000 11.4000 146.9000 ;
	    RECT 12.6000 146.8000 14.6000 146.9000 ;
	    RECT 8.6000 146.1000 9.0000 146.2000 ;
	    RECT 7.7000 145.8000 9.0000 146.1000 ;
	    RECT 5.4000 145.1000 5.8000 145.2000 ;
	    RECT 7.7000 145.1000 8.0000 145.8000 ;
	    RECT 11.1000 145.2000 11.4000 146.8000 ;
	    RECT 8.6000 145.1000 9.0000 145.2000 ;
	    RECT 1.4000 144.7000 2.3000 145.1000 ;
	    RECT 1.9000 142.2000 2.3000 144.7000 ;
	    RECT 1.4000 141.8000 2.3000 142.2000 ;
	    RECT 1.9000 141.1000 2.3000 141.8000 ;
	    RECT 4.3000 144.8000 4.8000 145.1000 ;
	    RECT 5.1000 144.8000 5.8000 145.1000 ;
	    RECT 7.5000 144.8000 8.0000 145.1000 ;
	    RECT 8.3000 144.8000 9.0000 145.1000 ;
	    RECT 10.2000 145.1000 11.4000 145.2000 ;
	    RECT 13.4000 145.1000 13.8000 145.2000 ;
	    RECT 14.2000 145.1000 14.6000 146.8000 ;
	    RECT 15.1000 146.9000 16.0000 147.1000 ;
	    RECT 15.1000 146.8000 15.9000 146.9000 ;
	    RECT 15.1000 145.2000 15.4000 146.8000 ;
	    RECT 16.2000 145.8000 17.0000 146.2000 ;
	    RECT 19.0000 146.1000 19.4000 147.9000 ;
	    RECT 20.7000 147.7000 22.5000 147.9000 ;
	    RECT 21.0000 147.2000 21.4000 147.4000 ;
	    RECT 23.0000 147.2000 23.3000 147.9000 ;
	    RECT 20.6000 146.9000 21.4000 147.2000 ;
	    RECT 20.6000 146.8000 21.0000 146.9000 ;
	    RECT 22.1000 146.8000 23.4000 147.2000 ;
	    RECT 17.4000 145.8000 19.4000 146.1000 ;
	    RECT 21.4000 145.8000 21.8000 146.6000 ;
	    RECT 10.2000 144.8000 11.7000 145.1000 ;
	    RECT 13.4000 144.8000 14.6000 145.1000 ;
	    RECT 15.0000 144.8000 15.4000 145.2000 ;
	    RECT 17.4000 144.8000 17.8000 145.8000 ;
	    RECT 4.3000 141.1000 4.7000 144.8000 ;
	    RECT 5.1000 144.2000 5.4000 144.8000 ;
	    RECT 5.0000 143.8000 5.4000 144.2000 ;
	    RECT 7.5000 141.1000 7.9000 144.8000 ;
	    RECT 8.3000 144.2000 8.6000 144.8000 ;
	    RECT 8.2000 143.8000 8.6000 144.2000 ;
	    RECT 10.7000 141.1000 11.7000 144.8000 ;
	    RECT 14.2000 141.1000 14.6000 144.8000 ;
	    RECT 15.1000 143.5000 15.4000 144.8000 ;
	    RECT 15.8000 143.8000 16.2000 144.6000 ;
	    RECT 18.2000 144.4000 18.6000 145.2000 ;
	    RECT 15.1000 143.2000 16.9000 143.5000 ;
	    RECT 15.1000 143.1000 15.4000 143.2000 ;
	    RECT 15.0000 141.1000 15.4000 143.1000 ;
	    RECT 16.6000 143.1000 16.9000 143.2000 ;
	    RECT 16.6000 141.1000 17.0000 143.1000 ;
	    RECT 19.0000 141.1000 19.4000 145.8000 ;
	    RECT 22.1000 145.1000 22.4000 146.8000 ;
	    RECT 23.0000 146.2000 23.3000 146.8000 ;
	    RECT 24.6000 146.4000 25.0000 147.2000 ;
	    RECT 23.0000 145.8000 23.4000 146.2000 ;
	    RECT 23.8000 146.1000 24.2000 146.2000 ;
	    RECT 25.4000 146.1000 25.7000 147.9000 ;
	    RECT 26.2000 147.8000 26.6000 148.2000 ;
	    RECT 28.6000 147.9000 29.0000 149.9000 ;
	    RECT 29.3000 148.2000 29.7000 148.6000 ;
	    RECT 27.8000 146.4000 28.2000 147.2000 ;
	    RECT 26.2000 146.1000 26.6000 146.2000 ;
	    RECT 23.8000 145.8000 24.6000 146.1000 ;
	    RECT 25.4000 145.8000 26.6000 146.1000 ;
	    RECT 27.0000 146.1000 27.4000 146.2000 ;
	    RECT 28.6000 146.1000 28.9000 147.9000 ;
	    RECT 29.4000 147.8000 29.8000 148.2000 ;
	    RECT 30.2000 147.5000 30.6000 149.9000 ;
	    RECT 32.4000 149.2000 32.8000 149.9000 ;
	    RECT 31.8000 148.9000 32.8000 149.2000 ;
	    RECT 34.6000 148.9000 35.0000 149.9000 ;
	    RECT 36.7000 149.2000 37.3000 149.9000 ;
	    RECT 36.6000 148.9000 37.3000 149.2000 ;
	    RECT 31.8000 148.5000 32.2000 148.9000 ;
	    RECT 34.6000 148.6000 34.9000 148.9000 ;
	    RECT 32.6000 148.2000 33.0000 148.6000 ;
	    RECT 33.5000 148.3000 34.9000 148.6000 ;
	    RECT 36.6000 148.5000 37.0000 148.9000 ;
	    RECT 33.5000 148.2000 33.9000 148.3000 ;
	    RECT 30.6000 147.1000 31.4000 147.2000 ;
	    RECT 32.7000 147.1000 33.0000 148.2000 ;
	    RECT 39.0000 148.1000 39.4000 149.9000 ;
	    RECT 39.8000 148.1000 40.2000 148.6000 ;
	    RECT 39.0000 147.8000 40.2000 148.1000 ;
	    RECT 37.5000 147.7000 37.9000 147.8000 ;
	    RECT 39.0000 147.7000 39.4000 147.8000 ;
	    RECT 37.5000 147.4000 39.4000 147.7000 ;
	    RECT 35.5000 147.1000 35.9000 147.2000 ;
	    RECT 30.6000 146.8000 36.1000 147.1000 ;
	    RECT 32.1000 146.7000 32.5000 146.8000 ;
	    RECT 31.3000 146.2000 31.7000 146.3000 ;
	    RECT 32.6000 146.2000 33.0000 146.3000 ;
	    RECT 35.8000 146.2000 36.1000 146.8000 ;
	    RECT 36.6000 146.4000 37.0000 146.5000 ;
	    RECT 29.4000 146.1000 29.8000 146.2000 ;
	    RECT 27.0000 145.8000 27.8000 146.1000 ;
	    RECT 28.6000 145.8000 29.8000 146.1000 ;
	    RECT 31.3000 145.9000 33.8000 146.2000 ;
	    RECT 33.4000 145.8000 33.8000 145.9000 ;
	    RECT 35.8000 145.8000 36.2000 146.2000 ;
	    RECT 36.6000 146.1000 38.5000 146.4000 ;
	    RECT 38.1000 146.0000 38.5000 146.1000 ;
	    RECT 24.2000 145.6000 24.6000 145.8000 ;
	    RECT 23.0000 145.1000 23.4000 145.2000 ;
	    RECT 26.2000 145.1000 26.5000 145.8000 ;
	    RECT 27.4000 145.6000 27.8000 145.8000 ;
	    RECT 29.4000 145.1000 29.7000 145.8000 ;
	    RECT 30.2000 145.5000 33.0000 145.6000 ;
	    RECT 30.2000 145.4000 33.1000 145.5000 ;
	    RECT 30.2000 145.3000 35.1000 145.4000 ;
	    RECT 21.9000 144.8000 22.4000 145.1000 ;
	    RECT 22.7000 144.8000 23.4000 145.1000 ;
	    RECT 23.8000 144.8000 25.8000 145.1000 ;
	    RECT 21.9000 141.1000 22.3000 144.8000 ;
	    RECT 22.7000 144.2000 23.0000 144.8000 ;
	    RECT 22.6000 143.8000 23.0000 144.2000 ;
	    RECT 23.8000 141.1000 24.2000 144.8000 ;
	    RECT 25.4000 141.1000 25.8000 144.8000 ;
	    RECT 26.2000 141.1000 26.6000 145.1000 ;
	    RECT 27.0000 144.8000 29.0000 145.1000 ;
	    RECT 27.0000 141.1000 27.4000 144.8000 ;
	    RECT 28.6000 141.1000 29.0000 144.8000 ;
	    RECT 29.4000 141.1000 29.8000 145.1000 ;
	    RECT 30.2000 141.1000 30.6000 145.3000 ;
	    RECT 32.7000 145.1000 35.1000 145.3000 ;
	    RECT 31.8000 144.5000 34.5000 144.8000 ;
	    RECT 31.8000 144.4000 32.2000 144.5000 ;
	    RECT 34.1000 144.4000 34.5000 144.5000 ;
	    RECT 34.8000 144.5000 35.1000 145.1000 ;
	    RECT 35.8000 145.2000 36.1000 145.8000 ;
	    RECT 37.3000 145.7000 37.7000 145.8000 ;
	    RECT 39.0000 145.7000 39.4000 147.4000 ;
	    RECT 37.3000 145.4000 39.4000 145.7000 ;
	    RECT 35.8000 144.9000 37.0000 145.2000 ;
	    RECT 35.5000 144.5000 35.9000 144.6000 ;
	    RECT 34.8000 144.2000 35.9000 144.5000 ;
	    RECT 36.7000 144.4000 37.0000 144.9000 ;
	    RECT 36.7000 144.0000 37.4000 144.4000 ;
	    RECT 33.5000 143.7000 33.9000 143.8000 ;
	    RECT 34.9000 143.7000 35.3000 143.8000 ;
	    RECT 31.8000 143.1000 32.2000 143.5000 ;
	    RECT 33.5000 143.4000 35.3000 143.7000 ;
	    RECT 34.6000 143.1000 34.9000 143.4000 ;
	    RECT 36.6000 143.1000 37.0000 143.5000 ;
	    RECT 31.8000 142.8000 32.8000 143.1000 ;
	    RECT 32.4000 141.1000 32.8000 142.8000 ;
	    RECT 34.6000 141.1000 35.0000 143.1000 ;
	    RECT 36.7000 141.1000 37.3000 143.1000 ;
	    RECT 39.0000 141.1000 39.4000 145.4000 ;
	    RECT 40.6000 147.1000 41.0000 149.9000 ;
	    RECT 41.4000 148.0000 41.8000 149.9000 ;
	    RECT 43.0000 149.6000 45.0000 149.9000 ;
	    RECT 43.0000 148.0000 43.4000 149.6000 ;
	    RECT 41.4000 147.9000 43.4000 148.0000 ;
	    RECT 41.5000 147.7000 43.3000 147.9000 ;
	    RECT 43.8000 147.8000 44.2000 149.3000 ;
	    RECT 44.6000 147.9000 45.0000 149.6000 ;
	    RECT 41.8000 147.2000 42.2000 147.4000 ;
	    RECT 43.9000 147.2000 44.2000 147.8000 ;
	    RECT 41.4000 147.1000 42.2000 147.2000 ;
	    RECT 40.6000 146.9000 42.2000 147.1000 ;
	    RECT 43.0000 146.9000 44.2000 147.2000 ;
	    RECT 44.6000 147.1000 45.0000 147.2000 ;
	    RECT 45.4000 147.1000 45.8000 149.9000 ;
	    RECT 49.4000 148.9000 49.8000 149.9000 ;
	    RECT 51.0000 149.2000 51.4000 149.9000 ;
	    RECT 49.2000 148.8000 49.8000 148.9000 ;
	    RECT 50.9000 148.8000 51.4000 149.2000 ;
	    RECT 46.2000 147.8000 46.6000 148.6000 ;
	    RECT 49.2000 148.5000 51.2000 148.8000 ;
	    RECT 40.6000 146.8000 41.8000 146.9000 ;
	    RECT 43.0000 146.8000 43.4000 146.9000 ;
	    RECT 44.6000 146.8000 45.8000 147.1000 ;
	    RECT 40.6000 141.1000 41.0000 146.8000 ;
	    RECT 42.2000 145.8000 42.6000 146.6000 ;
	    RECT 43.0000 145.1000 43.3000 146.8000 ;
	    RECT 43.8000 145.8000 44.2000 146.6000 ;
	    RECT 44.6000 146.4000 45.0000 146.8000 ;
	    RECT 42.7000 141.1000 43.7000 145.1000 ;
	    RECT 45.4000 141.1000 45.8000 146.8000 ;
	    RECT 49.2000 145.2000 49.5000 148.5000 ;
	    RECT 51.0000 147.8000 52.2000 148.2000 ;
	    RECT 53.4000 147.9000 53.8000 149.9000 ;
	    RECT 54.2000 148.0000 54.6000 149.9000 ;
	    RECT 55.8000 148.0000 56.2000 149.9000 ;
	    RECT 54.2000 147.9000 56.2000 148.0000 ;
	    RECT 53.5000 147.2000 53.8000 147.9000 ;
	    RECT 54.3000 147.7000 56.1000 147.9000 ;
	    RECT 55.4000 147.2000 55.8000 147.4000 ;
	    RECT 50.6000 147.1000 51.4000 147.2000 ;
	    RECT 53.4000 147.1000 54.7000 147.2000 ;
	    RECT 50.6000 146.8000 54.7000 147.1000 ;
	    RECT 55.4000 147.1000 56.2000 147.2000 ;
	    RECT 56.6000 147.1000 57.0000 149.9000 ;
	    RECT 57.4000 147.8000 57.8000 148.6000 ;
	    RECT 55.4000 146.9000 57.0000 147.1000 ;
	    RECT 55.8000 146.8000 57.0000 146.9000 ;
	    RECT 49.8000 145.8000 50.6000 146.2000 ;
	    RECT 47.8000 144.9000 49.5000 145.2000 ;
	    RECT 53.4000 145.1000 53.8000 145.2000 ;
	    RECT 54.4000 145.1000 54.7000 146.8000 ;
	    RECT 55.0000 145.8000 55.4000 146.6000 ;
	    RECT 47.8000 144.8000 48.2000 144.9000 ;
	    RECT 53.4000 144.8000 54.1000 145.1000 ;
	    RECT 54.4000 144.8000 54.9000 145.1000 ;
	    RECT 47.9000 144.5000 48.2000 144.8000 ;
	    RECT 48.7000 144.5000 50.5000 144.6000 ;
	    RECT 47.0000 141.5000 47.4000 144.5000 ;
	    RECT 47.8000 141.7000 48.2000 144.5000 ;
	    RECT 48.6000 144.3000 50.5000 144.5000 ;
	    RECT 47.1000 141.4000 47.4000 141.5000 ;
	    RECT 48.6000 141.5000 49.0000 144.3000 ;
	    RECT 50.2000 144.1000 50.5000 144.3000 ;
	    RECT 51.1000 144.4000 52.9000 144.7000 ;
	    RECT 51.1000 144.1000 51.4000 144.4000 ;
	    RECT 48.6000 141.4000 48.9000 141.5000 ;
	    RECT 47.1000 141.1000 48.9000 141.4000 ;
	    RECT 49.4000 141.4000 49.8000 144.0000 ;
	    RECT 50.2000 141.7000 50.6000 144.1000 ;
	    RECT 51.0000 141.4000 51.4000 144.1000 ;
	    RECT 49.4000 141.1000 51.4000 141.4000 ;
	    RECT 52.6000 144.1000 52.9000 144.4000 ;
	    RECT 53.8000 144.2000 54.1000 144.8000 ;
	    RECT 52.6000 141.1000 53.0000 144.1000 ;
	    RECT 53.8000 143.8000 54.2000 144.2000 ;
	    RECT 54.5000 141.1000 54.9000 144.8000 ;
	    RECT 56.6000 141.1000 57.0000 146.8000 ;
	    RECT 59.8000 146.1000 60.2000 149.9000 ;
	    RECT 60.6000 147.8000 61.0000 148.6000 ;
	    RECT 63.0000 147.9000 63.4000 149.9000 ;
	    RECT 63.7000 148.2000 64.1000 148.6000 ;
	    RECT 61.4000 147.1000 61.8000 147.2000 ;
	    RECT 62.2000 147.1000 62.6000 147.2000 ;
	    RECT 61.4000 146.8000 62.6000 147.1000 ;
	    RECT 62.2000 146.4000 62.6000 146.8000 ;
	    RECT 61.4000 146.1000 61.8000 146.2000 ;
	    RECT 63.0000 146.1000 63.3000 147.9000 ;
	    RECT 63.8000 147.8000 64.2000 148.2000 ;
	    RECT 64.6000 147.5000 65.0000 149.9000 ;
	    RECT 66.8000 149.2000 67.2000 149.9000 ;
	    RECT 66.2000 148.9000 67.2000 149.2000 ;
	    RECT 69.0000 148.9000 69.4000 149.9000 ;
	    RECT 71.1000 149.2000 71.7000 149.9000 ;
	    RECT 71.0000 148.9000 71.7000 149.2000 ;
	    RECT 66.2000 148.5000 66.6000 148.9000 ;
	    RECT 69.0000 148.6000 69.3000 148.9000 ;
	    RECT 67.0000 148.2000 67.4000 148.6000 ;
	    RECT 67.9000 148.3000 69.3000 148.6000 ;
	    RECT 71.0000 148.5000 71.4000 148.9000 ;
	    RECT 67.9000 148.2000 68.3000 148.3000 ;
	    RECT 65.0000 147.1000 65.8000 147.2000 ;
	    RECT 67.1000 147.1000 67.4000 148.2000 ;
	    RECT 71.9000 147.7000 72.3000 147.8000 ;
	    RECT 73.4000 147.7000 73.8000 149.9000 ;
	    RECT 71.9000 147.4000 73.8000 147.7000 ;
	    RECT 69.9000 147.1000 70.3000 147.2000 ;
	    RECT 65.0000 146.8000 70.5000 147.1000 ;
	    RECT 66.5000 146.7000 66.9000 146.8000 ;
	    RECT 65.7000 146.2000 66.1000 146.3000 ;
	    RECT 70.2000 146.2000 70.5000 146.8000 ;
	    RECT 71.0000 146.4000 71.4000 146.5000 ;
	    RECT 63.8000 146.1000 64.2000 146.2000 ;
	    RECT 59.8000 145.8000 62.2000 146.1000 ;
	    RECT 63.0000 145.8000 64.2000 146.1000 ;
	    RECT 65.7000 145.9000 68.2000 146.2000 ;
	    RECT 67.8000 145.8000 68.2000 145.9000 ;
	    RECT 70.2000 145.8000 70.6000 146.2000 ;
	    RECT 71.0000 146.1000 72.9000 146.4000 ;
	    RECT 72.5000 146.0000 72.9000 146.1000 ;
	    RECT 59.8000 141.1000 60.2000 145.8000 ;
	    RECT 61.8000 145.6000 62.2000 145.8000 ;
	    RECT 63.8000 145.1000 64.1000 145.8000 ;
	    RECT 64.6000 145.5000 67.4000 145.6000 ;
	    RECT 64.6000 145.4000 67.5000 145.5000 ;
	    RECT 64.6000 145.3000 69.5000 145.4000 ;
	    RECT 61.4000 144.8000 63.4000 145.1000 ;
	    RECT 61.4000 141.1000 61.8000 144.8000 ;
	    RECT 63.0000 141.1000 63.4000 144.8000 ;
	    RECT 63.8000 141.1000 64.2000 145.1000 ;
	    RECT 64.6000 141.1000 65.0000 145.3000 ;
	    RECT 67.1000 145.1000 69.5000 145.3000 ;
	    RECT 66.2000 144.5000 68.9000 144.8000 ;
	    RECT 66.2000 144.4000 66.6000 144.5000 ;
	    RECT 68.5000 144.4000 68.9000 144.5000 ;
	    RECT 69.2000 144.5000 69.5000 145.1000 ;
	    RECT 70.2000 145.2000 70.5000 145.8000 ;
	    RECT 71.7000 145.7000 72.1000 145.8000 ;
	    RECT 73.4000 145.7000 73.8000 147.4000 ;
	    RECT 71.7000 145.4000 73.8000 145.7000 ;
	    RECT 70.2000 144.9000 71.4000 145.2000 ;
	    RECT 69.9000 144.5000 70.3000 144.6000 ;
	    RECT 69.2000 144.2000 70.3000 144.5000 ;
	    RECT 71.1000 144.4000 71.4000 144.9000 ;
	    RECT 71.1000 144.0000 71.8000 144.4000 ;
	    RECT 67.9000 143.7000 68.3000 143.8000 ;
	    RECT 69.3000 143.7000 69.7000 143.8000 ;
	    RECT 66.2000 143.1000 66.6000 143.5000 ;
	    RECT 67.9000 143.4000 69.7000 143.7000 ;
	    RECT 69.0000 143.1000 69.3000 143.4000 ;
	    RECT 71.0000 143.1000 71.4000 143.5000 ;
	    RECT 66.2000 142.8000 67.2000 143.1000 ;
	    RECT 66.8000 141.1000 67.2000 142.8000 ;
	    RECT 69.0000 141.1000 69.4000 143.1000 ;
	    RECT 71.1000 141.1000 71.7000 143.1000 ;
	    RECT 73.4000 141.1000 73.8000 145.4000 ;
	    RECT 74.2000 147.7000 74.6000 149.9000 ;
	    RECT 76.3000 149.2000 76.9000 149.9000 ;
	    RECT 76.3000 148.9000 77.0000 149.2000 ;
	    RECT 78.6000 148.9000 79.0000 149.9000 ;
	    RECT 80.8000 149.2000 81.2000 149.9000 ;
	    RECT 80.8000 148.9000 81.8000 149.2000 ;
	    RECT 76.6000 148.5000 77.0000 148.9000 ;
	    RECT 78.7000 148.6000 79.0000 148.9000 ;
	    RECT 78.7000 148.3000 80.1000 148.6000 ;
	    RECT 79.7000 148.2000 80.1000 148.3000 ;
	    RECT 80.6000 148.2000 81.0000 148.6000 ;
	    RECT 81.4000 148.5000 81.8000 148.9000 ;
	    RECT 75.7000 147.7000 76.1000 147.8000 ;
	    RECT 74.2000 147.4000 76.1000 147.7000 ;
	    RECT 74.2000 145.7000 74.6000 147.4000 ;
	    RECT 77.7000 147.1000 78.1000 147.2000 ;
	    RECT 80.6000 147.1000 80.9000 148.2000 ;
	    RECT 83.0000 147.5000 83.4000 149.9000 ;
	    RECT 84.1000 149.2000 84.5000 149.9000 ;
	    RECT 84.1000 148.8000 85.0000 149.2000 ;
	    RECT 84.1000 148.2000 84.5000 148.8000 ;
	    RECT 84.1000 147.9000 85.0000 148.2000 ;
	    RECT 82.2000 147.1000 83.0000 147.2000 ;
	    RECT 77.5000 146.8000 83.0000 147.1000 ;
	    RECT 76.6000 146.4000 77.0000 146.5000 ;
	    RECT 75.1000 146.1000 77.0000 146.4000 ;
	    RECT 77.5000 146.2000 77.8000 146.8000 ;
	    RECT 81.1000 146.7000 81.5000 146.8000 ;
	    RECT 81.9000 146.2000 82.3000 146.3000 ;
	    RECT 75.1000 146.0000 75.5000 146.1000 ;
	    RECT 77.4000 145.8000 77.8000 146.2000 ;
	    RECT 79.8000 145.9000 82.3000 146.2000 ;
	    RECT 79.8000 145.8000 80.2000 145.9000 ;
	    RECT 75.9000 145.7000 76.3000 145.8000 ;
	    RECT 74.2000 145.4000 76.3000 145.7000 ;
	    RECT 74.2000 141.1000 74.6000 145.4000 ;
	    RECT 77.5000 145.2000 77.8000 145.8000 ;
	    RECT 80.6000 145.5000 83.4000 145.6000 ;
	    RECT 80.5000 145.4000 83.4000 145.5000 ;
	    RECT 76.6000 144.9000 77.8000 145.2000 ;
	    RECT 78.5000 145.3000 83.4000 145.4000 ;
	    RECT 78.5000 145.1000 80.9000 145.3000 ;
	    RECT 76.6000 144.4000 76.9000 144.9000 ;
	    RECT 76.2000 144.0000 76.9000 144.4000 ;
	    RECT 77.7000 144.5000 78.1000 144.6000 ;
	    RECT 78.5000 144.5000 78.8000 145.1000 ;
	    RECT 77.7000 144.2000 78.8000 144.5000 ;
	    RECT 79.1000 144.5000 81.8000 144.8000 ;
	    RECT 79.1000 144.4000 79.5000 144.5000 ;
	    RECT 81.4000 144.4000 81.8000 144.5000 ;
	    RECT 78.3000 143.7000 78.7000 143.8000 ;
	    RECT 79.7000 143.7000 80.1000 143.8000 ;
	    RECT 76.6000 143.1000 77.0000 143.5000 ;
	    RECT 78.3000 143.4000 80.1000 143.7000 ;
	    RECT 78.7000 143.1000 79.0000 143.4000 ;
	    RECT 81.4000 143.1000 81.8000 143.5000 ;
	    RECT 76.3000 141.1000 76.9000 143.1000 ;
	    RECT 78.6000 141.1000 79.0000 143.1000 ;
	    RECT 80.8000 142.8000 81.8000 143.1000 ;
	    RECT 80.8000 141.1000 81.2000 142.8000 ;
	    RECT 83.0000 141.1000 83.4000 145.3000 ;
	    RECT 83.8000 143.8000 84.2000 145.2000 ;
	    RECT 84.6000 141.1000 85.0000 147.9000 ;
	    RECT 85.4000 146.8000 85.8000 147.6000 ;
	    RECT 86.2000 147.5000 86.6000 149.9000 ;
	    RECT 88.4000 149.2000 88.8000 149.9000 ;
	    RECT 87.8000 148.9000 88.8000 149.2000 ;
	    RECT 90.6000 148.9000 91.0000 149.9000 ;
	    RECT 92.7000 149.2000 93.3000 149.9000 ;
	    RECT 92.6000 148.9000 93.3000 149.2000 ;
	    RECT 87.8000 148.5000 88.2000 148.9000 ;
	    RECT 90.6000 148.6000 90.9000 148.9000 ;
	    RECT 88.6000 148.2000 89.0000 148.6000 ;
	    RECT 89.5000 148.3000 90.9000 148.6000 ;
	    RECT 92.6000 148.5000 93.0000 148.9000 ;
	    RECT 89.5000 148.2000 89.9000 148.3000 ;
	    RECT 86.6000 147.1000 87.4000 147.2000 ;
	    RECT 88.7000 147.1000 89.0000 148.2000 ;
	    RECT 93.5000 147.7000 93.9000 147.8000 ;
	    RECT 95.0000 147.7000 95.4000 149.9000 ;
	    RECT 96.6000 148.9000 97.0000 149.9000 ;
	    RECT 95.8000 147.8000 96.2000 148.6000 ;
	    RECT 93.5000 147.4000 95.4000 147.7000 ;
	    RECT 91.5000 147.1000 91.9000 147.2000 ;
	    RECT 86.6000 146.8000 92.1000 147.1000 ;
	    RECT 88.1000 146.7000 88.5000 146.8000 ;
	    RECT 87.3000 146.2000 87.7000 146.3000 ;
	    RECT 91.8000 146.2000 92.1000 146.8000 ;
	    RECT 92.6000 146.4000 93.0000 146.5000 ;
	    RECT 87.3000 145.9000 89.8000 146.2000 ;
	    RECT 89.4000 145.8000 89.8000 145.9000 ;
	    RECT 91.8000 145.8000 92.2000 146.2000 ;
	    RECT 92.6000 146.1000 94.5000 146.4000 ;
	    RECT 94.1000 146.0000 94.5000 146.1000 ;
	    RECT 86.2000 145.5000 89.0000 145.6000 ;
	    RECT 86.2000 145.4000 89.1000 145.5000 ;
	    RECT 86.2000 145.3000 91.1000 145.4000 ;
	    RECT 86.2000 141.1000 86.6000 145.3000 ;
	    RECT 88.7000 145.1000 91.1000 145.3000 ;
	    RECT 87.8000 144.5000 90.5000 144.8000 ;
	    RECT 87.8000 144.4000 88.2000 144.5000 ;
	    RECT 90.1000 144.4000 90.5000 144.5000 ;
	    RECT 90.8000 144.5000 91.1000 145.1000 ;
	    RECT 91.8000 145.2000 92.1000 145.8000 ;
	    RECT 93.3000 145.7000 93.7000 145.8000 ;
	    RECT 95.0000 145.7000 95.4000 147.4000 ;
	    RECT 96.7000 147.2000 97.0000 148.9000 ;
	    RECT 98.2000 147.9000 98.6000 149.9000 ;
	    RECT 99.0000 148.0000 99.4000 149.9000 ;
	    RECT 100.6000 148.0000 101.0000 149.9000 ;
	    RECT 99.0000 147.9000 101.0000 148.0000 ;
	    RECT 98.3000 147.2000 98.6000 147.9000 ;
	    RECT 99.1000 147.7000 100.9000 147.9000 ;
	    RECT 100.2000 147.2000 100.6000 147.4000 ;
	    RECT 95.8000 146.8000 96.2000 147.2000 ;
	    RECT 96.6000 146.8000 97.0000 147.2000 ;
	    RECT 98.2000 146.8000 99.5000 147.2000 ;
	    RECT 100.2000 147.1000 101.0000 147.2000 ;
	    RECT 101.4000 147.1000 101.8000 149.9000 ;
	    RECT 102.2000 147.8000 102.6000 148.6000 ;
	    RECT 104.8000 148.2000 105.2000 149.9000 ;
	    RECT 106.5000 148.2000 106.9000 149.9000 ;
	    RECT 111.0000 148.9000 111.4000 149.9000 ;
	    RECT 113.4000 148.9000 113.8000 149.9000 ;
	    RECT 104.8000 147.8000 105.8000 148.2000 ;
	    RECT 106.5000 147.9000 107.4000 148.2000 ;
	    RECT 100.2000 146.9000 101.8000 147.1000 ;
	    RECT 104.8000 147.1000 105.2000 147.8000 ;
	    RECT 104.8000 146.9000 105.7000 147.1000 ;
	    RECT 100.6000 146.8000 101.8000 146.9000 ;
	    RECT 104.9000 146.8000 105.7000 146.9000 ;
	    RECT 95.8000 146.1000 96.1000 146.8000 ;
	    RECT 96.7000 146.1000 97.0000 146.8000 ;
	    RECT 95.8000 145.8000 97.0000 146.1000 ;
	    RECT 93.3000 145.4000 95.4000 145.7000 ;
	    RECT 91.8000 144.9000 93.0000 145.2000 ;
	    RECT 91.5000 144.5000 91.9000 144.6000 ;
	    RECT 90.8000 144.2000 91.9000 144.5000 ;
	    RECT 92.7000 144.4000 93.0000 144.9000 ;
	    RECT 92.7000 144.0000 93.4000 144.4000 ;
	    RECT 89.5000 143.7000 89.9000 143.8000 ;
	    RECT 90.9000 143.7000 91.3000 143.8000 ;
	    RECT 87.8000 143.1000 88.2000 143.5000 ;
	    RECT 89.5000 143.4000 91.3000 143.7000 ;
	    RECT 90.6000 143.1000 90.9000 143.4000 ;
	    RECT 92.6000 143.1000 93.0000 143.5000 ;
	    RECT 87.8000 142.8000 88.8000 143.1000 ;
	    RECT 88.4000 141.1000 88.8000 142.8000 ;
	    RECT 90.6000 141.1000 91.0000 143.1000 ;
	    RECT 92.7000 141.1000 93.3000 143.1000 ;
	    RECT 95.0000 141.1000 95.4000 145.4000 ;
	    RECT 96.7000 145.1000 97.0000 145.8000 ;
	    RECT 97.4000 146.1000 97.8000 146.2000 ;
	    RECT 99.2000 146.1000 99.5000 146.8000 ;
	    RECT 97.4000 145.8000 99.5000 146.1000 ;
	    RECT 99.8000 145.8000 100.2000 146.6000 ;
	    RECT 97.4000 145.4000 97.8000 145.8000 ;
	    RECT 98.2000 145.1000 98.6000 145.2000 ;
	    RECT 99.2000 145.1000 99.5000 145.8000 ;
	    RECT 96.6000 144.7000 97.5000 145.1000 ;
	    RECT 98.2000 144.8000 98.9000 145.1000 ;
	    RECT 99.2000 144.8000 99.7000 145.1000 ;
	    RECT 97.1000 141.1000 97.5000 144.7000 ;
	    RECT 98.6000 144.2000 98.9000 144.8000 ;
	    RECT 98.6000 143.8000 99.0000 144.2000 ;
	    RECT 99.3000 141.1000 99.7000 144.8000 ;
	    RECT 101.4000 141.1000 101.8000 146.8000 ;
	    RECT 103.8000 145.8000 104.6000 146.2000 ;
	    RECT 103.0000 144.8000 103.4000 145.6000 ;
	    RECT 105.4000 145.2000 105.7000 146.8000 ;
	    RECT 107.0000 146.1000 107.4000 147.9000 ;
	    RECT 110.2000 147.8000 110.6000 148.6000 ;
	    RECT 107.8000 147.1000 108.2000 147.6000 ;
	    RECT 111.1000 147.2000 111.4000 148.9000 ;
	    RECT 111.8000 148.1000 112.2000 148.2000 ;
	    RECT 112.6000 148.1000 113.0000 148.6000 ;
	    RECT 111.8000 147.8000 113.0000 148.1000 ;
	    RECT 113.5000 147.2000 113.8000 148.9000 ;
	    RECT 116.3000 148.2000 116.7000 149.9000 ;
	    RECT 115.8000 147.9000 116.7000 148.2000 ;
	    RECT 109.4000 147.1000 109.8000 147.2000 ;
	    RECT 107.8000 146.8000 109.8000 147.1000 ;
	    RECT 111.0000 147.1000 111.4000 147.2000 ;
	    RECT 112.6000 147.1000 113.0000 147.2000 ;
	    RECT 111.0000 146.8000 113.0000 147.1000 ;
	    RECT 113.4000 146.8000 113.8000 147.2000 ;
	    RECT 115.0000 146.8000 115.4000 147.6000 ;
	    RECT 107.8000 146.1000 108.2000 146.2000 ;
	    RECT 107.0000 145.8000 108.2000 146.1000 ;
	    RECT 105.4000 144.8000 105.8000 145.2000 ;
	    RECT 102.2000 144.1000 102.6000 144.2000 ;
	    RECT 104.6000 144.1000 105.0000 144.6000 ;
	    RECT 102.2000 143.8000 105.0000 144.1000 ;
	    RECT 105.4000 143.5000 105.7000 144.8000 ;
	    RECT 106.2000 144.4000 106.6000 145.2000 ;
	    RECT 103.9000 143.2000 105.7000 143.5000 ;
	    RECT 103.9000 143.1000 104.2000 143.2000 ;
	    RECT 103.8000 141.1000 104.2000 143.1000 ;
	    RECT 105.4000 143.1000 105.7000 143.2000 ;
	    RECT 105.4000 141.1000 105.8000 143.1000 ;
	    RECT 107.0000 141.1000 107.4000 145.8000 ;
	    RECT 111.1000 145.1000 111.4000 146.8000 ;
	    RECT 111.8000 145.4000 112.2000 146.2000 ;
	    RECT 113.5000 145.1000 113.8000 146.8000 ;
	    RECT 114.2000 146.1000 114.6000 146.2000 ;
	    RECT 115.8000 146.1000 116.2000 147.9000 ;
	    RECT 119.2000 147.1000 119.6000 149.9000 ;
	    RECT 119.2000 146.9000 120.1000 147.1000 ;
	    RECT 119.3000 146.8000 120.1000 146.9000 ;
	    RECT 114.2000 145.8000 116.2000 146.1000 ;
	    RECT 118.2000 145.8000 119.0000 146.2000 ;
	    RECT 114.2000 145.4000 114.6000 145.8000 ;
	    RECT 111.0000 144.7000 111.9000 145.1000 ;
	    RECT 113.4000 144.7000 114.3000 145.1000 ;
	    RECT 111.5000 141.1000 111.9000 144.7000 ;
	    RECT 113.9000 142.2000 114.3000 144.7000 ;
	    RECT 113.4000 141.8000 114.3000 142.2000 ;
	    RECT 113.9000 141.1000 114.3000 141.8000 ;
	    RECT 115.8000 141.1000 116.2000 145.8000 ;
	    RECT 116.6000 144.1000 117.0000 145.2000 ;
	    RECT 117.4000 144.8000 117.8000 145.6000 ;
	    RECT 119.8000 145.2000 120.1000 146.8000 ;
	    RECT 119.8000 144.8000 120.2000 145.2000 ;
	    RECT 118.2000 144.1000 118.6000 144.2000 ;
	    RECT 116.6000 143.8000 118.6000 144.1000 ;
	    RECT 119.0000 143.8000 119.4000 144.6000 ;
	    RECT 119.8000 143.5000 120.1000 144.8000 ;
	    RECT 118.3000 143.2000 120.1000 143.5000 ;
	    RECT 118.3000 143.1000 118.6000 143.2000 ;
	    RECT 118.2000 141.1000 118.6000 143.1000 ;
	    RECT 119.8000 143.1000 120.1000 143.2000 ;
	    RECT 119.8000 141.1000 120.2000 143.1000 ;
	    RECT 120.6000 141.1000 121.0000 149.9000 ;
	    RECT 121.4000 147.8000 121.8000 148.6000 ;
	    RECT 122.2000 147.7000 122.6000 149.9000 ;
	    RECT 124.3000 149.2000 124.9000 149.9000 ;
	    RECT 124.3000 148.9000 125.0000 149.2000 ;
	    RECT 126.6000 148.9000 127.0000 149.9000 ;
	    RECT 128.8000 149.2000 129.2000 149.9000 ;
	    RECT 128.8000 148.9000 129.8000 149.2000 ;
	    RECT 124.6000 148.5000 125.0000 148.9000 ;
	    RECT 126.7000 148.6000 127.0000 148.9000 ;
	    RECT 126.7000 148.3000 128.1000 148.6000 ;
	    RECT 127.7000 148.2000 128.1000 148.3000 ;
	    RECT 128.6000 147.8000 129.0000 148.6000 ;
	    RECT 129.4000 148.5000 129.8000 148.9000 ;
	    RECT 123.7000 147.7000 124.1000 147.8000 ;
	    RECT 122.2000 147.4000 124.1000 147.7000 ;
	    RECT 122.2000 145.7000 122.6000 147.4000 ;
	    RECT 125.7000 147.1000 126.1000 147.2000 ;
	    RECT 128.6000 147.1000 128.9000 147.8000 ;
	    RECT 131.0000 147.5000 131.4000 149.9000 ;
	    RECT 130.2000 147.1000 131.0000 147.2000 ;
	    RECT 125.5000 146.8000 131.0000 147.1000 ;
	    RECT 131.8000 146.8000 132.2000 147.6000 ;
	    RECT 124.6000 146.4000 125.0000 146.5000 ;
	    RECT 123.1000 146.1000 125.0000 146.4000 ;
	    RECT 123.1000 146.0000 123.5000 146.1000 ;
	    RECT 123.9000 145.7000 124.3000 145.8000 ;
	    RECT 122.2000 145.4000 124.3000 145.7000 ;
	    RECT 122.2000 141.1000 122.6000 145.4000 ;
	    RECT 125.5000 145.2000 125.8000 146.8000 ;
	    RECT 129.1000 146.7000 129.5000 146.8000 ;
	    RECT 129.9000 146.2000 130.3000 146.3000 ;
	    RECT 127.8000 145.9000 130.3000 146.2000 ;
	    RECT 132.6000 146.1000 133.0000 149.9000 ;
	    RECT 135.0000 147.9000 135.4000 149.9000 ;
	    RECT 135.7000 148.2000 136.1000 148.6000 ;
	    RECT 134.2000 146.4000 134.6000 147.2000 ;
	    RECT 133.4000 146.1000 133.8000 146.2000 ;
	    RECT 135.0000 146.1000 135.3000 147.9000 ;
	    RECT 135.8000 147.8000 136.2000 148.2000 ;
	    RECT 136.6000 147.8000 137.0000 148.6000 ;
	    RECT 135.8000 146.1000 136.2000 146.2000 ;
	    RECT 127.8000 145.8000 128.2000 145.9000 ;
	    RECT 132.6000 145.8000 134.2000 146.1000 ;
	    RECT 135.0000 145.8000 136.2000 146.1000 ;
	    RECT 137.4000 146.1000 137.8000 149.9000 ;
	    RECT 139.7000 147.9000 140.5000 149.9000 ;
	    RECT 143.5000 147.9000 144.3000 149.9000 ;
	    RECT 138.2000 147.1000 138.6000 147.2000 ;
	    RECT 139.0000 147.1000 139.4000 147.2000 ;
	    RECT 138.2000 146.8000 139.4000 147.1000 ;
	    RECT 139.0000 146.4000 139.4000 146.8000 ;
	    RECT 139.9000 146.2000 140.2000 147.9000 ;
	    RECT 140.6000 146.8000 141.0000 147.2000 ;
	    RECT 143.0000 146.8000 143.4000 147.2000 ;
	    RECT 140.6000 146.6000 140.9000 146.8000 ;
	    RECT 140.5000 146.2000 140.9000 146.6000 ;
	    RECT 143.1000 146.6000 143.4000 146.8000 ;
	    RECT 143.1000 146.2000 143.5000 146.6000 ;
	    RECT 143.8000 146.2000 144.1000 147.9000 ;
	    RECT 144.6000 146.4000 145.0000 147.2000 ;
	    RECT 138.2000 146.1000 138.6000 146.2000 ;
	    RECT 137.4000 145.8000 139.0000 146.1000 ;
	    RECT 139.8000 145.8000 140.2000 146.2000 ;
	    RECT 128.6000 145.5000 131.4000 145.6000 ;
	    RECT 128.5000 145.4000 131.4000 145.5000 ;
	    RECT 124.6000 144.9000 125.8000 145.2000 ;
	    RECT 126.5000 145.3000 131.4000 145.4000 ;
	    RECT 126.5000 145.1000 128.9000 145.3000 ;
	    RECT 124.6000 144.4000 124.9000 144.9000 ;
	    RECT 124.2000 144.0000 124.9000 144.4000 ;
	    RECT 125.7000 144.5000 126.1000 144.6000 ;
	    RECT 126.5000 144.5000 126.8000 145.1000 ;
	    RECT 125.7000 144.2000 126.8000 144.5000 ;
	    RECT 127.1000 144.5000 129.8000 144.8000 ;
	    RECT 127.1000 144.4000 127.5000 144.5000 ;
	    RECT 129.4000 144.4000 129.8000 144.5000 ;
	    RECT 126.3000 143.7000 126.7000 143.8000 ;
	    RECT 127.7000 143.7000 128.1000 143.8000 ;
	    RECT 124.6000 143.1000 125.0000 143.5000 ;
	    RECT 126.3000 143.4000 128.1000 143.7000 ;
	    RECT 126.7000 143.1000 127.0000 143.4000 ;
	    RECT 129.4000 143.1000 129.8000 143.5000 ;
	    RECT 124.3000 141.1000 124.9000 143.1000 ;
	    RECT 126.6000 141.1000 127.0000 143.1000 ;
	    RECT 128.8000 142.8000 129.8000 143.1000 ;
	    RECT 128.8000 141.1000 129.2000 142.8000 ;
	    RECT 131.0000 141.1000 131.4000 145.3000 ;
	    RECT 132.6000 141.1000 133.0000 145.8000 ;
	    RECT 133.8000 145.6000 134.2000 145.8000 ;
	    RECT 135.8000 145.1000 136.1000 145.8000 ;
	    RECT 133.4000 144.8000 135.4000 145.1000 ;
	    RECT 133.4000 141.1000 133.8000 144.8000 ;
	    RECT 135.0000 141.1000 135.4000 144.8000 ;
	    RECT 135.8000 141.1000 136.2000 145.1000 ;
	    RECT 137.4000 141.1000 137.8000 145.8000 ;
	    RECT 138.6000 145.6000 139.0000 145.8000 ;
	    RECT 139.9000 145.7000 140.2000 145.8000 ;
	    RECT 141.4000 146.1000 141.8000 146.2000 ;
	    RECT 142.2000 146.1000 142.6000 146.2000 ;
	    RECT 141.4000 145.8000 142.6000 146.1000 ;
	    RECT 139.9000 145.4000 140.9000 145.7000 ;
	    RECT 141.4000 145.4000 141.8000 145.8000 ;
	    RECT 142.2000 145.4000 142.6000 145.8000 ;
	    RECT 143.8000 145.8000 144.2000 146.2000 ;
	    RECT 145.4000 146.1000 145.8000 146.2000 ;
	    RECT 146.2000 146.1000 146.6000 149.9000 ;
	    RECT 147.0000 148.1000 147.4000 148.6000 ;
	    RECT 147.8000 148.1000 148.2000 149.9000 ;
	    RECT 149.9000 149.2000 150.5000 149.9000 ;
	    RECT 149.9000 148.9000 150.6000 149.2000 ;
	    RECT 152.2000 148.9000 152.6000 149.9000 ;
	    RECT 154.4000 149.2000 154.8000 149.9000 ;
	    RECT 154.4000 148.9000 155.4000 149.2000 ;
	    RECT 150.2000 148.5000 150.6000 148.9000 ;
	    RECT 152.3000 148.6000 152.6000 148.9000 ;
	    RECT 152.3000 148.3000 153.7000 148.6000 ;
	    RECT 153.3000 148.2000 153.7000 148.3000 ;
	    RECT 154.2000 148.2000 154.6000 148.6000 ;
	    RECT 155.0000 148.5000 155.4000 148.9000 ;
	    RECT 147.0000 147.8000 148.2000 148.1000 ;
	    RECT 149.4000 147.8000 149.8000 148.2000 ;
	    RECT 145.0000 145.8000 146.6000 146.1000 ;
	    RECT 143.8000 145.7000 144.1000 145.8000 ;
	    RECT 143.1000 145.4000 144.1000 145.7000 ;
	    RECT 145.0000 145.6000 145.4000 145.8000 ;
	    RECT 140.6000 145.1000 140.9000 145.4000 ;
	    RECT 143.1000 145.1000 143.4000 145.4000 ;
	    RECT 138.2000 144.8000 140.2000 145.1000 ;
	    RECT 138.2000 141.1000 138.6000 144.8000 ;
	    RECT 139.8000 141.4000 140.2000 144.8000 ;
	    RECT 140.6000 141.7000 141.0000 145.1000 ;
	    RECT 141.4000 141.4000 141.8000 145.1000 ;
	    RECT 139.8000 141.1000 141.8000 141.4000 ;
	    RECT 142.2000 141.4000 142.6000 145.1000 ;
	    RECT 143.0000 141.7000 143.4000 145.1000 ;
	    RECT 143.8000 144.8000 145.8000 145.1000 ;
	    RECT 143.8000 141.4000 144.2000 144.8000 ;
	    RECT 142.2000 141.1000 144.2000 141.4000 ;
	    RECT 145.4000 141.1000 145.8000 144.8000 ;
	    RECT 146.2000 141.1000 146.6000 145.8000 ;
	    RECT 147.8000 147.7000 148.2000 147.8000 ;
	    RECT 149.3000 147.7000 149.8000 147.8000 ;
	    RECT 147.8000 147.4000 149.8000 147.7000 ;
	    RECT 147.8000 145.7000 148.2000 147.4000 ;
	    RECT 151.3000 147.1000 151.7000 147.2000 ;
	    RECT 154.2000 147.1000 154.5000 148.2000 ;
	    RECT 156.6000 147.5000 157.0000 149.9000 ;
	    RECT 158.2000 148.2000 158.6000 149.9000 ;
	    RECT 158.1000 147.9000 158.6000 148.2000 ;
	    RECT 158.1000 147.2000 158.4000 147.9000 ;
	    RECT 159.8000 147.6000 160.2000 149.9000 ;
	    RECT 158.9000 147.3000 160.2000 147.6000 ;
	    RECT 162.2000 147.5000 162.6000 149.9000 ;
	    RECT 164.4000 149.2000 164.8000 149.9000 ;
	    RECT 163.8000 148.9000 164.8000 149.2000 ;
	    RECT 166.6000 148.9000 167.0000 149.9000 ;
	    RECT 168.7000 149.2000 169.3000 149.9000 ;
	    RECT 168.6000 148.9000 169.3000 149.2000 ;
	    RECT 163.8000 148.5000 164.2000 148.9000 ;
	    RECT 166.6000 148.6000 166.9000 148.9000 ;
	    RECT 164.6000 148.2000 165.0000 148.6000 ;
	    RECT 165.5000 148.3000 166.9000 148.6000 ;
	    RECT 168.6000 148.5000 169.0000 148.9000 ;
	    RECT 165.5000 148.2000 165.9000 148.3000 ;
	    RECT 155.8000 147.1000 156.6000 147.2000 ;
	    RECT 151.1000 146.8000 156.6000 147.1000 ;
	    RECT 158.1000 146.8000 158.6000 147.2000 ;
	    RECT 150.2000 146.4000 150.6000 146.5000 ;
	    RECT 148.7000 146.1000 150.6000 146.4000 ;
	    RECT 151.1000 146.1000 151.4000 146.8000 ;
	    RECT 154.7000 146.7000 155.1000 146.8000 ;
	    RECT 155.5000 146.2000 155.9000 146.3000 ;
	    RECT 151.8000 146.1000 152.2000 146.2000 ;
	    RECT 148.7000 146.0000 149.1000 146.1000 ;
	    RECT 151.0000 145.8000 152.2000 146.1000 ;
	    RECT 153.4000 145.9000 155.9000 146.2000 ;
	    RECT 153.4000 145.8000 153.8000 145.9000 ;
	    RECT 149.5000 145.7000 149.9000 145.8000 ;
	    RECT 147.8000 145.4000 149.9000 145.7000 ;
	    RECT 147.8000 141.1000 148.2000 145.4000 ;
	    RECT 151.1000 145.2000 151.4000 145.8000 ;
	    RECT 154.2000 145.5000 157.0000 145.6000 ;
	    RECT 154.1000 145.4000 157.0000 145.5000 ;
	    RECT 150.2000 144.9000 151.4000 145.2000 ;
	    RECT 152.1000 145.3000 157.0000 145.4000 ;
	    RECT 152.1000 145.1000 154.5000 145.3000 ;
	    RECT 150.2000 144.4000 150.5000 144.9000 ;
	    RECT 149.8000 144.0000 150.5000 144.4000 ;
	    RECT 151.3000 144.5000 151.7000 144.6000 ;
	    RECT 152.1000 144.5000 152.4000 145.1000 ;
	    RECT 151.3000 144.2000 152.4000 144.5000 ;
	    RECT 152.7000 144.5000 155.4000 144.8000 ;
	    RECT 152.7000 144.4000 153.1000 144.5000 ;
	    RECT 155.0000 144.4000 155.4000 144.5000 ;
	    RECT 151.9000 143.7000 152.3000 143.8000 ;
	    RECT 153.3000 143.7000 153.7000 143.8000 ;
	    RECT 150.2000 143.1000 150.6000 143.5000 ;
	    RECT 151.9000 143.4000 153.7000 143.7000 ;
	    RECT 152.3000 143.1000 152.6000 143.4000 ;
	    RECT 155.0000 143.1000 155.4000 143.5000 ;
	    RECT 149.9000 141.1000 150.5000 143.1000 ;
	    RECT 152.2000 141.1000 152.6000 143.1000 ;
	    RECT 154.4000 142.8000 155.4000 143.1000 ;
	    RECT 154.4000 141.1000 154.8000 142.8000 ;
	    RECT 156.6000 141.1000 157.0000 145.3000 ;
	    RECT 158.1000 145.1000 158.4000 146.8000 ;
	    RECT 158.9000 146.5000 159.2000 147.3000 ;
	    RECT 162.6000 147.1000 163.4000 147.2000 ;
	    RECT 164.7000 147.1000 165.0000 148.2000 ;
	    RECT 169.5000 147.7000 169.9000 147.8000 ;
	    RECT 171.0000 147.7000 171.4000 149.9000 ;
	    RECT 171.8000 147.8000 172.2000 148.6000 ;
	    RECT 172.6000 148.1000 173.0000 149.9000 ;
	    RECT 174.2000 148.9000 174.6000 149.9000 ;
	    RECT 173.4000 148.1000 173.8000 148.6000 ;
	    RECT 172.6000 147.8000 173.8000 148.1000 ;
	    RECT 169.5000 147.4000 171.4000 147.7000 ;
	    RECT 167.5000 147.1000 167.9000 147.2000 ;
	    RECT 162.6000 146.8000 168.1000 147.1000 ;
	    RECT 164.1000 146.7000 164.5000 146.8000 ;
	    RECT 158.7000 146.1000 159.2000 146.5000 ;
	    RECT 158.9000 145.1000 159.2000 146.1000 ;
	    RECT 159.7000 146.2000 160.1000 146.6000 ;
	    RECT 163.3000 146.2000 163.7000 146.3000 ;
	    RECT 159.7000 145.8000 160.2000 146.2000 ;
	    RECT 163.3000 145.9000 165.8000 146.2000 ;
	    RECT 165.4000 145.8000 165.8000 145.9000 ;
	    RECT 167.0000 146.1000 167.4000 146.2000 ;
	    RECT 167.8000 146.1000 168.1000 146.8000 ;
	    RECT 168.6000 146.4000 169.0000 146.5000 ;
	    RECT 168.6000 146.1000 170.5000 146.4000 ;
	    RECT 167.0000 145.8000 168.1000 146.1000 ;
	    RECT 170.1000 146.0000 170.5000 146.1000 ;
	    RECT 162.2000 145.5000 165.0000 145.6000 ;
	    RECT 162.2000 145.4000 165.1000 145.5000 ;
	    RECT 162.2000 145.3000 167.1000 145.4000 ;
	    RECT 158.1000 144.6000 158.6000 145.1000 ;
	    RECT 158.9000 144.8000 160.2000 145.1000 ;
	    RECT 158.2000 141.1000 158.6000 144.6000 ;
	    RECT 159.8000 141.1000 160.2000 144.8000 ;
	    RECT 162.2000 141.1000 162.6000 145.3000 ;
	    RECT 164.7000 145.1000 167.1000 145.3000 ;
	    RECT 163.8000 144.5000 166.5000 144.8000 ;
	    RECT 163.8000 144.4000 164.2000 144.5000 ;
	    RECT 166.1000 144.4000 166.5000 144.5000 ;
	    RECT 166.8000 144.5000 167.1000 145.1000 ;
	    RECT 167.8000 145.2000 168.1000 145.8000 ;
	    RECT 169.3000 145.7000 169.7000 145.8000 ;
	    RECT 171.0000 145.7000 171.4000 147.4000 ;
	    RECT 169.3000 145.4000 171.4000 145.7000 ;
	    RECT 167.8000 144.9000 169.0000 145.2000 ;
	    RECT 167.5000 144.5000 167.9000 144.6000 ;
	    RECT 166.8000 144.2000 167.9000 144.5000 ;
	    RECT 168.7000 144.4000 169.0000 144.9000 ;
	    RECT 168.7000 144.0000 169.4000 144.4000 ;
	    RECT 165.5000 143.7000 165.9000 143.8000 ;
	    RECT 166.9000 143.7000 167.3000 143.8000 ;
	    RECT 163.8000 143.1000 164.2000 143.5000 ;
	    RECT 165.5000 143.4000 167.3000 143.7000 ;
	    RECT 166.6000 143.1000 166.9000 143.4000 ;
	    RECT 168.6000 143.1000 169.0000 143.5000 ;
	    RECT 163.8000 142.8000 164.8000 143.1000 ;
	    RECT 164.4000 141.1000 164.8000 142.8000 ;
	    RECT 166.6000 141.1000 167.0000 143.1000 ;
	    RECT 168.7000 141.1000 169.3000 143.1000 ;
	    RECT 171.0000 141.1000 171.4000 145.4000 ;
	    RECT 172.6000 141.1000 173.0000 147.8000 ;
	    RECT 174.3000 147.2000 174.6000 148.9000 ;
	    RECT 175.8000 147.9000 176.2000 149.9000 ;
	    RECT 176.6000 148.0000 177.0000 149.9000 ;
	    RECT 178.2000 148.0000 178.6000 149.9000 ;
	    RECT 179.3000 148.4000 179.7000 149.9000 ;
	    RECT 176.6000 147.9000 178.6000 148.0000 ;
	    RECT 179.0000 147.9000 179.7000 148.4000 ;
	    RECT 181.4000 147.9000 181.8000 149.9000 ;
	    RECT 175.9000 147.2000 176.2000 147.9000 ;
	    RECT 176.7000 147.7000 178.5000 147.9000 ;
	    RECT 177.8000 147.2000 178.2000 147.4000 ;
	    RECT 173.4000 146.8000 173.8000 147.2000 ;
	    RECT 174.2000 146.8000 174.6000 147.2000 ;
	    RECT 175.8000 146.8000 177.1000 147.2000 ;
	    RECT 177.8000 146.9000 178.6000 147.2000 ;
	    RECT 178.2000 146.8000 178.6000 146.9000 ;
	    RECT 173.4000 146.1000 173.7000 146.8000 ;
	    RECT 174.3000 146.1000 174.6000 146.8000 ;
	    RECT 173.4000 145.8000 174.6000 146.1000 ;
	    RECT 174.3000 145.1000 174.6000 145.8000 ;
	    RECT 175.0000 146.1000 175.4000 146.2000 ;
	    RECT 176.8000 146.1000 177.1000 146.8000 ;
	    RECT 175.0000 145.8000 177.1000 146.1000 ;
	    RECT 177.4000 145.8000 177.8000 146.6000 ;
	    RECT 179.0000 146.2000 179.3000 147.9000 ;
	    RECT 181.4000 147.8000 181.7000 147.9000 ;
	    RECT 182.2000 147.8000 182.6000 148.6000 ;
	    RECT 180.8000 147.6000 181.7000 147.8000 ;
	    RECT 179.6000 147.5000 181.7000 147.6000 ;
	    RECT 179.6000 147.3000 181.1000 147.5000 ;
	    RECT 179.6000 147.2000 180.0000 147.3000 ;
	    RECT 179.0000 145.8000 179.4000 146.2000 ;
	    RECT 175.0000 145.4000 175.4000 145.8000 ;
	    RECT 175.8000 145.1000 176.2000 145.2000 ;
	    RECT 176.8000 145.1000 177.1000 145.8000 ;
	    RECT 179.0000 145.1000 179.3000 145.8000 ;
	    RECT 179.7000 145.5000 180.0000 147.2000 ;
	    RECT 180.4000 146.6000 181.0000 147.0000 ;
	    RECT 180.6000 146.2000 180.9000 146.6000 ;
	    RECT 181.4000 146.4000 181.8000 147.2000 ;
	    RECT 180.6000 145.8000 181.0000 146.2000 ;
	    RECT 183.0000 146.1000 183.4000 149.9000 ;
	    RECT 184.6000 148.9000 185.0000 149.9000 ;
	    RECT 187.0000 148.9000 187.4000 149.9000 ;
	    RECT 184.6000 147.2000 184.9000 148.9000 ;
	    RECT 185.4000 147.8000 185.8000 148.6000 ;
	    RECT 186.2000 147.8000 186.6000 148.6000 ;
	    RECT 187.1000 147.2000 187.4000 148.9000 ;
	    RECT 188.6000 148.0000 189.0000 149.9000 ;
	    RECT 190.2000 148.0000 190.6000 149.9000 ;
	    RECT 188.6000 147.9000 190.6000 148.0000 ;
	    RECT 191.0000 147.9000 191.4000 149.9000 ;
	    RECT 192.6000 148.9000 193.0000 149.9000 ;
	    RECT 188.7000 147.7000 190.5000 147.9000 ;
	    RECT 189.0000 147.2000 189.4000 147.4000 ;
	    RECT 191.0000 147.2000 191.3000 147.9000 ;
	    RECT 191.8000 147.8000 192.2000 148.6000 ;
	    RECT 192.7000 147.2000 193.0000 148.9000 ;
	    RECT 194.2000 148.0000 194.6000 149.9000 ;
	    RECT 195.8000 148.0000 196.2000 149.9000 ;
	    RECT 194.2000 147.9000 196.2000 148.0000 ;
	    RECT 196.6000 147.9000 197.0000 149.9000 ;
	    RECT 194.3000 147.7000 196.1000 147.9000 ;
	    RECT 194.6000 147.2000 195.0000 147.4000 ;
	    RECT 196.6000 147.2000 196.9000 147.9000 ;
	    RECT 197.4000 147.7000 197.8000 149.9000 ;
	    RECT 199.5000 149.2000 200.1000 149.9000 ;
	    RECT 199.5000 148.9000 200.2000 149.2000 ;
	    RECT 201.8000 148.9000 202.2000 149.9000 ;
	    RECT 204.0000 149.2000 204.4000 149.9000 ;
	    RECT 204.0000 148.9000 205.0000 149.2000 ;
	    RECT 199.8000 148.5000 200.2000 148.9000 ;
	    RECT 201.9000 148.6000 202.2000 148.9000 ;
	    RECT 201.9000 148.3000 203.3000 148.6000 ;
	    RECT 202.9000 148.2000 203.3000 148.3000 ;
	    RECT 203.8000 148.2000 204.2000 148.6000 ;
	    RECT 204.6000 148.5000 205.0000 148.9000 ;
	    RECT 198.9000 147.7000 199.3000 147.8000 ;
	    RECT 197.4000 147.4000 199.3000 147.7000 ;
	    RECT 184.6000 147.1000 185.0000 147.2000 ;
	    RECT 185.4000 147.1000 185.8000 147.2000 ;
	    RECT 184.6000 146.8000 185.8000 147.1000 ;
	    RECT 187.0000 146.8000 187.4000 147.2000 ;
	    RECT 188.6000 146.9000 189.4000 147.2000 ;
	    RECT 188.6000 146.8000 189.0000 146.9000 ;
	    RECT 190.1000 146.8000 191.4000 147.2000 ;
	    RECT 192.6000 146.8000 193.0000 147.2000 ;
	    RECT 193.4000 147.1000 193.8000 147.2000 ;
	    RECT 194.2000 147.1000 195.0000 147.2000 ;
	    RECT 193.4000 146.9000 195.0000 147.1000 ;
	    RECT 193.4000 146.8000 194.6000 146.9000 ;
	    RECT 195.7000 146.8000 197.0000 147.2000 ;
	    RECT 183.8000 146.1000 184.2000 146.2000 ;
	    RECT 183.0000 145.8000 184.2000 146.1000 ;
	    RECT 179.7000 145.2000 180.9000 145.5000 ;
	    RECT 174.2000 144.7000 175.1000 145.1000 ;
	    RECT 175.8000 144.8000 176.5000 145.1000 ;
	    RECT 176.8000 144.8000 177.3000 145.1000 ;
	    RECT 174.7000 141.1000 175.1000 144.7000 ;
	    RECT 176.2000 144.2000 176.5000 144.8000 ;
	    RECT 176.2000 143.8000 176.6000 144.2000 ;
	    RECT 176.9000 141.1000 177.3000 144.8000 ;
	    RECT 179.0000 141.1000 179.4000 145.1000 ;
	    RECT 180.6000 143.1000 180.9000 145.2000 ;
	    RECT 180.6000 141.1000 181.0000 143.1000 ;
	    RECT 183.0000 141.1000 183.4000 145.8000 ;
	    RECT 183.8000 145.4000 184.2000 145.8000 ;
	    RECT 184.6000 145.1000 184.9000 146.8000 ;
	    RECT 187.1000 145.1000 187.4000 146.8000 ;
	    RECT 187.8000 145.4000 188.2000 146.2000 ;
	    RECT 189.4000 145.8000 189.8000 146.6000 ;
	    RECT 190.1000 145.1000 190.4000 146.8000 ;
	    RECT 191.0000 146.2000 191.3000 146.8000 ;
	    RECT 191.0000 145.8000 191.4000 146.2000 ;
	    RECT 191.0000 145.1000 191.4000 145.2000 ;
	    RECT 192.7000 145.1000 193.0000 146.8000 ;
	    RECT 193.4000 145.4000 193.8000 146.2000 ;
	    RECT 194.2000 146.1000 194.6000 146.2000 ;
	    RECT 195.0000 146.1000 195.4000 146.6000 ;
	    RECT 194.2000 145.8000 195.4000 146.1000 ;
	    RECT 195.7000 146.1000 196.0000 146.8000 ;
	    RECT 196.6000 146.1000 197.0000 146.2000 ;
	    RECT 195.7000 145.8000 197.0000 146.1000 ;
	    RECT 195.7000 145.1000 196.0000 145.8000 ;
	    RECT 197.4000 145.7000 197.8000 147.4000 ;
	    RECT 200.9000 147.1000 201.3000 147.2000 ;
	    RECT 203.0000 147.1000 203.4000 147.2000 ;
	    RECT 203.8000 147.1000 204.1000 148.2000 ;
	    RECT 206.2000 147.5000 206.6000 149.9000 ;
	    RECT 207.1000 148.2000 207.5000 148.6000 ;
	    RECT 207.0000 147.8000 207.4000 148.2000 ;
	    RECT 207.8000 147.8000 208.2000 149.9000 ;
	    RECT 210.5000 148.2000 210.9000 149.9000 ;
	    RECT 210.5000 147.9000 211.4000 148.2000 ;
	    RECT 205.4000 147.1000 206.2000 147.2000 ;
	    RECT 200.7000 146.8000 206.2000 147.1000 ;
	    RECT 199.8000 146.4000 200.2000 146.5000 ;
	    RECT 198.3000 146.1000 200.2000 146.4000 ;
	    RECT 198.3000 146.0000 198.7000 146.1000 ;
	    RECT 199.1000 145.7000 199.5000 145.8000 ;
	    RECT 197.4000 145.4000 199.5000 145.7000 ;
	    RECT 196.6000 145.1000 197.0000 145.2000 ;
	    RECT 197.4000 145.1000 197.8000 145.4000 ;
	    RECT 200.7000 145.2000 201.0000 146.8000 ;
	    RECT 204.3000 146.7000 204.7000 146.8000 ;
	    RECT 203.8000 146.2000 204.2000 146.3000 ;
	    RECT 205.1000 146.2000 205.5000 146.3000 ;
	    RECT 203.0000 145.9000 205.5000 146.2000 ;
	    RECT 207.0000 146.1000 207.4000 146.2000 ;
	    RECT 207.9000 146.1000 208.2000 147.8000 ;
	    RECT 208.6000 147.1000 209.0000 147.2000 ;
	    RECT 211.0000 147.1000 211.4000 147.9000 ;
	    RECT 215.8000 147.9000 216.2000 149.9000 ;
	    RECT 216.5000 148.2000 216.9000 148.6000 ;
	    RECT 208.6000 146.8000 211.4000 147.1000 ;
	    RECT 211.8000 146.8000 212.2000 147.6000 ;
	    RECT 213.4000 147.1000 213.8000 147.2000 ;
	    RECT 215.0000 147.1000 215.4000 147.2000 ;
	    RECT 213.4000 146.8000 215.4000 147.1000 ;
	    RECT 208.6000 146.4000 209.0000 146.8000 ;
	    RECT 209.4000 146.1000 209.8000 146.2000 ;
	    RECT 203.0000 145.8000 203.4000 145.9000 ;
	    RECT 207.0000 145.8000 208.2000 146.1000 ;
	    RECT 209.0000 145.8000 209.8000 146.1000 ;
	    RECT 203.8000 145.5000 206.6000 145.6000 ;
	    RECT 203.7000 145.4000 206.6000 145.5000 ;
	    RECT 184.1000 144.7000 185.0000 145.1000 ;
	    RECT 187.0000 144.7000 187.9000 145.1000 ;
	    RECT 184.1000 141.1000 184.5000 144.7000 ;
	    RECT 187.5000 144.2000 187.9000 144.7000 ;
	    RECT 189.9000 144.8000 190.4000 145.1000 ;
	    RECT 190.7000 144.8000 191.4000 145.1000 ;
	    RECT 187.5000 143.8000 188.2000 144.2000 ;
	    RECT 187.5000 141.1000 187.9000 143.8000 ;
	    RECT 189.9000 141.1000 190.3000 144.8000 ;
	    RECT 190.7000 144.2000 191.0000 144.8000 ;
	    RECT 192.6000 144.7000 193.5000 145.1000 ;
	    RECT 190.6000 143.8000 191.0000 144.2000 ;
	    RECT 193.1000 143.2000 193.5000 144.7000 ;
	    RECT 195.5000 144.8000 196.0000 145.1000 ;
	    RECT 196.3000 144.8000 197.8000 145.1000 ;
	    RECT 193.1000 142.8000 193.8000 143.2000 ;
	    RECT 193.1000 141.1000 193.5000 142.8000 ;
	    RECT 195.5000 141.1000 195.9000 144.8000 ;
	    RECT 196.3000 144.2000 196.6000 144.8000 ;
	    RECT 196.2000 143.8000 196.6000 144.2000 ;
	    RECT 197.4000 141.1000 197.8000 144.8000 ;
	    RECT 199.8000 144.9000 201.0000 145.2000 ;
	    RECT 201.7000 145.3000 206.6000 145.4000 ;
	    RECT 201.7000 145.1000 204.1000 145.3000 ;
	    RECT 199.8000 144.4000 200.1000 144.9000 ;
	    RECT 199.4000 144.0000 200.1000 144.4000 ;
	    RECT 200.9000 144.5000 201.3000 144.6000 ;
	    RECT 201.7000 144.5000 202.0000 145.1000 ;
	    RECT 200.9000 144.2000 202.0000 144.5000 ;
	    RECT 202.3000 144.5000 205.0000 144.8000 ;
	    RECT 202.3000 144.4000 202.7000 144.5000 ;
	    RECT 204.6000 144.4000 205.0000 144.5000 ;
	    RECT 201.5000 143.7000 201.9000 143.8000 ;
	    RECT 202.9000 143.7000 203.3000 143.8000 ;
	    RECT 199.8000 143.1000 200.2000 143.5000 ;
	    RECT 201.5000 143.4000 203.3000 143.7000 ;
	    RECT 201.9000 143.1000 202.2000 143.4000 ;
	    RECT 204.6000 143.1000 205.0000 143.5000 ;
	    RECT 199.5000 141.1000 200.1000 143.1000 ;
	    RECT 201.8000 141.1000 202.2000 143.1000 ;
	    RECT 204.0000 142.8000 205.0000 143.1000 ;
	    RECT 204.0000 141.1000 204.4000 142.8000 ;
	    RECT 206.2000 141.1000 206.6000 145.3000 ;
	    RECT 207.1000 145.1000 207.4000 145.8000 ;
	    RECT 209.0000 145.6000 209.4000 145.8000 ;
	    RECT 207.0000 141.1000 207.4000 145.1000 ;
	    RECT 207.8000 144.8000 209.8000 145.1000 ;
	    RECT 207.8000 141.1000 208.2000 144.8000 ;
	    RECT 209.4000 141.1000 209.8000 144.8000 ;
	    RECT 210.2000 144.4000 210.6000 145.2000 ;
	    RECT 211.0000 141.1000 211.4000 146.8000 ;
	    RECT 215.0000 146.4000 215.4000 146.8000 ;
	    RECT 214.2000 146.1000 214.6000 146.2000 ;
	    RECT 215.8000 146.1000 216.1000 147.9000 ;
	    RECT 216.6000 147.8000 217.0000 148.2000 ;
	    RECT 219.0000 147.9000 219.4000 149.9000 ;
	    RECT 219.7000 148.2000 220.1000 148.6000 ;
	    RECT 219.8000 148.1000 220.2000 148.2000 ;
	    RECT 220.6000 148.1000 221.0000 149.9000 ;
	    RECT 218.2000 146.4000 218.6000 147.2000 ;
	    RECT 216.6000 146.1000 217.0000 146.2000 ;
	    RECT 217.4000 146.1000 217.8000 146.2000 ;
	    RECT 219.0000 146.1000 219.3000 147.9000 ;
	    RECT 219.8000 147.8000 221.0000 148.1000 ;
	    RECT 221.4000 148.0000 221.8000 149.9000 ;
	    RECT 223.0000 148.0000 223.4000 149.9000 ;
	    RECT 221.4000 147.9000 223.4000 148.0000 ;
	    RECT 224.6000 148.9000 225.0000 149.9000 ;
	    RECT 227.0000 148.9000 227.4000 149.9000 ;
	    RECT 220.7000 147.2000 221.0000 147.8000 ;
	    RECT 221.5000 147.7000 223.3000 147.9000 ;
	    RECT 222.6000 147.2000 223.0000 147.4000 ;
	    RECT 224.6000 147.2000 224.9000 148.9000 ;
	    RECT 225.4000 148.1000 225.8000 148.6000 ;
	    RECT 226.2000 148.1000 226.6000 148.6000 ;
	    RECT 225.4000 147.8000 226.6000 148.1000 ;
	    RECT 227.1000 147.2000 227.4000 148.9000 ;
	    RECT 229.4000 148.9000 229.8000 149.9000 ;
	    RECT 229.4000 147.2000 229.7000 148.9000 ;
	    RECT 230.2000 147.8000 230.6000 148.6000 ;
	    RECT 231.0000 147.6000 231.4000 149.9000 ;
	    RECT 232.6000 148.2000 233.0000 149.9000 ;
	    RECT 232.6000 147.9000 233.1000 148.2000 ;
	    RECT 231.0000 147.3000 232.3000 147.6000 ;
	    RECT 220.6000 146.8000 221.9000 147.2000 ;
	    RECT 222.6000 146.9000 223.4000 147.2000 ;
	    RECT 223.0000 146.8000 223.4000 146.9000 ;
	    RECT 224.6000 146.8000 225.0000 147.2000 ;
	    RECT 225.4000 147.1000 225.8000 147.2000 ;
	    RECT 227.0000 147.1000 227.4000 147.2000 ;
	    RECT 225.4000 146.8000 227.4000 147.1000 ;
	    RECT 228.6000 147.1000 229.0000 147.2000 ;
	    RECT 229.4000 147.1000 229.8000 147.2000 ;
	    RECT 228.6000 146.8000 229.8000 147.1000 ;
	    RECT 219.8000 146.1000 220.2000 146.2000 ;
	    RECT 214.2000 145.8000 215.0000 146.1000 ;
	    RECT 215.8000 145.8000 218.2000 146.1000 ;
	    RECT 219.0000 145.8000 220.2000 146.1000 ;
	    RECT 214.6000 145.6000 215.0000 145.8000 ;
	    RECT 216.6000 145.1000 216.9000 145.8000 ;
	    RECT 217.8000 145.6000 218.2000 145.8000 ;
	    RECT 219.8000 145.1000 220.1000 145.8000 ;
	    RECT 220.6000 145.1000 221.0000 145.2000 ;
	    RECT 221.6000 145.1000 221.9000 146.8000 ;
	    RECT 222.2000 145.8000 222.6000 146.6000 ;
	    RECT 223.0000 146.1000 223.4000 146.2000 ;
	    RECT 223.8000 146.1000 224.2000 146.2000 ;
	    RECT 223.0000 145.8000 224.2000 146.1000 ;
	    RECT 223.8000 145.4000 224.2000 145.8000 ;
	    RECT 224.6000 145.1000 224.9000 146.8000 ;
	    RECT 227.1000 145.1000 227.4000 146.8000 ;
	    RECT 227.8000 145.4000 228.2000 146.2000 ;
	    RECT 228.6000 145.4000 229.0000 146.2000 ;
	    RECT 229.4000 145.1000 229.7000 146.8000 ;
	    RECT 231.1000 146.2000 231.5000 146.6000 ;
	    RECT 231.0000 145.8000 231.5000 146.2000 ;
	    RECT 232.0000 146.5000 232.3000 147.3000 ;
	    RECT 232.8000 147.2000 233.1000 147.9000 ;
	    RECT 234.2000 147.6000 234.6000 149.9000 ;
	    RECT 235.8000 148.2000 236.2000 149.9000 ;
	    RECT 238.2000 148.8000 238.6000 149.9000 ;
	    RECT 235.8000 147.9000 236.3000 148.2000 ;
	    RECT 234.2000 147.3000 235.5000 147.6000 ;
	    RECT 232.6000 146.8000 233.1000 147.2000 ;
	    RECT 232.0000 146.1000 232.5000 146.5000 ;
	    RECT 232.0000 145.1000 232.3000 146.1000 ;
	    RECT 232.8000 145.1000 233.1000 146.8000 ;
	    RECT 233.4000 146.8000 233.8000 147.2000 ;
	    RECT 233.4000 146.1000 233.7000 146.8000 ;
	    RECT 234.3000 146.2000 234.7000 146.6000 ;
	    RECT 234.2000 146.1000 234.7000 146.2000 ;
	    RECT 233.4000 145.8000 234.7000 146.1000 ;
	    RECT 235.2000 146.5000 235.5000 147.3000 ;
	    RECT 236.0000 147.2000 236.3000 147.9000 ;
	    RECT 235.8000 146.8000 236.3000 147.2000 ;
	    RECT 235.2000 146.1000 235.7000 146.5000 ;
	    RECT 235.2000 145.1000 235.5000 146.1000 ;
	    RECT 236.0000 145.1000 236.3000 146.8000 ;
	    RECT 238.2000 147.2000 238.5000 148.8000 ;
	    RECT 239.0000 147.8000 239.4000 148.6000 ;
	    RECT 239.8000 147.8000 240.2000 148.6000 ;
	    RECT 238.2000 146.8000 238.6000 147.2000 ;
	    RECT 237.4000 145.4000 237.8000 146.2000 ;
	    RECT 238.2000 145.1000 238.5000 146.8000 ;
	    RECT 239.8000 145.1000 240.2000 145.2000 ;
	    RECT 240.6000 145.1000 241.0000 149.9000 ;
	    RECT 242.2000 148.9000 242.6000 149.9000 ;
	    RECT 242.2000 147.2000 242.5000 148.9000 ;
	    RECT 243.0000 147.8000 243.4000 148.6000 ;
	    RECT 242.2000 146.8000 242.6000 147.2000 ;
	    RECT 245.6000 147.1000 246.0000 149.9000 ;
	    RECT 247.8000 148.8000 248.2000 149.9000 ;
	    RECT 247.8000 147.2000 248.1000 148.8000 ;
	    RECT 248.6000 147.8000 249.0000 148.6000 ;
	    RECT 249.4000 147.9000 249.8000 149.9000 ;
	    RECT 250.2000 148.0000 250.6000 149.9000 ;
	    RECT 251.8000 148.0000 252.2000 149.9000 ;
	    RECT 250.2000 147.9000 252.2000 148.0000 ;
	    RECT 252.6000 147.9000 253.0000 149.9000 ;
	    RECT 253.4000 148.0000 253.8000 149.9000 ;
	    RECT 255.0000 148.0000 255.4000 149.9000 ;
	    RECT 256.1000 148.4000 256.5000 149.9000 ;
	    RECT 253.4000 147.9000 255.4000 148.0000 ;
	    RECT 255.8000 147.9000 256.5000 148.4000 ;
	    RECT 258.2000 147.9000 258.6000 149.9000 ;
	    RECT 259.8000 148.9000 260.2000 149.9000 ;
	    RECT 249.5000 147.2000 249.8000 147.9000 ;
	    RECT 250.3000 147.7000 252.1000 147.9000 ;
	    RECT 251.4000 147.2000 251.8000 147.4000 ;
	    RECT 252.7000 147.2000 253.0000 147.9000 ;
	    RECT 253.5000 147.7000 255.3000 147.9000 ;
	    RECT 254.6000 147.2000 255.0000 147.4000 ;
	    RECT 245.6000 146.9000 246.5000 147.1000 ;
	    RECT 245.7000 146.8000 246.5000 146.9000 ;
	    RECT 241.4000 145.4000 241.8000 146.2000 ;
	    RECT 242.2000 146.1000 242.5000 146.8000 ;
	    RECT 243.0000 146.1000 243.4000 146.2000 ;
	    RECT 242.2000 145.8000 243.4000 146.1000 ;
	    RECT 244.6000 145.8000 245.4000 146.2000 ;
	    RECT 242.2000 145.1000 242.5000 145.8000 ;
	    RECT 214.2000 144.8000 216.2000 145.1000 ;
	    RECT 214.2000 141.1000 214.6000 144.8000 ;
	    RECT 215.8000 141.1000 216.2000 144.8000 ;
	    RECT 216.6000 141.1000 217.0000 145.1000 ;
	    RECT 217.4000 144.8000 219.4000 145.1000 ;
	    RECT 217.4000 141.1000 217.8000 144.8000 ;
	    RECT 219.0000 141.1000 219.4000 144.8000 ;
	    RECT 219.8000 141.1000 220.2000 145.1000 ;
	    RECT 220.6000 144.8000 221.3000 145.1000 ;
	    RECT 221.6000 144.8000 222.1000 145.1000 ;
	    RECT 221.0000 144.2000 221.3000 144.8000 ;
	    RECT 221.0000 143.8000 221.4000 144.2000 ;
	    RECT 221.7000 141.1000 222.1000 144.8000 ;
	    RECT 224.1000 144.7000 225.0000 145.1000 ;
	    RECT 227.0000 144.7000 227.9000 145.1000 ;
	    RECT 224.1000 144.2000 224.5000 144.7000 ;
	    RECT 223.8000 143.8000 224.5000 144.2000 ;
	    RECT 224.1000 141.1000 224.5000 143.8000 ;
	    RECT 227.5000 141.1000 227.9000 144.7000 ;
	    RECT 228.9000 144.7000 229.8000 145.1000 ;
	    RECT 231.0000 144.8000 232.3000 145.1000 ;
	    RECT 228.9000 141.1000 229.3000 144.7000 ;
	    RECT 231.0000 141.1000 231.4000 144.8000 ;
	    RECT 232.6000 144.6000 233.1000 145.1000 ;
	    RECT 234.2000 144.8000 235.5000 145.1000 ;
	    RECT 232.6000 141.1000 233.0000 144.6000 ;
	    RECT 234.2000 141.1000 234.6000 144.8000 ;
	    RECT 235.8000 144.6000 236.3000 145.1000 ;
	    RECT 237.7000 144.7000 238.6000 145.1000 ;
	    RECT 239.8000 144.8000 241.0000 145.1000 ;
	    RECT 235.8000 141.1000 236.2000 144.6000 ;
	    RECT 237.7000 141.1000 238.1000 144.7000 ;
	    RECT 240.6000 141.1000 241.0000 144.8000 ;
	    RECT 241.7000 144.7000 242.6000 145.1000 ;
	    RECT 243.8000 144.8000 244.2000 145.6000 ;
	    RECT 246.2000 145.2000 246.5000 146.8000 ;
	    RECT 247.8000 146.8000 248.2000 147.2000 ;
	    RECT 249.4000 146.8000 250.7000 147.2000 ;
	    RECT 251.4000 146.9000 252.2000 147.2000 ;
	    RECT 251.8000 146.8000 252.2000 146.9000 ;
	    RECT 252.6000 146.8000 253.9000 147.2000 ;
	    RECT 254.6000 146.9000 255.4000 147.2000 ;
	    RECT 247.0000 145.4000 247.4000 146.2000 ;
	    RECT 246.2000 144.8000 246.6000 145.2000 ;
	    RECT 247.8000 145.1000 248.1000 146.8000 ;
	    RECT 249.4000 145.1000 249.8000 145.2000 ;
	    RECT 250.4000 145.1000 250.7000 146.8000 ;
	    RECT 251.0000 145.8000 251.4000 146.6000 ;
	    RECT 252.6000 145.1000 253.0000 145.2000 ;
	    RECT 253.6000 145.1000 253.9000 146.8000 ;
	    RECT 255.0000 146.8000 255.4000 146.9000 ;
	    RECT 254.2000 145.8000 254.6000 146.6000 ;
	    RECT 255.0000 146.1000 255.3000 146.8000 ;
	    RECT 255.8000 146.2000 256.1000 147.9000 ;
	    RECT 258.2000 147.8000 258.5000 147.9000 ;
	    RECT 259.0000 147.8000 259.4000 148.6000 ;
	    RECT 257.6000 147.6000 258.5000 147.8000 ;
	    RECT 256.4000 147.5000 258.5000 147.6000 ;
	    RECT 256.4000 147.3000 257.9000 147.5000 ;
	    RECT 256.4000 147.2000 256.8000 147.3000 ;
	    RECT 259.9000 147.2000 260.2000 148.9000 ;
	    RECT 261.4000 147.9000 261.8000 149.9000 ;
	    RECT 262.2000 148.0000 262.6000 149.9000 ;
	    RECT 263.8000 148.0000 264.2000 149.9000 ;
	    RECT 265.4000 148.9000 265.8000 149.9000 ;
	    RECT 262.2000 147.9000 264.2000 148.0000 ;
	    RECT 261.5000 147.2000 261.8000 147.9000 ;
	    RECT 262.3000 147.7000 264.1000 147.9000 ;
	    RECT 264.6000 147.8000 265.0000 148.2000 ;
	    RECT 263.4000 147.2000 263.8000 147.4000 ;
	    RECT 255.8000 146.1000 256.2000 146.2000 ;
	    RECT 255.0000 145.8000 256.2000 146.1000 ;
	    RECT 255.8000 145.1000 256.1000 145.8000 ;
	    RECT 256.5000 145.5000 256.8000 147.2000 ;
	    RECT 257.2000 146.6000 257.8000 147.0000 ;
	    RECT 257.4000 146.2000 257.7000 146.6000 ;
	    RECT 258.2000 146.4000 258.6000 147.2000 ;
	    RECT 259.8000 147.1000 260.2000 147.2000 ;
	    RECT 259.0000 146.8000 260.2000 147.1000 ;
	    RECT 261.4000 146.8000 262.7000 147.2000 ;
	    RECT 263.4000 146.9000 264.2000 147.2000 ;
	    RECT 263.8000 146.8000 264.2000 146.9000 ;
	    RECT 264.6000 147.1000 264.9000 147.8000 ;
	    RECT 265.4000 147.2000 265.7000 148.9000 ;
	    RECT 266.2000 147.8000 266.6000 148.6000 ;
	    RECT 268.3000 148.2000 268.7000 149.9000 ;
	    RECT 267.8000 147.8000 268.9000 148.2000 ;
	    RECT 266.2000 147.2000 266.5000 147.8000 ;
	    RECT 265.4000 147.1000 265.8000 147.2000 ;
	    RECT 264.6000 146.8000 265.8000 147.1000 ;
	    RECT 266.2000 147.1000 266.6000 147.2000 ;
	    RECT 267.0000 147.1000 267.4000 147.6000 ;
	    RECT 266.2000 146.8000 267.4000 147.1000 ;
	    RECT 259.0000 146.2000 259.3000 146.8000 ;
	    RECT 257.4000 145.8000 257.8000 146.2000 ;
	    RECT 259.0000 145.8000 259.4000 146.2000 ;
	    RECT 256.5000 145.2000 257.7000 145.5000 ;
	    RECT 241.7000 141.1000 242.1000 144.7000 ;
	    RECT 245.4000 143.8000 245.8000 144.6000 ;
	    RECT 246.2000 143.5000 246.5000 144.8000 ;
	    RECT 244.7000 143.2000 246.5000 143.5000 ;
	    RECT 244.7000 143.1000 245.0000 143.2000 ;
	    RECT 244.6000 141.1000 245.0000 143.1000 ;
	    RECT 246.2000 143.1000 246.5000 143.2000 ;
	    RECT 247.3000 144.7000 248.2000 145.1000 ;
	    RECT 249.4000 144.8000 250.1000 145.1000 ;
	    RECT 250.4000 144.8000 250.9000 145.1000 ;
	    RECT 252.6000 144.8000 253.3000 145.1000 ;
	    RECT 253.6000 144.8000 254.1000 145.1000 ;
	    RECT 246.2000 141.1000 246.6000 143.1000 ;
	    RECT 247.3000 141.1000 247.7000 144.7000 ;
	    RECT 249.8000 144.2000 250.1000 144.8000 ;
	    RECT 250.5000 144.2000 250.9000 144.8000 ;
	    RECT 253.0000 144.2000 253.3000 144.8000 ;
	    RECT 249.8000 143.8000 250.2000 144.2000 ;
	    RECT 250.5000 143.8000 251.4000 144.2000 ;
	    RECT 253.0000 143.8000 253.4000 144.2000 ;
	    RECT 250.5000 141.1000 250.9000 143.8000 ;
	    RECT 253.7000 141.1000 254.1000 144.8000 ;
	    RECT 255.8000 141.1000 256.2000 145.1000 ;
	    RECT 257.4000 143.1000 257.7000 145.2000 ;
	    RECT 259.9000 145.1000 260.2000 146.8000 ;
	    RECT 262.4000 146.2000 262.7000 146.8000 ;
	    RECT 260.6000 146.1000 261.0000 146.2000 ;
	    RECT 261.4000 146.1000 261.8000 146.2000 ;
	    RECT 260.6000 145.8000 261.8000 146.1000 ;
	    RECT 262.2000 145.8000 262.7000 146.2000 ;
	    RECT 263.0000 145.8000 263.4000 146.6000 ;
	    RECT 260.6000 145.4000 261.0000 145.8000 ;
	    RECT 261.4000 145.1000 261.8000 145.2000 ;
	    RECT 262.4000 145.1000 262.7000 145.8000 ;
	    RECT 264.6000 145.4000 265.0000 146.2000 ;
	    RECT 265.4000 145.1000 265.7000 146.8000 ;
	    RECT 259.8000 144.7000 260.7000 145.1000 ;
	    RECT 261.4000 144.8000 262.1000 145.1000 ;
	    RECT 262.4000 144.8000 262.9000 145.1000 ;
	    RECT 257.4000 141.1000 257.8000 143.1000 ;
	    RECT 260.3000 141.1000 260.7000 144.7000 ;
	    RECT 261.8000 144.2000 262.1000 144.8000 ;
	    RECT 261.8000 143.8000 262.2000 144.2000 ;
	    RECT 262.5000 141.1000 262.9000 144.8000 ;
	    RECT 264.9000 144.7000 265.8000 145.1000 ;
	    RECT 264.9000 141.1000 265.3000 144.7000 ;
	    RECT 267.8000 141.1000 268.2000 147.8000 ;
	    RECT 268.6000 147.2000 268.9000 147.8000 ;
	    RECT 268.6000 146.8000 269.0000 147.2000 ;
	    RECT 268.6000 144.4000 269.0000 145.2000 ;
	    RECT 269.4000 141.1000 269.8000 149.9000 ;
	    RECT 270.2000 147.8000 270.6000 148.6000 ;
	    RECT 0.6000 137.9000 1.0000 139.9000 ;
	    RECT 0.7000 137.8000 1.0000 137.9000 ;
	    RECT 2.2000 137.9000 2.6000 139.9000 ;
	    RECT 2.2000 137.8000 2.5000 137.9000 ;
	    RECT 0.7000 137.5000 2.5000 137.8000 ;
	    RECT 0.7000 136.2000 1.0000 137.5000 ;
	    RECT 1.4000 136.4000 1.8000 137.2000 ;
	    RECT 4.1000 136.2000 4.5000 139.9000 ;
	    RECT 0.6000 135.8000 1.0000 136.2000 ;
	    RECT 0.7000 134.2000 1.0000 135.8000 ;
	    RECT 3.0000 136.1000 3.4000 136.2000 ;
	    RECT 3.8000 136.1000 4.5000 136.2000 ;
	    RECT 3.0000 135.9000 4.5000 136.1000 ;
	    RECT 3.0000 135.8000 4.1000 135.9000 ;
	    RECT 3.0000 135.4000 3.4000 135.8000 ;
	    RECT 3.8000 135.2000 4.1000 135.8000 ;
	    RECT 6.2000 135.6000 6.6000 139.9000 ;
	    RECT 7.0000 135.8000 7.4000 136.6000 ;
	    RECT 4.6000 135.4000 6.6000 135.6000 ;
	    RECT 4.5000 135.3000 6.6000 135.4000 ;
	    RECT 1.8000 134.8000 2.6000 135.2000 ;
	    RECT 3.8000 134.8000 4.2000 135.2000 ;
	    RECT 4.5000 135.0000 4.9000 135.3000 ;
	    RECT 0.7000 134.1000 1.5000 134.2000 ;
	    RECT 0.7000 133.9000 1.6000 134.1000 ;
	    RECT 1.2000 131.1000 1.6000 133.9000 ;
	    RECT 3.8000 133.1000 4.1000 134.8000 ;
	    RECT 4.5000 133.5000 4.8000 135.0000 ;
	    RECT 7.0000 133.8000 7.4000 134.2000 ;
	    RECT 4.5000 133.2000 5.7000 133.5000 ;
	    RECT 7.0000 133.2000 7.3000 133.8000 ;
	    RECT 7.8000 133.2000 8.2000 139.9000 ;
	    RECT 9.7000 136.3000 10.1000 139.9000 ;
	    RECT 9.7000 135.9000 10.6000 136.3000 ;
	    RECT 9.4000 134.8000 9.8000 135.6000 ;
	    RECT 10.2000 134.2000 10.5000 135.9000 ;
	    RECT 11.8000 135.1000 12.2000 139.9000 ;
	    RECT 14.2000 136.1000 14.6000 139.9000 ;
	    RECT 15.0000 136.8000 15.4000 137.2000 ;
	    RECT 15.0000 136.1000 15.3000 136.8000 ;
	    RECT 14.2000 135.8000 15.3000 136.1000 ;
	    RECT 12.6000 135.1000 13.0000 135.2000 ;
	    RECT 11.8000 134.8000 13.0000 135.1000 ;
	    RECT 10.2000 133.8000 10.6000 134.2000 ;
	    RECT 3.8000 131.1000 4.2000 133.1000 ;
	    RECT 5.4000 132.1000 5.7000 133.2000 ;
	    RECT 6.2000 132.4000 6.6000 133.2000 ;
	    RECT 7.0000 132.8000 8.2000 133.2000 ;
	    RECT 9.4000 133.1000 9.8000 133.2000 ;
	    RECT 10.2000 133.1000 10.5000 133.8000 ;
	    RECT 9.4000 132.8000 10.5000 133.1000 ;
	    RECT 5.4000 131.1000 5.8000 132.1000 ;
	    RECT 7.3000 131.1000 7.7000 132.8000 ;
	    RECT 10.2000 132.1000 10.5000 132.8000 ;
	    RECT 10.2000 131.1000 10.6000 132.1000 ;
	    RECT 11.8000 131.1000 12.2000 134.8000 ;
	    RECT 14.2000 131.1000 14.6000 135.8000 ;
	    RECT 15.8000 135.1000 16.2000 139.9000 ;
	    RECT 16.6000 135.8000 17.0000 136.6000 ;
	    RECT 17.4000 135.6000 17.8000 139.9000 ;
	    RECT 19.5000 136.2000 19.9000 139.9000 ;
	    RECT 21.4000 137.9000 21.8000 139.9000 ;
	    RECT 21.5000 137.8000 21.8000 137.9000 ;
	    RECT 23.0000 137.9000 23.4000 139.9000 ;
	    RECT 23.0000 137.8000 23.3000 137.9000 ;
	    RECT 21.5000 137.5000 23.3000 137.8000 ;
	    RECT 22.2000 136.4000 22.6000 137.2000 ;
	    RECT 23.0000 136.2000 23.3000 137.5000 ;
	    RECT 24.1000 136.3000 24.5000 139.9000 ;
	    RECT 19.5000 136.1000 20.2000 136.2000 ;
	    RECT 20.6000 136.1000 21.0000 136.2000 ;
	    RECT 19.5000 135.9000 21.0000 136.1000 ;
	    RECT 19.8000 135.8000 21.0000 135.9000 ;
	    RECT 17.4000 135.4000 19.4000 135.6000 ;
	    RECT 17.4000 135.3000 19.5000 135.4000 ;
	    RECT 15.8000 134.8000 16.9000 135.1000 ;
	    RECT 19.1000 135.0000 19.5000 135.3000 ;
	    RECT 19.9000 135.2000 20.2000 135.8000 ;
	    RECT 20.6000 135.4000 21.0000 135.8000 ;
	    RECT 23.0000 135.8000 23.4000 136.2000 ;
	    RECT 24.1000 135.9000 25.0000 136.3000 ;
	    RECT 26.2000 135.9000 26.6000 139.9000 ;
	    RECT 27.8000 137.9000 28.2000 139.9000 ;
	    RECT 15.8000 133.1000 16.2000 134.8000 ;
	    RECT 16.6000 134.2000 16.9000 134.8000 ;
	    RECT 16.6000 133.8000 17.0000 134.2000 ;
	    RECT 19.2000 133.5000 19.5000 135.0000 ;
	    RECT 19.8000 134.8000 20.2000 135.2000 ;
	    RECT 21.4000 134.8000 22.2000 135.2000 ;
	    RECT 23.0000 135.1000 23.3000 135.8000 ;
	    RECT 23.8000 135.1000 24.2000 135.6000 ;
	    RECT 23.0000 134.8000 24.2000 135.1000 ;
	    RECT 18.3000 133.2000 19.5000 133.5000 ;
	    RECT 15.8000 132.8000 16.7000 133.1000 ;
	    RECT 16.3000 131.1000 16.7000 132.8000 ;
	    RECT 17.4000 132.4000 17.8000 133.2000 ;
	    RECT 18.3000 132.1000 18.6000 133.2000 ;
	    RECT 19.9000 133.1000 20.2000 134.8000 ;
	    RECT 23.0000 134.2000 23.3000 134.8000 ;
	    RECT 22.5000 134.1000 23.3000 134.2000 ;
	    RECT 18.2000 131.1000 18.6000 132.1000 ;
	    RECT 19.8000 131.1000 20.2000 133.1000 ;
	    RECT 22.4000 133.9000 23.3000 134.1000 ;
	    RECT 24.6000 134.2000 24.9000 135.9000 ;
	    RECT 26.2000 135.2000 26.5000 135.9000 ;
	    RECT 27.8000 135.8000 28.1000 137.9000 ;
	    RECT 26.9000 135.5000 28.1000 135.8000 ;
	    RECT 26.2000 134.8000 26.6000 135.2000 ;
	    RECT 22.4000 131.1000 22.8000 133.9000 ;
	    RECT 24.6000 133.8000 25.0000 134.2000 ;
	    RECT 24.6000 132.2000 24.9000 133.8000 ;
	    RECT 25.4000 132.4000 25.8000 133.2000 ;
	    RECT 26.2000 133.1000 26.5000 134.8000 ;
	    RECT 26.9000 133.8000 27.2000 135.5000 ;
	    RECT 27.8000 134.8000 28.2000 135.2000 ;
	    RECT 30.2000 135.1000 30.6000 139.9000 ;
	    RECT 31.0000 135.8000 31.4000 136.6000 ;
	    RECT 33.1000 136.2000 33.5000 139.9000 ;
	    RECT 33.8000 136.8000 34.2000 137.2000 ;
	    RECT 33.9000 136.2000 34.2000 136.8000 ;
	    RECT 35.4000 136.8000 35.8000 137.2000 ;
	    RECT 35.4000 136.2000 35.7000 136.8000 ;
	    RECT 36.1000 136.2000 36.5000 139.9000 ;
	    RECT 33.1000 135.9000 33.6000 136.2000 ;
	    RECT 33.9000 135.9000 34.6000 136.2000 ;
	    RECT 32.6000 135.1000 33.0000 135.2000 ;
	    RECT 30.2000 134.8000 33.0000 135.1000 ;
	    RECT 27.8000 134.4000 28.1000 134.8000 ;
	    RECT 27.6000 134.1000 28.1000 134.4000 ;
	    RECT 27.6000 134.0000 28.0000 134.1000 ;
	    RECT 28.6000 133.8000 29.0000 134.6000 ;
	    RECT 26.8000 133.7000 27.2000 133.8000 ;
	    RECT 26.8000 133.5000 28.3000 133.7000 ;
	    RECT 26.8000 133.4000 28.9000 133.5000 ;
	    RECT 29.4000 133.4000 29.8000 134.2000 ;
	    RECT 28.0000 133.2000 28.9000 133.4000 ;
	    RECT 28.6000 133.1000 28.9000 133.2000 ;
	    RECT 30.2000 133.1000 30.6000 134.8000 ;
	    RECT 32.6000 134.4000 33.0000 134.8000 ;
	    RECT 33.3000 135.1000 33.6000 135.9000 ;
	    RECT 34.2000 135.8000 34.6000 135.9000 ;
	    RECT 35.0000 135.9000 35.7000 136.2000 ;
	    RECT 36.0000 135.9000 36.5000 136.2000 ;
	    RECT 35.0000 135.8000 35.4000 135.9000 ;
	    RECT 35.0000 135.1000 35.3000 135.8000 ;
	    RECT 36.0000 135.2000 36.3000 135.9000 ;
	    RECT 33.3000 134.8000 35.3000 135.1000 ;
	    RECT 35.8000 134.8000 36.3000 135.2000 ;
	    RECT 33.3000 134.2000 33.6000 134.8000 ;
	    RECT 36.0000 134.2000 36.3000 134.8000 ;
	    RECT 36.6000 135.1000 37.0000 135.2000 ;
	    RECT 38.2000 135.1000 38.6000 139.9000 ;
	    RECT 39.8000 135.7000 40.2000 139.9000 ;
	    RECT 42.0000 138.2000 42.4000 139.9000 ;
	    RECT 41.4000 137.9000 42.4000 138.2000 ;
	    RECT 44.2000 137.9000 44.6000 139.9000 ;
	    RECT 46.3000 137.9000 46.9000 139.9000 ;
	    RECT 41.4000 137.5000 41.8000 137.9000 ;
	    RECT 44.2000 137.6000 44.5000 137.9000 ;
	    RECT 43.1000 137.3000 44.9000 137.6000 ;
	    RECT 46.2000 137.5000 46.6000 137.9000 ;
	    RECT 43.1000 137.2000 43.5000 137.3000 ;
	    RECT 44.5000 137.2000 44.9000 137.3000 ;
	    RECT 41.4000 136.5000 41.8000 136.6000 ;
	    RECT 43.7000 136.5000 44.1000 136.6000 ;
	    RECT 41.4000 136.2000 44.1000 136.5000 ;
	    RECT 44.4000 136.5000 45.5000 136.8000 ;
	    RECT 44.4000 135.9000 44.7000 136.5000 ;
	    RECT 45.1000 136.4000 45.5000 136.5000 ;
	    RECT 46.3000 136.6000 47.0000 137.0000 ;
	    RECT 46.3000 136.1000 46.6000 136.6000 ;
	    RECT 42.3000 135.7000 44.7000 135.9000 ;
	    RECT 39.8000 135.6000 44.7000 135.7000 ;
	    RECT 45.4000 135.8000 46.6000 136.1000 ;
	    RECT 39.8000 135.5000 42.7000 135.6000 ;
	    RECT 39.8000 135.4000 42.6000 135.5000 ;
	    RECT 45.4000 135.2000 45.7000 135.8000 ;
	    RECT 48.6000 135.6000 49.0000 139.9000 ;
	    RECT 50.7000 136.3000 51.1000 139.9000 ;
	    RECT 52.6000 137.9000 53.0000 139.9000 ;
	    RECT 50.2000 135.9000 51.1000 136.3000 ;
	    RECT 50.2000 135.8000 50.6000 135.9000 ;
	    RECT 46.9000 135.3000 49.0000 135.6000 ;
	    RECT 46.9000 135.2000 47.3000 135.3000 ;
	    RECT 43.0000 135.1000 43.4000 135.2000 ;
	    RECT 36.6000 134.8000 38.6000 135.1000 ;
	    RECT 36.6000 134.4000 37.0000 134.8000 ;
	    RECT 31.8000 134.1000 32.2000 134.2000 ;
	    RECT 31.8000 133.8000 32.6000 134.1000 ;
	    RECT 33.3000 133.8000 34.6000 134.2000 ;
	    RECT 35.0000 133.8000 36.3000 134.2000 ;
	    RECT 37.4000 134.1000 37.8000 134.2000 ;
	    RECT 37.0000 133.8000 37.8000 134.1000 ;
	    RECT 32.2000 133.6000 32.6000 133.8000 ;
	    RECT 31.9000 133.1000 33.7000 133.3000 ;
	    RECT 34.2000 133.1000 34.5000 133.8000 ;
	    RECT 35.1000 133.1000 35.4000 133.8000 ;
	    RECT 37.0000 133.6000 37.4000 133.8000 ;
	    RECT 35.9000 133.1000 37.7000 133.3000 ;
	    RECT 26.2000 132.6000 26.9000 133.1000 ;
	    RECT 26.5000 132.2000 26.9000 132.6000 ;
	    RECT 24.6000 131.1000 25.0000 132.2000 ;
	    RECT 26.2000 131.8000 26.9000 132.2000 ;
	    RECT 26.5000 131.1000 26.9000 131.8000 ;
	    RECT 28.6000 131.1000 29.0000 133.1000 ;
	    RECT 30.2000 132.8000 31.1000 133.1000 ;
	    RECT 30.7000 132.2000 31.1000 132.8000 ;
	    RECT 30.2000 131.8000 31.1000 132.2000 ;
	    RECT 30.7000 131.1000 31.1000 131.8000 ;
	    RECT 31.8000 133.0000 33.8000 133.1000 ;
	    RECT 31.8000 131.1000 32.2000 133.0000 ;
	    RECT 33.4000 131.1000 33.8000 133.0000 ;
	    RECT 34.2000 131.1000 34.6000 133.1000 ;
	    RECT 35.0000 131.1000 35.4000 133.1000 ;
	    RECT 35.8000 133.0000 37.8000 133.1000 ;
	    RECT 35.8000 131.1000 36.2000 133.0000 ;
	    RECT 37.4000 131.1000 37.8000 133.0000 ;
	    RECT 38.2000 131.1000 38.6000 134.8000 ;
	    RECT 40.9000 134.8000 43.4000 135.1000 ;
	    RECT 45.4000 134.8000 45.8000 135.2000 ;
	    RECT 47.7000 134.9000 48.1000 135.0000 ;
	    RECT 40.9000 134.7000 41.3000 134.8000 ;
	    RECT 42.2000 134.7000 42.6000 134.8000 ;
	    RECT 41.7000 134.2000 42.1000 134.3000 ;
	    RECT 45.4000 134.2000 45.7000 134.8000 ;
	    RECT 46.2000 134.6000 48.1000 134.9000 ;
	    RECT 46.2000 134.5000 46.6000 134.6000 ;
	    RECT 39.0000 133.8000 39.4000 134.2000 ;
	    RECT 40.2000 133.9000 45.7000 134.2000 ;
	    RECT 40.2000 133.8000 41.0000 133.9000 ;
	    RECT 39.0000 133.2000 39.3000 133.8000 ;
	    RECT 39.0000 132.4000 39.4000 133.2000 ;
	    RECT 39.8000 131.1000 40.2000 133.5000 ;
	    RECT 42.3000 132.8000 42.6000 133.9000 ;
	    RECT 45.1000 133.8000 45.5000 133.9000 ;
	    RECT 48.6000 133.6000 49.0000 135.3000 ;
	    RECT 50.3000 134.2000 50.6000 135.8000 ;
	    RECT 52.7000 135.8000 53.0000 137.9000 ;
	    RECT 54.2000 135.9000 54.6000 139.9000 ;
	    RECT 56.3000 139.2000 57.3000 139.9000 ;
	    RECT 55.8000 138.8000 57.3000 139.2000 ;
	    RECT 56.3000 135.9000 57.3000 138.8000 ;
	    RECT 51.0000 134.8000 51.4000 135.6000 ;
	    RECT 52.7000 135.5000 53.9000 135.8000 ;
	    RECT 52.6000 134.8000 53.0000 135.2000 ;
	    RECT 50.2000 133.8000 50.6000 134.2000 ;
	    RECT 51.8000 133.8000 52.2000 134.6000 ;
	    RECT 52.7000 134.4000 53.0000 134.8000 ;
	    RECT 52.6000 134.0000 53.2000 134.4000 ;
	    RECT 53.6000 133.8000 53.9000 135.5000 ;
	    RECT 54.3000 135.2000 54.6000 135.9000 ;
	    RECT 54.2000 135.1000 54.6000 135.2000 ;
	    RECT 54.2000 134.8000 55.4000 135.1000 ;
	    RECT 47.1000 133.3000 49.0000 133.6000 ;
	    RECT 47.1000 133.2000 47.5000 133.3000 ;
	    RECT 48.6000 133.1000 49.0000 133.3000 ;
	    RECT 49.4000 133.1000 49.8000 133.2000 ;
	    RECT 48.6000 132.8000 49.8000 133.1000 ;
	    RECT 41.4000 132.1000 41.8000 132.5000 ;
	    RECT 42.2000 132.4000 42.6000 132.8000 ;
	    RECT 43.1000 132.7000 43.5000 132.8000 ;
	    RECT 43.1000 132.4000 44.5000 132.7000 ;
	    RECT 44.2000 132.1000 44.5000 132.4000 ;
	    RECT 46.2000 132.1000 46.6000 132.5000 ;
	    RECT 41.4000 131.8000 42.4000 132.1000 ;
	    RECT 42.0000 131.1000 42.4000 131.8000 ;
	    RECT 44.2000 131.1000 44.6000 132.1000 ;
	    RECT 46.2000 131.8000 46.9000 132.1000 ;
	    RECT 46.3000 131.1000 46.9000 131.8000 ;
	    RECT 48.6000 131.1000 49.0000 132.8000 ;
	    RECT 49.4000 132.4000 49.8000 132.8000 ;
	    RECT 50.3000 132.1000 50.6000 133.8000 ;
	    RECT 53.6000 133.7000 54.0000 133.8000 ;
	    RECT 52.5000 133.5000 54.0000 133.7000 ;
	    RECT 51.9000 133.4000 54.0000 133.5000 ;
	    RECT 51.9000 133.2000 52.8000 133.4000 ;
	    RECT 51.9000 133.1000 52.2000 133.2000 ;
	    RECT 54.3000 133.1000 54.6000 134.8000 ;
	    RECT 55.0000 133.8000 55.4000 134.8000 ;
	    RECT 55.8000 134.4000 56.2000 135.2000 ;
	    RECT 56.7000 134.2000 57.0000 135.9000 ;
	    RECT 57.4000 135.1000 57.8000 135.2000 ;
	    RECT 61.4000 135.1000 61.8000 139.9000 ;
	    RECT 57.4000 134.8000 61.8000 135.1000 ;
	    RECT 57.4000 134.4000 57.8000 134.8000 ;
	    RECT 56.6000 134.1000 57.0000 134.2000 ;
	    RECT 58.2000 134.1000 58.6000 134.2000 ;
	    RECT 55.8000 133.8000 57.0000 134.1000 ;
	    RECT 57.8000 133.8000 58.6000 134.1000 ;
	    RECT 55.8000 133.1000 56.1000 133.8000 ;
	    RECT 57.8000 133.6000 58.2000 133.8000 ;
	    RECT 56.7000 133.1000 58.5000 133.3000 ;
	    RECT 50.2000 131.1000 50.6000 132.1000 ;
	    RECT 51.8000 131.1000 52.2000 133.1000 ;
	    RECT 53.9000 132.6000 54.6000 133.1000 ;
	    RECT 53.9000 131.1000 54.3000 132.6000 ;
	    RECT 55.0000 131.4000 55.4000 133.1000 ;
	    RECT 55.8000 131.7000 56.2000 133.1000 ;
	    RECT 56.6000 133.0000 58.6000 133.1000 ;
	    RECT 56.6000 131.4000 57.0000 133.0000 ;
	    RECT 55.0000 131.1000 57.0000 131.4000 ;
	    RECT 58.2000 131.1000 58.6000 133.0000 ;
	    RECT 60.6000 132.4000 61.0000 133.2000 ;
	    RECT 61.4000 131.1000 61.8000 134.8000 ;
	    RECT 62.2000 135.6000 62.6000 139.9000 ;
	    RECT 64.3000 137.9000 64.9000 139.9000 ;
	    RECT 66.6000 137.9000 67.0000 139.9000 ;
	    RECT 68.8000 138.2000 69.2000 139.9000 ;
	    RECT 68.8000 137.9000 69.8000 138.2000 ;
	    RECT 64.6000 137.5000 65.0000 137.9000 ;
	    RECT 66.7000 137.6000 67.0000 137.9000 ;
	    RECT 66.3000 137.3000 68.1000 137.6000 ;
	    RECT 69.4000 137.5000 69.8000 137.9000 ;
	    RECT 66.3000 137.2000 66.7000 137.3000 ;
	    RECT 67.7000 137.2000 68.1000 137.3000 ;
	    RECT 64.2000 136.6000 64.9000 137.0000 ;
	    RECT 64.6000 136.1000 64.9000 136.6000 ;
	    RECT 65.7000 136.5000 66.8000 136.8000 ;
	    RECT 65.7000 136.4000 66.1000 136.5000 ;
	    RECT 64.6000 135.8000 65.8000 136.1000 ;
	    RECT 62.2000 135.3000 64.3000 135.6000 ;
	    RECT 62.2000 133.6000 62.6000 135.3000 ;
	    RECT 63.9000 135.2000 64.3000 135.3000 ;
	    RECT 63.1000 134.9000 63.5000 135.0000 ;
	    RECT 63.1000 134.6000 65.0000 134.9000 ;
	    RECT 64.6000 134.5000 65.0000 134.6000 ;
	    RECT 65.5000 134.2000 65.8000 135.8000 ;
	    RECT 66.5000 135.9000 66.8000 136.5000 ;
	    RECT 67.1000 136.5000 67.5000 136.6000 ;
	    RECT 69.4000 136.5000 69.8000 136.6000 ;
	    RECT 67.1000 136.2000 69.8000 136.5000 ;
	    RECT 66.5000 135.7000 68.9000 135.9000 ;
	    RECT 71.0000 135.7000 71.4000 139.9000 ;
	    RECT 72.6000 136.4000 73.0000 139.9000 ;
	    RECT 66.5000 135.6000 71.4000 135.7000 ;
	    RECT 68.5000 135.5000 71.4000 135.6000 ;
	    RECT 68.6000 135.4000 71.4000 135.5000 ;
	    RECT 72.5000 135.9000 73.0000 136.4000 ;
	    RECT 74.2000 136.2000 74.6000 139.9000 ;
	    RECT 73.3000 135.9000 74.6000 136.2000 ;
	    RECT 67.0000 135.1000 67.4000 135.2000 ;
	    RECT 67.8000 135.1000 68.2000 135.2000 ;
	    RECT 67.0000 134.8000 70.3000 135.1000 ;
	    RECT 69.9000 134.7000 70.3000 134.8000 ;
	    RECT 69.1000 134.2000 69.5000 134.3000 ;
	    RECT 72.5000 134.2000 72.8000 135.9000 ;
	    RECT 73.3000 134.9000 73.6000 135.9000 ;
	    RECT 73.1000 134.5000 73.6000 134.9000 ;
	    RECT 65.5000 133.9000 71.0000 134.2000 ;
	    RECT 65.7000 133.8000 66.1000 133.9000 ;
	    RECT 62.2000 133.3000 64.1000 133.6000 ;
	    RECT 62.2000 131.1000 62.6000 133.3000 ;
	    RECT 63.7000 133.2000 64.1000 133.3000 ;
	    RECT 68.6000 132.8000 68.9000 133.9000 ;
	    RECT 70.2000 133.8000 71.0000 133.9000 ;
	    RECT 72.5000 133.8000 73.0000 134.2000 ;
	    RECT 67.7000 132.7000 68.1000 132.8000 ;
	    RECT 64.6000 132.1000 65.0000 132.5000 ;
	    RECT 66.7000 132.4000 68.1000 132.7000 ;
	    RECT 68.6000 132.4000 69.0000 132.8000 ;
	    RECT 66.7000 132.1000 67.0000 132.4000 ;
	    RECT 69.4000 132.1000 69.8000 132.5000 ;
	    RECT 64.3000 131.8000 65.0000 132.1000 ;
	    RECT 64.3000 131.1000 64.9000 131.8000 ;
	    RECT 66.6000 131.1000 67.0000 132.1000 ;
	    RECT 68.8000 131.8000 69.8000 132.1000 ;
	    RECT 68.8000 131.1000 69.2000 131.8000 ;
	    RECT 71.0000 131.1000 71.4000 133.5000 ;
	    RECT 72.5000 133.1000 72.8000 133.8000 ;
	    RECT 73.3000 133.7000 73.6000 134.5000 ;
	    RECT 75.0000 135.6000 75.4000 139.9000 ;
	    RECT 77.1000 137.9000 77.7000 139.9000 ;
	    RECT 79.4000 137.9000 79.8000 139.9000 ;
	    RECT 81.6000 138.2000 82.0000 139.9000 ;
	    RECT 81.6000 137.9000 82.6000 138.2000 ;
	    RECT 77.4000 137.5000 77.8000 137.9000 ;
	    RECT 79.5000 137.6000 79.8000 137.9000 ;
	    RECT 79.1000 137.3000 80.9000 137.6000 ;
	    RECT 82.2000 137.5000 82.6000 137.9000 ;
	    RECT 79.1000 137.2000 79.5000 137.3000 ;
	    RECT 80.5000 137.2000 80.9000 137.3000 ;
	    RECT 76.6000 137.0000 77.3000 137.2000 ;
	    RECT 76.6000 136.8000 77.7000 137.0000 ;
	    RECT 77.0000 136.6000 77.7000 136.8000 ;
	    RECT 77.4000 136.1000 77.7000 136.6000 ;
	    RECT 78.5000 136.5000 79.6000 136.8000 ;
	    RECT 78.5000 136.4000 78.9000 136.5000 ;
	    RECT 77.4000 135.8000 78.6000 136.1000 ;
	    RECT 75.0000 135.3000 77.1000 135.6000 ;
	    RECT 73.3000 133.4000 74.6000 133.7000 ;
	    RECT 72.5000 132.8000 73.0000 133.1000 ;
	    RECT 72.6000 131.1000 73.0000 132.8000 ;
	    RECT 74.2000 131.1000 74.6000 133.4000 ;
	    RECT 75.0000 133.6000 75.4000 135.3000 ;
	    RECT 76.7000 135.2000 77.1000 135.3000 ;
	    RECT 75.9000 134.9000 76.3000 135.0000 ;
	    RECT 75.9000 134.6000 77.8000 134.9000 ;
	    RECT 77.4000 134.5000 77.8000 134.6000 ;
	    RECT 78.3000 134.2000 78.6000 135.8000 ;
	    RECT 79.3000 135.9000 79.6000 136.5000 ;
	    RECT 79.9000 136.5000 80.3000 136.6000 ;
	    RECT 82.2000 136.5000 82.6000 136.6000 ;
	    RECT 79.9000 136.2000 82.6000 136.5000 ;
	    RECT 79.3000 135.7000 81.7000 135.9000 ;
	    RECT 83.8000 135.7000 84.2000 139.9000 ;
	    RECT 85.4000 136.4000 85.8000 139.9000 ;
	    RECT 79.3000 135.6000 84.2000 135.7000 ;
	    RECT 81.3000 135.5000 84.2000 135.6000 ;
	    RECT 81.4000 135.4000 84.2000 135.5000 ;
	    RECT 85.3000 135.9000 85.8000 136.4000 ;
	    RECT 87.0000 136.2000 87.4000 139.9000 ;
	    RECT 86.1000 135.9000 87.4000 136.2000 ;
	    RECT 79.0000 135.1000 79.4000 135.2000 ;
	    RECT 80.6000 135.1000 81.0000 135.2000 ;
	    RECT 79.0000 134.8000 83.1000 135.1000 ;
	    RECT 82.7000 134.7000 83.1000 134.8000 ;
	    RECT 81.9000 134.2000 82.3000 134.3000 ;
	    RECT 85.3000 134.2000 85.6000 135.9000 ;
	    RECT 86.1000 134.9000 86.4000 135.9000 ;
	    RECT 85.9000 134.5000 86.4000 134.9000 ;
	    RECT 78.3000 133.9000 83.8000 134.2000 ;
	    RECT 78.5000 133.8000 78.9000 133.9000 ;
	    RECT 75.0000 133.3000 76.9000 133.6000 ;
	    RECT 75.0000 131.1000 75.4000 133.3000 ;
	    RECT 76.5000 133.2000 76.9000 133.3000 ;
	    RECT 81.4000 132.8000 81.7000 133.9000 ;
	    RECT 83.0000 133.8000 83.8000 133.9000 ;
	    RECT 85.3000 133.8000 85.8000 134.2000 ;
	    RECT 80.5000 132.7000 80.9000 132.8000 ;
	    RECT 77.4000 132.1000 77.8000 132.5000 ;
	    RECT 79.5000 132.4000 80.9000 132.7000 ;
	    RECT 81.4000 132.4000 81.8000 132.8000 ;
	    RECT 79.5000 132.1000 79.8000 132.4000 ;
	    RECT 82.2000 132.1000 82.6000 132.5000 ;
	    RECT 77.1000 131.8000 77.8000 132.1000 ;
	    RECT 77.1000 131.1000 77.7000 131.8000 ;
	    RECT 79.4000 131.1000 79.8000 132.1000 ;
	    RECT 81.6000 131.8000 82.6000 132.1000 ;
	    RECT 81.6000 131.1000 82.0000 131.8000 ;
	    RECT 83.8000 131.1000 84.2000 133.5000 ;
	    RECT 85.3000 133.1000 85.6000 133.8000 ;
	    RECT 86.1000 133.7000 86.4000 134.5000 ;
	    RECT 86.9000 134.8000 87.4000 135.2000 ;
	    RECT 86.9000 134.4000 87.3000 134.8000 ;
	    RECT 86.1000 133.4000 87.4000 133.7000 ;
	    RECT 85.3000 132.8000 85.8000 133.1000 ;
	    RECT 85.4000 131.1000 85.8000 132.8000 ;
	    RECT 87.0000 131.1000 87.4000 133.4000 ;
	    RECT 87.8000 132.4000 88.2000 133.2000 ;
	    RECT 88.6000 131.1000 89.0000 139.9000 ;
	    RECT 89.4000 136.2000 89.8000 139.9000 ;
	    RECT 89.4000 135.9000 90.5000 136.2000 ;
	    RECT 91.0000 135.9000 91.4000 139.9000 ;
	    RECT 90.2000 135.6000 90.5000 135.9000 ;
	    RECT 90.2000 135.2000 90.8000 135.6000 ;
	    RECT 90.2000 133.7000 90.5000 135.2000 ;
	    RECT 91.1000 134.8000 91.4000 135.9000 ;
	    RECT 92.6000 135.6000 93.0000 139.9000 ;
	    RECT 94.2000 135.6000 94.6000 139.9000 ;
	    RECT 95.8000 135.6000 96.2000 139.9000 ;
	    RECT 97.4000 135.6000 97.8000 139.9000 ;
	    RECT 89.4000 133.4000 90.5000 133.7000 ;
	    RECT 89.4000 131.1000 89.8000 133.4000 ;
	    RECT 91.0000 131.1000 91.4000 134.8000 ;
	    RECT 91.8000 135.2000 93.0000 135.6000 ;
	    RECT 93.5000 135.2000 94.6000 135.6000 ;
	    RECT 95.1000 135.2000 96.2000 135.6000 ;
	    RECT 96.9000 135.2000 97.8000 135.6000 ;
	    RECT 91.8000 133.8000 92.2000 135.2000 ;
	    RECT 93.5000 134.5000 93.9000 135.2000 ;
	    RECT 95.1000 134.5000 95.5000 135.2000 ;
	    RECT 96.9000 134.5000 97.3000 135.2000 ;
	    RECT 92.6000 134.1000 93.9000 134.5000 ;
	    RECT 94.3000 134.1000 95.5000 134.5000 ;
	    RECT 96.0000 134.1000 97.3000 134.5000 ;
	    RECT 93.5000 133.8000 93.9000 134.1000 ;
	    RECT 95.1000 133.8000 95.5000 134.1000 ;
	    RECT 96.9000 133.8000 97.3000 134.1000 ;
	    RECT 91.8000 133.4000 93.0000 133.8000 ;
	    RECT 93.5000 133.4000 94.6000 133.8000 ;
	    RECT 95.1000 133.4000 96.2000 133.8000 ;
	    RECT 96.9000 133.4000 97.8000 133.8000 ;
	    RECT 92.6000 131.1000 93.0000 133.4000 ;
	    RECT 94.2000 131.1000 94.6000 133.4000 ;
	    RECT 95.8000 131.1000 96.2000 133.4000 ;
	    RECT 97.4000 131.1000 97.8000 133.4000 ;
	    RECT 99.0000 132.4000 99.4000 133.2000 ;
	    RECT 99.8000 131.1000 100.2000 139.9000 ;
	    RECT 100.6000 133.4000 101.0000 134.2000 ;
	    RECT 101.4000 133.1000 101.8000 139.9000 ;
	    RECT 103.1000 139.6000 104.9000 139.9000 ;
	    RECT 103.1000 139.5000 103.4000 139.6000 ;
	    RECT 102.2000 135.8000 102.6000 136.6000 ;
	    RECT 103.0000 136.5000 103.4000 139.5000 ;
	    RECT 104.6000 139.5000 104.9000 139.6000 ;
	    RECT 105.4000 139.6000 107.4000 139.9000 ;
	    RECT 103.8000 136.5000 104.2000 139.3000 ;
	    RECT 104.6000 136.7000 105.0000 139.5000 ;
	    RECT 105.4000 137.0000 105.8000 139.6000 ;
	    RECT 106.2000 136.9000 106.6000 139.3000 ;
	    RECT 107.0000 136.9000 107.4000 139.6000 ;
	    RECT 106.2000 136.7000 106.5000 136.9000 ;
	    RECT 104.6000 136.5000 106.5000 136.7000 ;
	    RECT 103.9000 136.2000 104.2000 136.5000 ;
	    RECT 104.7000 136.4000 106.5000 136.5000 ;
	    RECT 107.1000 136.6000 107.4000 136.9000 ;
	    RECT 108.6000 136.9000 109.0000 139.9000 ;
	    RECT 108.6000 136.6000 108.9000 136.9000 ;
	    RECT 107.1000 136.3000 108.9000 136.6000 ;
	    RECT 111.3000 136.3000 111.7000 139.9000 ;
	    RECT 114.2000 137.9000 114.6000 139.9000 ;
	    RECT 103.8000 136.1000 104.2000 136.2000 ;
	    RECT 103.8000 135.8000 105.5000 136.1000 ;
	    RECT 111.3000 135.9000 112.2000 136.3000 ;
	    RECT 103.0000 133.1000 103.4000 133.2000 ;
	    RECT 101.4000 132.8000 103.4000 133.1000 ;
	    RECT 101.9000 131.1000 102.3000 132.8000 ;
	    RECT 105.2000 132.5000 105.5000 135.8000 ;
	    RECT 105.8000 134.8000 106.6000 135.2000 ;
	    RECT 110.2000 135.1000 110.6000 135.2000 ;
	    RECT 111.0000 135.1000 111.4000 135.6000 ;
	    RECT 110.2000 134.8000 111.4000 135.1000 ;
	    RECT 111.8000 134.2000 112.1000 135.9000 ;
	    RECT 114.3000 135.8000 114.6000 137.9000 ;
	    RECT 115.8000 135.9000 116.2000 139.9000 ;
	    RECT 116.9000 136.3000 117.3000 139.9000 ;
	    RECT 116.9000 135.9000 117.8000 136.3000 ;
	    RECT 114.3000 135.5000 115.5000 135.8000 ;
	    RECT 112.6000 135.1000 113.0000 135.2000 ;
	    RECT 112.6000 134.8000 113.8000 135.1000 ;
	    RECT 114.2000 134.8000 114.6000 135.2000 ;
	    RECT 106.6000 133.8000 107.4000 134.2000 ;
	    RECT 111.8000 133.8000 112.2000 134.2000 ;
	    RECT 113.4000 133.8000 113.8000 134.8000 ;
	    RECT 114.3000 134.4000 114.6000 134.8000 ;
	    RECT 114.2000 134.0000 114.8000 134.4000 ;
	    RECT 115.2000 133.8000 115.5000 135.5000 ;
	    RECT 115.9000 135.2000 116.2000 135.9000 ;
	    RECT 115.8000 134.8000 116.2000 135.2000 ;
	    RECT 116.6000 134.8000 117.0000 135.6000 ;
	    RECT 107.3000 132.8000 108.2000 133.2000 ;
	    RECT 111.0000 133.1000 111.4000 133.2000 ;
	    RECT 111.8000 133.1000 112.1000 133.8000 ;
	    RECT 115.2000 133.7000 115.6000 133.8000 ;
	    RECT 114.1000 133.5000 115.6000 133.7000 ;
	    RECT 113.5000 133.4000 115.6000 133.5000 ;
	    RECT 113.5000 133.2000 114.4000 133.4000 ;
	    RECT 111.0000 132.8000 112.1000 133.1000 ;
	    RECT 105.2000 132.2000 107.2000 132.5000 ;
	    RECT 105.2000 132.1000 105.8000 132.2000 ;
	    RECT 105.4000 131.1000 105.8000 132.1000 ;
	    RECT 106.9000 132.1000 107.2000 132.2000 ;
	    RECT 111.8000 132.1000 112.1000 132.8000 ;
	    RECT 112.6000 132.4000 113.0000 133.2000 ;
	    RECT 113.5000 133.1000 113.8000 133.2000 ;
	    RECT 115.9000 133.1000 116.2000 134.8000 ;
	    RECT 106.9000 131.8000 107.4000 132.1000 ;
	    RECT 107.0000 131.1000 107.4000 131.8000 ;
	    RECT 111.8000 131.1000 112.2000 132.1000 ;
	    RECT 113.4000 131.1000 113.8000 133.1000 ;
	    RECT 115.5000 132.6000 116.2000 133.1000 ;
	    RECT 117.4000 134.2000 117.7000 135.9000 ;
	    RECT 119.0000 135.6000 119.4000 139.9000 ;
	    RECT 121.1000 137.9000 121.7000 139.9000 ;
	    RECT 123.4000 137.9000 123.8000 139.9000 ;
	    RECT 125.6000 138.2000 126.0000 139.9000 ;
	    RECT 125.6000 137.9000 126.6000 138.2000 ;
	    RECT 121.4000 137.5000 121.8000 137.9000 ;
	    RECT 123.5000 137.6000 123.8000 137.9000 ;
	    RECT 123.1000 137.3000 124.9000 137.6000 ;
	    RECT 126.2000 137.5000 126.6000 137.9000 ;
	    RECT 123.1000 137.2000 123.5000 137.3000 ;
	    RECT 124.5000 137.2000 124.9000 137.3000 ;
	    RECT 121.0000 136.6000 121.7000 137.0000 ;
	    RECT 121.4000 136.1000 121.7000 136.6000 ;
	    RECT 122.5000 136.5000 123.6000 136.8000 ;
	    RECT 122.5000 136.4000 122.9000 136.5000 ;
	    RECT 121.4000 135.8000 122.6000 136.1000 ;
	    RECT 119.0000 135.3000 121.1000 135.6000 ;
	    RECT 117.4000 133.8000 117.8000 134.2000 ;
	    RECT 118.2000 133.8000 118.6000 134.2000 ;
	    RECT 115.5000 132.2000 115.9000 132.6000 ;
	    RECT 117.4000 132.2000 117.7000 133.8000 ;
	    RECT 118.2000 133.2000 118.5000 133.8000 ;
	    RECT 119.0000 133.6000 119.4000 135.3000 ;
	    RECT 120.7000 135.2000 121.1000 135.3000 ;
	    RECT 119.9000 134.9000 120.3000 135.0000 ;
	    RECT 119.9000 134.6000 121.8000 134.9000 ;
	    RECT 121.4000 134.5000 121.8000 134.6000 ;
	    RECT 122.3000 134.2000 122.6000 135.8000 ;
	    RECT 123.3000 135.9000 123.6000 136.5000 ;
	    RECT 123.9000 136.5000 124.3000 136.6000 ;
	    RECT 126.2000 136.5000 126.6000 136.6000 ;
	    RECT 123.9000 136.2000 126.6000 136.5000 ;
	    RECT 123.3000 135.7000 125.7000 135.9000 ;
	    RECT 127.8000 135.7000 128.2000 139.9000 ;
	    RECT 123.3000 135.6000 128.2000 135.7000 ;
	    RECT 125.3000 135.5000 128.2000 135.6000 ;
	    RECT 125.4000 135.4000 128.2000 135.5000 ;
	    RECT 128.6000 135.6000 129.0000 139.9000 ;
	    RECT 130.7000 137.9000 131.3000 139.9000 ;
	    RECT 133.0000 137.9000 133.4000 139.9000 ;
	    RECT 135.2000 138.2000 135.6000 139.9000 ;
	    RECT 135.2000 137.9000 136.2000 138.2000 ;
	    RECT 131.0000 137.5000 131.4000 137.9000 ;
	    RECT 133.1000 137.6000 133.4000 137.9000 ;
	    RECT 132.7000 137.3000 134.5000 137.6000 ;
	    RECT 135.8000 137.5000 136.2000 137.9000 ;
	    RECT 132.7000 137.2000 133.1000 137.3000 ;
	    RECT 134.1000 137.2000 134.5000 137.3000 ;
	    RECT 130.6000 136.6000 131.3000 137.0000 ;
	    RECT 131.0000 136.1000 131.3000 136.6000 ;
	    RECT 132.1000 136.5000 133.2000 136.8000 ;
	    RECT 132.1000 136.4000 132.5000 136.5000 ;
	    RECT 131.0000 135.8000 132.2000 136.1000 ;
	    RECT 128.6000 135.3000 130.7000 135.6000 ;
	    RECT 124.6000 135.1000 125.0000 135.2000 ;
	    RECT 124.6000 134.8000 127.1000 135.1000 ;
	    RECT 126.7000 134.7000 127.1000 134.8000 ;
	    RECT 125.9000 134.2000 126.3000 134.3000 ;
	    RECT 122.3000 133.9000 127.8000 134.2000 ;
	    RECT 122.5000 133.8000 122.9000 133.9000 ;
	    RECT 119.0000 133.3000 120.9000 133.6000 ;
	    RECT 118.2000 132.4000 118.6000 133.2000 ;
	    RECT 115.5000 131.8000 116.2000 132.2000 ;
	    RECT 115.5000 131.1000 115.9000 131.8000 ;
	    RECT 117.4000 131.1000 117.8000 132.2000 ;
	    RECT 119.0000 131.1000 119.4000 133.3000 ;
	    RECT 120.5000 133.2000 120.9000 133.3000 ;
	    RECT 125.4000 132.8000 125.7000 133.9000 ;
	    RECT 127.0000 133.8000 127.8000 133.9000 ;
	    RECT 128.6000 133.6000 129.0000 135.3000 ;
	    RECT 130.3000 135.2000 130.7000 135.3000 ;
	    RECT 129.5000 134.9000 129.9000 135.0000 ;
	    RECT 129.5000 134.6000 131.4000 134.9000 ;
	    RECT 131.0000 134.5000 131.4000 134.6000 ;
	    RECT 131.9000 134.2000 132.2000 135.8000 ;
	    RECT 132.9000 135.9000 133.2000 136.5000 ;
	    RECT 133.5000 136.5000 133.9000 136.6000 ;
	    RECT 135.8000 136.5000 136.2000 136.6000 ;
	    RECT 133.5000 136.2000 136.2000 136.5000 ;
	    RECT 132.9000 135.7000 135.3000 135.9000 ;
	    RECT 137.4000 135.7000 137.8000 139.9000 ;
	    RECT 132.9000 135.6000 137.8000 135.7000 ;
	    RECT 134.9000 135.5000 137.8000 135.6000 ;
	    RECT 135.0000 135.4000 137.8000 135.5000 ;
	    RECT 138.2000 135.6000 138.6000 139.9000 ;
	    RECT 140.3000 137.9000 140.9000 139.9000 ;
	    RECT 142.6000 137.9000 143.0000 139.9000 ;
	    RECT 144.8000 138.2000 145.2000 139.9000 ;
	    RECT 144.8000 137.9000 145.8000 138.2000 ;
	    RECT 140.6000 137.5000 141.0000 137.9000 ;
	    RECT 142.7000 137.6000 143.0000 137.9000 ;
	    RECT 142.3000 137.3000 144.1000 137.6000 ;
	    RECT 145.4000 137.5000 145.8000 137.9000 ;
	    RECT 142.3000 137.2000 142.7000 137.3000 ;
	    RECT 143.7000 137.2000 144.1000 137.3000 ;
	    RECT 140.2000 136.6000 140.9000 137.0000 ;
	    RECT 140.6000 136.1000 140.9000 136.6000 ;
	    RECT 141.7000 136.5000 142.8000 136.8000 ;
	    RECT 141.7000 136.4000 142.1000 136.5000 ;
	    RECT 140.6000 135.8000 141.8000 136.1000 ;
	    RECT 138.2000 135.3000 140.3000 135.6000 ;
	    RECT 134.2000 135.1000 134.6000 135.2000 ;
	    RECT 134.2000 134.8000 136.7000 135.1000 ;
	    RECT 136.3000 134.7000 136.7000 134.8000 ;
	    RECT 135.5000 134.2000 135.9000 134.3000 ;
	    RECT 131.9000 133.9000 137.4000 134.2000 ;
	    RECT 132.1000 133.8000 132.5000 133.9000 ;
	    RECT 124.5000 132.7000 124.9000 132.8000 ;
	    RECT 121.4000 132.1000 121.8000 132.5000 ;
	    RECT 123.5000 132.4000 124.9000 132.7000 ;
	    RECT 125.4000 132.4000 125.8000 132.8000 ;
	    RECT 123.5000 132.1000 123.8000 132.4000 ;
	    RECT 126.2000 132.1000 126.6000 132.5000 ;
	    RECT 121.1000 131.8000 121.8000 132.1000 ;
	    RECT 121.1000 131.1000 121.7000 131.8000 ;
	    RECT 123.4000 131.1000 123.8000 132.1000 ;
	    RECT 125.6000 131.8000 126.6000 132.1000 ;
	    RECT 125.6000 131.1000 126.0000 131.8000 ;
	    RECT 127.8000 131.1000 128.2000 133.5000 ;
	    RECT 128.6000 133.3000 130.5000 133.6000 ;
	    RECT 128.6000 131.1000 129.0000 133.3000 ;
	    RECT 130.1000 133.2000 130.5000 133.3000 ;
	    RECT 135.0000 133.2000 135.3000 133.9000 ;
	    RECT 136.6000 133.8000 137.4000 133.9000 ;
	    RECT 138.2000 133.6000 138.6000 135.3000 ;
	    RECT 139.9000 135.2000 140.3000 135.3000 ;
	    RECT 141.5000 135.2000 141.8000 135.8000 ;
	    RECT 142.5000 135.9000 142.8000 136.5000 ;
	    RECT 143.1000 136.5000 143.5000 136.6000 ;
	    RECT 145.4000 136.5000 145.8000 136.6000 ;
	    RECT 143.1000 136.2000 145.8000 136.5000 ;
	    RECT 142.5000 135.7000 144.9000 135.9000 ;
	    RECT 147.0000 135.7000 147.4000 139.9000 ;
	    RECT 147.8000 136.2000 148.2000 139.9000 ;
	    RECT 147.8000 135.9000 148.9000 136.2000 ;
	    RECT 149.4000 135.9000 149.8000 139.9000 ;
	    RECT 142.5000 135.6000 147.4000 135.7000 ;
	    RECT 144.5000 135.5000 147.4000 135.6000 ;
	    RECT 144.6000 135.4000 147.4000 135.5000 ;
	    RECT 148.6000 135.6000 148.9000 135.9000 ;
	    RECT 148.6000 135.2000 149.2000 135.6000 ;
	    RECT 139.1000 134.9000 139.5000 135.0000 ;
	    RECT 139.1000 134.6000 141.0000 134.9000 ;
	    RECT 141.4000 134.8000 141.8000 135.2000 ;
	    RECT 143.8000 135.1000 144.2000 135.2000 ;
	    RECT 143.8000 134.8000 146.3000 135.1000 ;
	    RECT 140.6000 134.5000 141.0000 134.6000 ;
	    RECT 141.5000 134.2000 141.8000 134.8000 ;
	    RECT 145.9000 134.7000 146.3000 134.8000 ;
	    RECT 145.1000 134.2000 145.5000 134.3000 ;
	    RECT 141.5000 133.9000 147.0000 134.2000 ;
	    RECT 141.7000 133.8000 142.1000 133.9000 ;
	    RECT 134.1000 132.7000 134.5000 132.8000 ;
	    RECT 131.0000 132.1000 131.4000 132.5000 ;
	    RECT 133.1000 132.4000 134.5000 132.7000 ;
	    RECT 135.0000 132.4000 135.4000 133.2000 ;
	    RECT 133.1000 132.1000 133.4000 132.4000 ;
	    RECT 135.8000 132.1000 136.2000 132.5000 ;
	    RECT 130.7000 131.8000 131.4000 132.1000 ;
	    RECT 130.7000 131.1000 131.3000 131.8000 ;
	    RECT 133.0000 131.1000 133.4000 132.1000 ;
	    RECT 135.2000 131.8000 136.2000 132.1000 ;
	    RECT 135.2000 131.1000 135.6000 131.8000 ;
	    RECT 137.4000 131.1000 137.8000 133.5000 ;
	    RECT 138.2000 133.3000 140.1000 133.6000 ;
	    RECT 138.2000 131.1000 138.6000 133.3000 ;
	    RECT 139.7000 133.2000 140.1000 133.3000 ;
	    RECT 144.6000 132.8000 144.9000 133.9000 ;
	    RECT 146.2000 133.8000 147.0000 133.9000 ;
	    RECT 148.6000 133.7000 148.9000 135.2000 ;
	    RECT 149.5000 134.8000 149.8000 135.9000 ;
	    RECT 143.7000 132.7000 144.1000 132.8000 ;
	    RECT 140.6000 132.1000 141.0000 132.5000 ;
	    RECT 142.7000 132.4000 144.1000 132.7000 ;
	    RECT 144.6000 132.4000 145.0000 132.8000 ;
	    RECT 142.7000 132.1000 143.0000 132.4000 ;
	    RECT 145.4000 132.1000 145.8000 132.5000 ;
	    RECT 140.3000 131.8000 141.0000 132.1000 ;
	    RECT 140.3000 131.1000 140.9000 131.8000 ;
	    RECT 142.6000 131.1000 143.0000 132.1000 ;
	    RECT 144.8000 131.8000 145.8000 132.1000 ;
	    RECT 144.8000 131.1000 145.2000 131.8000 ;
	    RECT 147.0000 131.1000 147.4000 133.5000 ;
	    RECT 147.8000 133.4000 148.9000 133.7000 ;
	    RECT 147.8000 131.1000 148.2000 133.4000 ;
	    RECT 149.4000 131.1000 149.8000 134.8000 ;
	    RECT 150.2000 135.6000 150.6000 139.9000 ;
	    RECT 152.3000 137.9000 152.9000 139.9000 ;
	    RECT 154.6000 137.9000 155.0000 139.9000 ;
	    RECT 156.8000 138.2000 157.2000 139.9000 ;
	    RECT 156.8000 137.9000 157.8000 138.2000 ;
	    RECT 152.6000 137.5000 153.0000 137.9000 ;
	    RECT 154.7000 137.6000 155.0000 137.9000 ;
	    RECT 154.3000 137.3000 156.1000 137.6000 ;
	    RECT 157.4000 137.5000 157.8000 137.9000 ;
	    RECT 154.3000 137.2000 154.7000 137.3000 ;
	    RECT 155.7000 137.2000 156.1000 137.3000 ;
	    RECT 151.8000 137.0000 152.5000 137.2000 ;
	    RECT 151.8000 136.8000 152.9000 137.0000 ;
	    RECT 152.2000 136.6000 152.9000 136.8000 ;
	    RECT 152.6000 136.1000 152.9000 136.6000 ;
	    RECT 153.7000 136.5000 154.8000 136.8000 ;
	    RECT 153.7000 136.4000 154.1000 136.5000 ;
	    RECT 152.6000 135.8000 153.8000 136.1000 ;
	    RECT 150.2000 135.3000 152.3000 135.6000 ;
	    RECT 150.2000 133.6000 150.6000 135.3000 ;
	    RECT 151.9000 135.2000 152.3000 135.3000 ;
	    RECT 151.1000 134.9000 151.5000 135.0000 ;
	    RECT 151.1000 134.6000 153.0000 134.9000 ;
	    RECT 152.6000 134.5000 153.0000 134.6000 ;
	    RECT 153.5000 134.2000 153.8000 135.8000 ;
	    RECT 154.5000 135.9000 154.8000 136.5000 ;
	    RECT 155.1000 136.5000 155.5000 136.6000 ;
	    RECT 157.4000 136.5000 157.8000 136.6000 ;
	    RECT 155.1000 136.2000 157.8000 136.5000 ;
	    RECT 154.5000 135.7000 156.9000 135.9000 ;
	    RECT 159.0000 135.7000 159.4000 139.9000 ;
	    RECT 154.5000 135.6000 159.4000 135.7000 ;
	    RECT 156.5000 135.5000 159.4000 135.6000 ;
	    RECT 156.6000 135.4000 159.4000 135.5000 ;
	    RECT 162.2000 135.6000 162.6000 139.9000 ;
	    RECT 163.8000 135.6000 164.2000 139.9000 ;
	    RECT 165.4000 135.6000 165.8000 139.9000 ;
	    RECT 167.0000 135.6000 167.4000 139.9000 ;
	    RECT 169.4000 135.6000 169.8000 139.9000 ;
	    RECT 171.0000 135.6000 171.4000 139.9000 ;
	    RECT 172.6000 135.6000 173.0000 139.9000 ;
	    RECT 174.2000 135.6000 174.6000 139.9000 ;
	    RECT 176.6000 137.9000 177.0000 139.9000 ;
	    RECT 176.7000 137.8000 177.0000 137.9000 ;
	    RECT 178.2000 137.9000 178.6000 139.9000 ;
	    RECT 178.2000 137.8000 178.5000 137.9000 ;
	    RECT 176.7000 137.5000 178.5000 137.8000 ;
	    RECT 177.4000 136.4000 177.8000 137.2000 ;
	    RECT 178.2000 136.2000 178.5000 137.5000 ;
	    RECT 179.0000 136.2000 179.4000 139.9000 ;
	    RECT 180.6000 136.4000 181.0000 139.9000 ;
	    RECT 162.2000 135.2000 163.1000 135.6000 ;
	    RECT 163.8000 135.2000 164.9000 135.6000 ;
	    RECT 165.4000 135.2000 166.5000 135.6000 ;
	    RECT 167.0000 135.2000 168.2000 135.6000 ;
	    RECT 169.4000 135.2000 170.3000 135.6000 ;
	    RECT 171.0000 135.2000 172.1000 135.6000 ;
	    RECT 172.6000 135.2000 173.7000 135.6000 ;
	    RECT 155.8000 135.1000 156.2000 135.2000 ;
	    RECT 155.8000 134.8000 158.3000 135.1000 ;
	    RECT 156.6000 134.7000 157.0000 134.8000 ;
	    RECT 157.9000 134.7000 158.3000 134.8000 ;
	    RECT 162.7000 134.5000 163.1000 135.2000 ;
	    RECT 164.5000 134.5000 164.9000 135.2000 ;
	    RECT 166.1000 134.5000 166.5000 135.2000 ;
	    RECT 157.1000 134.2000 157.5000 134.3000 ;
	    RECT 153.5000 133.9000 159.0000 134.2000 ;
	    RECT 153.7000 133.8000 154.1000 133.9000 ;
	    RECT 150.2000 133.3000 152.1000 133.6000 ;
	    RECT 150.2000 131.1000 150.6000 133.3000 ;
	    RECT 151.7000 133.2000 152.1000 133.3000 ;
	    RECT 156.6000 132.8000 156.9000 133.9000 ;
	    RECT 158.2000 133.8000 159.0000 133.9000 ;
	    RECT 162.7000 134.1000 164.0000 134.5000 ;
	    RECT 164.5000 134.1000 165.7000 134.5000 ;
	    RECT 166.1000 134.1000 167.4000 134.5000 ;
	    RECT 162.7000 133.8000 163.1000 134.1000 ;
	    RECT 164.5000 133.8000 164.9000 134.1000 ;
	    RECT 166.1000 133.8000 166.5000 134.1000 ;
	    RECT 167.8000 133.8000 168.2000 135.2000 ;
	    RECT 169.9000 134.5000 170.3000 135.2000 ;
	    RECT 171.7000 134.5000 172.1000 135.2000 ;
	    RECT 173.3000 134.5000 173.7000 135.2000 ;
	    RECT 174.2000 135.2000 175.4000 135.6000 ;
	    RECT 175.8000 135.4000 176.2000 136.2000 ;
	    RECT 178.2000 135.8000 178.6000 136.2000 ;
	    RECT 179.0000 135.9000 180.3000 136.2000 ;
	    RECT 180.6000 135.9000 181.1000 136.4000 ;
	    RECT 182.2000 136.2000 182.6000 139.9000 ;
	    RECT 183.8000 136.4000 184.2000 139.9000 ;
	    RECT 182.2000 135.9000 183.5000 136.2000 ;
	    RECT 183.8000 135.9000 184.3000 136.4000 ;
	    RECT 185.4000 136.2000 185.8000 139.9000 ;
	    RECT 187.0000 136.4000 187.4000 139.9000 ;
	    RECT 185.4000 135.9000 186.7000 136.2000 ;
	    RECT 187.0000 135.9000 187.5000 136.4000 ;
	    RECT 188.6000 136.2000 189.0000 139.9000 ;
	    RECT 190.2000 136.4000 190.6000 139.9000 ;
	    RECT 188.6000 135.9000 189.9000 136.2000 ;
	    RECT 190.2000 135.9000 190.7000 136.4000 ;
	    RECT 174.2000 134.8000 174.6000 135.2000 ;
	    RECT 169.9000 134.1000 171.2000 134.5000 ;
	    RECT 171.7000 134.1000 172.9000 134.5000 ;
	    RECT 173.3000 134.1000 174.6000 134.5000 ;
	    RECT 169.9000 133.8000 170.3000 134.1000 ;
	    RECT 171.7000 133.8000 172.1000 134.1000 ;
	    RECT 173.3000 133.8000 173.7000 134.1000 ;
	    RECT 175.0000 133.8000 175.4000 135.2000 ;
	    RECT 176.6000 134.8000 177.4000 135.2000 ;
	    RECT 178.2000 134.2000 178.5000 135.8000 ;
	    RECT 179.0000 134.8000 179.5000 135.2000 ;
	    RECT 179.1000 134.4000 179.5000 134.8000 ;
	    RECT 180.0000 134.9000 180.3000 135.9000 ;
	    RECT 180.0000 134.5000 180.5000 134.9000 ;
	    RECT 177.7000 134.1000 178.5000 134.2000 ;
	    RECT 155.7000 132.7000 156.1000 132.8000 ;
	    RECT 152.6000 132.1000 153.0000 132.5000 ;
	    RECT 154.7000 132.4000 156.1000 132.7000 ;
	    RECT 156.6000 132.4000 157.0000 132.8000 ;
	    RECT 154.7000 132.1000 155.0000 132.4000 ;
	    RECT 157.4000 132.1000 157.8000 132.5000 ;
	    RECT 152.3000 131.8000 153.0000 132.1000 ;
	    RECT 152.3000 131.1000 152.9000 131.8000 ;
	    RECT 154.6000 131.1000 155.0000 132.1000 ;
	    RECT 156.8000 131.8000 157.8000 132.1000 ;
	    RECT 156.8000 131.1000 157.2000 131.8000 ;
	    RECT 159.0000 131.1000 159.4000 133.5000 ;
	    RECT 162.2000 133.4000 163.1000 133.8000 ;
	    RECT 163.8000 133.4000 164.9000 133.8000 ;
	    RECT 165.4000 133.4000 166.5000 133.8000 ;
	    RECT 167.0000 133.4000 168.2000 133.8000 ;
	    RECT 169.4000 133.4000 170.3000 133.8000 ;
	    RECT 171.0000 133.4000 172.1000 133.8000 ;
	    RECT 172.6000 133.4000 173.7000 133.8000 ;
	    RECT 174.2000 133.4000 175.4000 133.8000 ;
	    RECT 177.6000 133.9000 178.5000 134.1000 ;
	    RECT 162.2000 131.1000 162.6000 133.4000 ;
	    RECT 163.8000 131.1000 164.2000 133.4000 ;
	    RECT 165.4000 131.1000 165.8000 133.4000 ;
	    RECT 167.0000 131.1000 167.4000 133.4000 ;
	    RECT 169.4000 131.1000 169.8000 133.4000 ;
	    RECT 171.0000 131.1000 171.4000 133.4000 ;
	    RECT 172.6000 131.1000 173.0000 133.4000 ;
	    RECT 174.2000 131.1000 174.6000 133.4000 ;
	    RECT 177.6000 131.1000 178.0000 133.9000 ;
	    RECT 180.0000 133.7000 180.3000 134.5000 ;
	    RECT 180.8000 134.2000 181.1000 135.9000 ;
	    RECT 182.2000 134.8000 182.7000 135.2000 ;
	    RECT 182.3000 134.4000 182.7000 134.8000 ;
	    RECT 183.2000 134.9000 183.5000 135.9000 ;
	    RECT 183.2000 134.5000 183.7000 134.9000 ;
	    RECT 180.6000 134.1000 181.1000 134.2000 ;
	    RECT 181.4000 134.1000 181.8000 134.2000 ;
	    RECT 180.6000 133.8000 181.8000 134.1000 ;
	    RECT 179.0000 133.4000 180.3000 133.7000 ;
	    RECT 179.0000 131.1000 179.4000 133.4000 ;
	    RECT 180.8000 133.1000 181.1000 133.8000 ;
	    RECT 183.2000 133.7000 183.5000 134.5000 ;
	    RECT 184.0000 134.2000 184.3000 135.9000 ;
	    RECT 185.4000 134.8000 185.9000 135.2000 ;
	    RECT 185.5000 134.4000 185.9000 134.8000 ;
	    RECT 186.4000 134.9000 186.7000 135.9000 ;
	    RECT 186.4000 134.5000 186.9000 134.9000 ;
	    RECT 183.8000 133.8000 184.3000 134.2000 ;
	    RECT 180.6000 132.8000 181.1000 133.1000 ;
	    RECT 182.2000 133.4000 183.5000 133.7000 ;
	    RECT 180.6000 131.1000 181.0000 132.8000 ;
	    RECT 182.2000 131.1000 182.6000 133.4000 ;
	    RECT 184.0000 133.1000 184.3000 133.8000 ;
	    RECT 186.4000 133.7000 186.7000 134.5000 ;
	    RECT 187.2000 134.2000 187.5000 135.9000 ;
	    RECT 188.6000 134.8000 189.1000 135.2000 ;
	    RECT 188.7000 134.4000 189.1000 134.8000 ;
	    RECT 189.6000 134.9000 189.9000 135.9000 ;
	    RECT 189.6000 134.5000 190.1000 134.9000 ;
	    RECT 187.0000 133.8000 187.5000 134.2000 ;
	    RECT 183.8000 132.8000 184.3000 133.1000 ;
	    RECT 185.4000 133.4000 186.7000 133.7000 ;
	    RECT 183.8000 131.1000 184.2000 132.8000 ;
	    RECT 185.4000 131.1000 185.8000 133.4000 ;
	    RECT 187.2000 133.1000 187.5000 133.8000 ;
	    RECT 189.6000 133.7000 189.9000 134.5000 ;
	    RECT 190.4000 134.2000 190.7000 135.9000 ;
	    RECT 190.2000 133.8000 190.7000 134.2000 ;
	    RECT 187.0000 132.8000 187.5000 133.1000 ;
	    RECT 188.6000 133.4000 189.9000 133.7000 ;
	    RECT 187.0000 131.1000 187.4000 132.8000 ;
	    RECT 188.6000 131.1000 189.0000 133.4000 ;
	    RECT 190.4000 133.1000 190.7000 133.8000 ;
	    RECT 190.2000 132.8000 190.7000 133.1000 ;
	    RECT 192.6000 135.1000 193.0000 139.9000 ;
	    RECT 195.5000 138.2000 195.9000 139.9000 ;
	    RECT 195.5000 137.8000 196.2000 138.2000 ;
	    RECT 197.4000 137.9000 197.8000 139.9000 ;
	    RECT 197.5000 137.8000 197.8000 137.9000 ;
	    RECT 199.0000 137.9000 199.4000 139.9000 ;
	    RECT 199.0000 137.8000 199.3000 137.9000 ;
	    RECT 195.5000 136.3000 195.9000 137.8000 ;
	    RECT 197.5000 137.5000 199.3000 137.8000 ;
	    RECT 198.2000 136.4000 198.6000 137.2000 ;
	    RECT 195.0000 135.9000 195.9000 136.3000 ;
	    RECT 199.0000 136.2000 199.3000 137.5000 ;
	    RECT 199.8000 137.1000 200.2000 139.9000 ;
	    RECT 200.6000 137.1000 201.0000 137.2000 ;
	    RECT 199.8000 136.8000 201.0000 137.1000 ;
	    RECT 194.2000 135.1000 194.6000 135.2000 ;
	    RECT 192.6000 134.8000 194.6000 135.1000 ;
	    RECT 190.2000 131.1000 190.6000 132.8000 ;
	    RECT 192.6000 131.1000 193.0000 134.8000 ;
	    RECT 195.1000 134.2000 195.4000 135.9000 ;
	    RECT 195.8000 134.8000 196.2000 135.6000 ;
	    RECT 196.6000 135.4000 197.0000 136.2000 ;
	    RECT 199.0000 135.8000 199.4000 136.2000 ;
	    RECT 197.4000 134.8000 198.2000 135.2000 ;
	    RECT 199.0000 134.2000 199.3000 135.8000 ;
	    RECT 193.4000 133.4000 193.8000 134.2000 ;
	    RECT 195.0000 133.8000 195.4000 134.2000 ;
	    RECT 198.2000 133.9000 199.3000 134.2000 ;
	    RECT 198.2000 133.8000 198.8000 133.9000 ;
	    RECT 194.2000 132.4000 194.6000 133.2000 ;
	    RECT 195.1000 132.1000 195.4000 133.8000 ;
	    RECT 195.0000 131.1000 195.4000 132.1000 ;
	    RECT 198.4000 131.1000 198.8000 133.8000 ;
	    RECT 199.8000 131.1000 200.2000 136.8000 ;
	    RECT 201.4000 135.8000 201.8000 136.6000 ;
	    RECT 200.6000 132.4000 201.0000 133.2000 ;
	    RECT 202.2000 133.1000 202.6000 139.9000 ;
	    RECT 204.6000 135.1000 205.0000 139.9000 ;
	    RECT 205.7000 136.3000 206.1000 139.9000 ;
	    RECT 208.2000 136.8000 208.6000 137.2000 ;
	    RECT 205.7000 135.9000 206.6000 136.3000 ;
	    RECT 208.2000 136.2000 208.5000 136.8000 ;
	    RECT 208.9000 136.2000 209.3000 139.9000 ;
	    RECT 206.2000 135.8000 206.6000 135.9000 ;
	    RECT 207.8000 135.9000 208.5000 136.2000 ;
	    RECT 208.8000 135.9000 209.3000 136.2000 ;
	    RECT 212.6000 135.9000 213.0000 139.9000 ;
	    RECT 213.4000 136.2000 213.8000 139.9000 ;
	    RECT 215.0000 136.2000 215.4000 139.9000 ;
	    RECT 213.4000 135.9000 215.4000 136.2000 ;
	    RECT 207.8000 135.8000 208.2000 135.9000 ;
	    RECT 205.4000 135.1000 205.8000 135.6000 ;
	    RECT 204.6000 134.8000 205.8000 135.1000 ;
	    RECT 201.7000 132.8000 202.6000 133.1000 ;
	    RECT 201.7000 131.1000 202.1000 132.8000 ;
	    RECT 203.8000 132.4000 204.2000 133.2000 ;
	    RECT 204.6000 133.1000 205.0000 134.8000 ;
	    RECT 206.2000 134.2000 206.5000 135.8000 ;
	    RECT 208.8000 134.2000 209.1000 135.9000 ;
	    RECT 212.7000 135.2000 213.0000 135.9000 ;
	    RECT 214.6000 135.2000 215.0000 135.4000 ;
	    RECT 209.4000 134.4000 209.8000 135.2000 ;
	    RECT 212.6000 134.9000 213.8000 135.2000 ;
	    RECT 214.6000 134.9000 215.4000 135.2000 ;
	    RECT 212.6000 134.8000 213.0000 134.9000 ;
	    RECT 206.2000 133.8000 206.6000 134.2000 ;
	    RECT 207.8000 133.8000 209.1000 134.2000 ;
	    RECT 210.2000 134.1000 210.6000 134.2000 ;
	    RECT 209.8000 133.8000 210.6000 134.1000 ;
	    RECT 205.4000 133.1000 205.8000 133.2000 ;
	    RECT 204.6000 132.8000 205.8000 133.1000 ;
	    RECT 204.6000 131.1000 205.0000 132.8000 ;
	    RECT 206.2000 132.1000 206.5000 133.8000 ;
	    RECT 207.0000 132.4000 207.4000 133.2000 ;
	    RECT 207.9000 133.1000 208.2000 133.8000 ;
	    RECT 209.8000 133.6000 210.2000 133.8000 ;
	    RECT 208.7000 133.1000 210.5000 133.3000 ;
	    RECT 206.2000 131.1000 206.6000 132.1000 ;
	    RECT 207.8000 131.1000 208.2000 133.1000 ;
	    RECT 208.6000 133.0000 210.6000 133.1000 ;
	    RECT 208.6000 131.1000 209.0000 133.0000 ;
	    RECT 210.2000 131.1000 210.6000 133.0000 ;
	    RECT 212.6000 132.8000 213.0000 133.2000 ;
	    RECT 213.5000 133.1000 213.8000 134.9000 ;
	    RECT 215.0000 134.8000 215.4000 134.9000 ;
	    RECT 214.2000 133.8000 214.6000 134.6000 ;
	    RECT 215.8000 133.4000 216.2000 134.2000 ;
	    RECT 212.7000 132.4000 213.1000 132.8000 ;
	    RECT 213.4000 131.1000 213.8000 133.1000 ;
	    RECT 216.6000 133.1000 217.0000 139.9000 ;
	    RECT 217.4000 135.8000 217.8000 136.6000 ;
	    RECT 218.2000 133.4000 218.6000 134.2000 ;
	    RECT 219.0000 133.1000 219.4000 139.9000 ;
	    RECT 219.8000 135.8000 220.2000 136.6000 ;
	    RECT 220.6000 135.1000 221.0000 135.2000 ;
	    RECT 221.4000 135.1000 221.8000 139.9000 ;
	    RECT 222.2000 135.8000 222.6000 136.6000 ;
	    RECT 220.6000 134.8000 221.8000 135.1000 ;
	    RECT 219.8000 134.1000 220.2000 134.2000 ;
	    RECT 220.6000 134.1000 221.0000 134.2000 ;
	    RECT 219.8000 133.8000 221.0000 134.1000 ;
	    RECT 220.6000 133.4000 221.0000 133.8000 ;
	    RECT 221.4000 133.1000 221.8000 134.8000 ;
	    RECT 216.6000 132.8000 217.5000 133.1000 ;
	    RECT 219.0000 132.8000 219.9000 133.1000 ;
	    RECT 221.4000 132.8000 222.3000 133.1000 ;
	    RECT 217.1000 131.1000 217.5000 132.8000 ;
	    RECT 219.5000 131.1000 219.9000 132.8000 ;
	    RECT 221.9000 131.1000 222.3000 132.8000 ;
	    RECT 223.0000 131.1000 223.4000 139.9000 ;
	    RECT 224.6000 133.4000 225.0000 134.2000 ;
	    RECT 223.8000 132.4000 224.2000 133.2000 ;
	    RECT 225.4000 133.1000 225.8000 139.9000 ;
	    RECT 226.2000 136.1000 226.6000 136.6000 ;
	    RECT 227.0000 136.1000 227.4000 136.2000 ;
	    RECT 226.2000 135.8000 227.4000 136.1000 ;
	    RECT 227.0000 133.4000 227.4000 134.2000 ;
	    RECT 227.8000 133.1000 228.2000 139.9000 ;
	    RECT 228.6000 135.8000 229.0000 136.6000 ;
	    RECT 228.6000 134.1000 229.0000 134.2000 ;
	    RECT 229.4000 134.1000 229.8000 134.2000 ;
	    RECT 228.6000 133.8000 229.8000 134.1000 ;
	    RECT 229.4000 133.4000 229.8000 133.8000 ;
	    RECT 230.2000 133.1000 230.6000 139.9000 ;
	    RECT 231.0000 135.8000 231.4000 136.6000 ;
	    RECT 231.8000 136.1000 232.2000 136.2000 ;
	    RECT 232.6000 136.1000 233.0000 139.9000 ;
	    RECT 234.2000 137.1000 234.6000 137.2000 ;
	    RECT 235.0000 137.1000 235.4000 139.9000 ;
	    RECT 234.2000 136.8000 235.4000 137.1000 ;
	    RECT 231.8000 135.8000 233.0000 136.1000 ;
	    RECT 233.4000 135.8000 233.8000 136.6000 ;
	    RECT 231.8000 133.4000 232.2000 134.2000 ;
	    RECT 232.6000 133.1000 233.0000 135.8000 ;
	    RECT 233.4000 134.1000 233.8000 134.2000 ;
	    RECT 234.2000 134.1000 234.6000 134.2000 ;
	    RECT 233.4000 133.8000 234.6000 134.1000 ;
	    RECT 234.2000 133.4000 234.6000 133.8000 ;
	    RECT 235.0000 133.1000 235.4000 136.8000 ;
	    RECT 237.9000 138.2000 238.3000 139.9000 ;
	    RECT 237.9000 137.8000 238.6000 138.2000 ;
	    RECT 235.8000 135.8000 236.2000 136.6000 ;
	    RECT 237.9000 136.3000 238.3000 137.8000 ;
	    RECT 240.3000 136.3000 240.7000 139.9000 ;
	    RECT 237.4000 135.9000 238.3000 136.3000 ;
	    RECT 239.8000 135.9000 240.7000 136.3000 ;
	    RECT 241.7000 136.3000 242.1000 139.9000 ;
	    RECT 244.2000 136.8000 244.6000 137.2000 ;
	    RECT 241.7000 135.9000 242.6000 136.3000 ;
	    RECT 244.2000 136.2000 244.5000 136.8000 ;
	    RECT 244.9000 136.2000 245.3000 139.9000 ;
	    RECT 248.3000 136.2000 248.7000 139.9000 ;
	    RECT 249.0000 136.8000 249.4000 137.2000 ;
	    RECT 249.1000 136.2000 249.4000 136.8000 ;
	    RECT 243.8000 135.9000 244.5000 136.2000 ;
	    RECT 237.5000 134.2000 237.8000 135.9000 ;
	    RECT 238.2000 134.8000 238.6000 135.6000 ;
	    RECT 239.9000 134.2000 240.2000 135.9000 ;
	    RECT 240.6000 134.8000 241.0000 135.6000 ;
	    RECT 241.4000 134.8000 241.8000 135.6000 ;
	    RECT 242.2000 135.1000 242.5000 135.9000 ;
	    RECT 243.8000 135.8000 244.2000 135.9000 ;
	    RECT 244.8000 135.8000 245.8000 136.2000 ;
	    RECT 248.3000 135.9000 248.8000 136.2000 ;
	    RECT 249.1000 135.9000 249.8000 136.2000 ;
	    RECT 251.5000 135.9000 252.5000 139.9000 ;
	    RECT 255.5000 139.2000 255.9000 139.9000 ;
	    RECT 255.0000 138.8000 255.9000 139.2000 ;
	    RECT 255.5000 136.2000 255.9000 138.8000 ;
	    RECT 258.5000 137.2000 258.9000 139.9000 ;
	    RECT 256.2000 136.8000 256.6000 137.2000 ;
	    RECT 256.3000 136.2000 256.6000 136.8000 ;
	    RECT 257.8000 136.8000 258.2000 137.2000 ;
	    RECT 258.5000 136.8000 259.4000 137.2000 ;
	    RECT 257.8000 136.2000 258.1000 136.8000 ;
	    RECT 258.5000 136.2000 258.9000 136.8000 ;
	    RECT 255.5000 135.9000 256.0000 136.2000 ;
	    RECT 256.3000 135.9000 257.0000 136.2000 ;
	    RECT 243.8000 135.1000 244.1000 135.8000 ;
	    RECT 242.2000 134.8000 244.1000 135.1000 ;
	    RECT 237.4000 133.8000 237.8000 134.2000 ;
	    RECT 239.8000 133.8000 240.2000 134.2000 ;
	    RECT 225.4000 132.8000 226.3000 133.1000 ;
	    RECT 227.8000 132.8000 228.7000 133.1000 ;
	    RECT 230.2000 132.8000 231.1000 133.1000 ;
	    RECT 232.6000 132.8000 233.5000 133.1000 ;
	    RECT 235.0000 132.8000 235.9000 133.1000 ;
	    RECT 225.9000 132.2000 226.3000 132.8000 ;
	    RECT 228.3000 132.2000 228.7000 132.8000 ;
	    RECT 230.7000 132.2000 231.1000 132.8000 ;
	    RECT 225.9000 131.8000 226.6000 132.2000 ;
	    RECT 227.8000 131.8000 228.7000 132.2000 ;
	    RECT 230.2000 131.8000 231.1000 132.2000 ;
	    RECT 225.9000 131.1000 226.3000 131.8000 ;
	    RECT 228.3000 131.1000 228.7000 131.8000 ;
	    RECT 230.7000 131.1000 231.1000 131.8000 ;
	    RECT 233.1000 131.1000 233.5000 132.8000 ;
	    RECT 235.5000 131.1000 235.9000 132.8000 ;
	    RECT 236.6000 132.4000 237.0000 133.2000 ;
	    RECT 237.5000 132.1000 237.8000 133.8000 ;
	    RECT 239.0000 132.4000 239.4000 133.2000 ;
	    RECT 239.9000 132.2000 240.2000 133.8000 ;
	    RECT 237.4000 131.1000 237.8000 132.1000 ;
	    RECT 239.8000 131.1000 240.2000 132.2000 ;
	    RECT 242.2000 134.2000 242.5000 134.8000 ;
	    RECT 244.8000 134.2000 245.1000 135.8000 ;
	    RECT 245.4000 134.4000 245.8000 135.2000 ;
	    RECT 247.8000 134.4000 248.2000 135.2000 ;
	    RECT 248.5000 135.1000 248.8000 135.9000 ;
	    RECT 249.4000 135.8000 249.8000 135.9000 ;
	    RECT 249.4000 135.1000 249.8000 135.2000 ;
	    RECT 248.5000 134.8000 249.8000 135.1000 ;
	    RECT 248.5000 134.2000 248.8000 134.8000 ;
	    RECT 251.0000 134.4000 251.4000 135.2000 ;
	    RECT 251.8000 134.2000 252.1000 135.9000 ;
	    RECT 252.6000 134.4000 253.0000 135.2000 ;
	    RECT 242.2000 133.8000 242.6000 134.2000 ;
	    RECT 243.8000 133.8000 245.1000 134.2000 ;
	    RECT 247.0000 134.1000 247.4000 134.2000 ;
	    RECT 247.0000 133.8000 247.8000 134.1000 ;
	    RECT 248.5000 133.8000 249.8000 134.2000 ;
	    RECT 250.2000 134.1000 250.6000 134.2000 ;
	    RECT 251.8000 134.1000 252.2000 134.2000 ;
	    RECT 250.2000 133.8000 251.0000 134.1000 ;
	    RECT 251.8000 133.8000 253.0000 134.1000 ;
	    RECT 253.4000 133.8000 253.8000 134.6000 ;
	    RECT 255.0000 134.4000 255.4000 135.2000 ;
	    RECT 255.7000 134.2000 256.0000 135.9000 ;
	    RECT 256.6000 135.8000 257.0000 135.9000 ;
	    RECT 257.4000 135.9000 258.1000 136.2000 ;
	    RECT 258.4000 135.9000 258.9000 136.2000 ;
	    RECT 260.9000 136.3000 261.3000 139.9000 ;
	    RECT 260.9000 135.9000 261.8000 136.3000 ;
	    RECT 263.0000 135.9000 263.4000 139.9000 ;
	    RECT 264.6000 137.9000 265.0000 139.9000 ;
	    RECT 257.4000 135.8000 257.8000 135.9000 ;
	    RECT 258.4000 134.2000 258.7000 135.9000 ;
	    RECT 259.0000 134.4000 259.4000 135.2000 ;
	    RECT 260.6000 134.8000 261.0000 135.6000 ;
	    RECT 261.4000 134.2000 261.7000 135.9000 ;
	    RECT 263.0000 135.2000 263.3000 135.9000 ;
	    RECT 264.6000 135.8000 264.9000 137.9000 ;
	    RECT 266.2000 136.2000 266.6000 139.9000 ;
	    RECT 267.8000 136.4000 268.2000 139.9000 ;
	    RECT 266.2000 135.9000 267.5000 136.2000 ;
	    RECT 267.8000 135.9000 268.3000 136.4000 ;
	    RECT 263.7000 135.5000 264.9000 135.8000 ;
	    RECT 262.2000 135.1000 262.6000 135.2000 ;
	    RECT 263.0000 135.1000 263.4000 135.2000 ;
	    RECT 262.2000 134.8000 263.4000 135.1000 ;
	    RECT 254.2000 134.1000 254.6000 134.2000 ;
	    RECT 254.2000 133.8000 255.0000 134.1000 ;
	    RECT 255.7000 133.8000 257.0000 134.2000 ;
	    RECT 257.4000 133.8000 258.7000 134.2000 ;
	    RECT 259.8000 134.1000 260.2000 134.2000 ;
	    RECT 259.4000 133.8000 260.2000 134.1000 ;
	    RECT 260.6000 133.8000 261.0000 134.2000 ;
	    RECT 261.4000 133.8000 261.8000 134.2000 ;
	    RECT 242.2000 132.1000 242.5000 133.8000 ;
	    RECT 243.0000 132.4000 243.4000 133.2000 ;
	    RECT 243.9000 133.1000 244.2000 133.8000 ;
	    RECT 247.4000 133.6000 247.8000 133.8000 ;
	    RECT 244.7000 133.1000 246.5000 133.3000 ;
	    RECT 247.1000 133.1000 248.9000 133.3000 ;
	    RECT 249.4000 133.1000 249.7000 133.8000 ;
	    RECT 250.6000 133.6000 251.0000 133.8000 ;
	    RECT 250.3000 133.1000 252.1000 133.3000 ;
	    RECT 252.7000 133.2000 253.0000 133.8000 ;
	    RECT 254.6000 133.6000 255.0000 133.8000 ;
	    RECT 242.2000 131.1000 242.6000 132.1000 ;
	    RECT 243.8000 131.1000 244.2000 133.1000 ;
	    RECT 244.6000 133.0000 246.6000 133.1000 ;
	    RECT 244.6000 131.1000 245.0000 133.0000 ;
	    RECT 246.2000 131.1000 246.6000 133.0000 ;
	    RECT 247.0000 133.0000 249.0000 133.1000 ;
	    RECT 247.0000 131.1000 247.4000 133.0000 ;
	    RECT 248.6000 131.1000 249.0000 133.0000 ;
	    RECT 249.4000 131.1000 249.8000 133.1000 ;
	    RECT 250.2000 133.0000 252.2000 133.1000 ;
	    RECT 250.2000 131.1000 250.6000 133.0000 ;
	    RECT 251.8000 131.4000 252.2000 133.0000 ;
	    RECT 252.6000 131.7000 253.0000 133.2000 ;
	    RECT 254.3000 133.1000 256.1000 133.3000 ;
	    RECT 256.6000 133.1000 256.9000 133.8000 ;
	    RECT 257.5000 133.1000 257.8000 133.8000 ;
	    RECT 259.4000 133.6000 259.8000 133.8000 ;
	    RECT 258.3000 133.1000 260.1000 133.3000 ;
	    RECT 260.6000 133.1000 260.9000 133.8000 ;
	    RECT 261.4000 133.1000 261.7000 133.8000 ;
	    RECT 253.4000 131.4000 253.8000 133.1000 ;
	    RECT 251.8000 131.1000 253.8000 131.4000 ;
	    RECT 254.2000 133.0000 256.2000 133.1000 ;
	    RECT 254.2000 131.1000 254.6000 133.0000 ;
	    RECT 255.8000 131.1000 256.2000 133.0000 ;
	    RECT 256.6000 131.1000 257.0000 133.1000 ;
	    RECT 257.4000 131.1000 257.8000 133.1000 ;
	    RECT 258.2000 133.0000 260.2000 133.1000 ;
	    RECT 258.2000 131.1000 258.6000 133.0000 ;
	    RECT 259.8000 131.1000 260.2000 133.0000 ;
	    RECT 260.6000 132.8000 261.7000 133.1000 ;
	    RECT 261.4000 132.1000 261.7000 132.8000 ;
	    RECT 263.0000 133.1000 263.3000 134.8000 ;
	    RECT 263.7000 133.8000 264.0000 135.5000 ;
	    RECT 266.2000 134.8000 266.7000 135.2000 ;
	    RECT 265.4000 133.8000 265.8000 134.6000 ;
	    RECT 266.3000 134.4000 266.7000 134.8000 ;
	    RECT 267.2000 134.9000 267.5000 135.9000 ;
	    RECT 267.2000 134.5000 267.7000 134.9000 ;
	    RECT 263.6000 133.7000 264.0000 133.8000 ;
	    RECT 267.2000 133.7000 267.5000 134.5000 ;
	    RECT 268.0000 134.2000 268.3000 135.9000 ;
	    RECT 267.8000 134.1000 268.3000 134.2000 ;
	    RECT 268.6000 134.1000 269.0000 134.2000 ;
	    RECT 267.8000 133.8000 269.0000 134.1000 ;
	    RECT 263.6000 133.5000 265.1000 133.7000 ;
	    RECT 263.6000 133.4000 265.7000 133.5000 ;
	    RECT 264.8000 133.2000 265.7000 133.4000 ;
	    RECT 265.4000 133.1000 265.7000 133.2000 ;
	    RECT 266.2000 133.4000 267.5000 133.7000 ;
	    RECT 263.0000 132.6000 263.7000 133.1000 ;
	    RECT 261.4000 131.1000 261.8000 132.1000 ;
	    RECT 263.3000 131.1000 263.7000 132.6000 ;
	    RECT 265.4000 131.1000 265.8000 133.1000 ;
	    RECT 266.2000 131.1000 266.6000 133.4000 ;
	    RECT 268.0000 133.1000 268.3000 133.8000 ;
	    RECT 267.8000 132.8000 268.3000 133.1000 ;
	    RECT 267.8000 131.1000 268.2000 132.8000 ;
	    RECT 0.6000 127.9000 1.0000 129.9000 ;
	    RECT 2.8000 129.2000 3.6000 129.9000 ;
	    RECT 2.8000 128.8000 4.2000 129.2000 ;
	    RECT 2.8000 128.1000 3.6000 128.8000 ;
	    RECT 0.6000 127.6000 1.7000 127.9000 ;
	    RECT 1.3000 127.5000 1.7000 127.6000 ;
	    RECT 2.6000 126.7000 3.0000 127.1000 ;
	    RECT 2.6000 126.4000 2.9000 126.7000 ;
	    RECT 1.6000 126.1000 2.9000 126.4000 ;
	    RECT 3.3000 126.4000 3.6000 128.1000 ;
	    RECT 5.4000 127.9000 5.8000 129.9000 ;
	    RECT 4.6000 127.6000 5.8000 127.9000 ;
	    RECT 7.8000 127.9000 8.2000 129.9000 ;
	    RECT 10.2000 128.9000 10.6000 129.9000 ;
	    RECT 8.5000 128.2000 8.9000 128.6000 ;
	    RECT 4.6000 127.5000 5.0000 127.6000 ;
	    RECT 7.0000 126.4000 7.4000 127.2000 ;
	    RECT 3.3000 126.2000 3.8000 126.4000 ;
	    RECT 3.3000 126.1000 4.2000 126.2000 ;
	    RECT 1.6000 126.0000 2.0000 126.1000 ;
	    RECT 3.5000 125.8000 4.2000 126.1000 ;
	    RECT 6.2000 126.1000 6.6000 126.2000 ;
	    RECT 7.8000 126.1000 8.1000 127.9000 ;
	    RECT 8.6000 127.8000 9.0000 128.2000 ;
	    RECT 8.6000 127.1000 8.9000 127.8000 ;
	    RECT 10.3000 127.2000 10.6000 128.9000 ;
	    RECT 10.2000 127.1000 10.6000 127.2000 ;
	    RECT 8.6000 126.8000 10.6000 127.1000 ;
	    RECT 8.6000 126.1000 9.0000 126.2000 ;
	    RECT 6.2000 125.8000 7.0000 126.1000 ;
	    RECT 7.8000 125.8000 9.0000 126.1000 ;
	    RECT 2.7000 125.7000 3.1000 125.8000 ;
	    RECT 1.4000 125.4000 3.1000 125.7000 ;
	    RECT 1.4000 125.1000 1.7000 125.4000 ;
	    RECT 3.5000 125.1000 3.8000 125.8000 ;
	    RECT 6.6000 125.6000 7.0000 125.8000 ;
	    RECT 8.6000 125.1000 8.9000 125.8000 ;
	    RECT 10.3000 125.1000 10.6000 126.8000 ;
	    RECT 11.0000 126.1000 11.4000 126.2000 ;
	    RECT 11.8000 126.1000 12.2000 129.9000 ;
	    RECT 13.4000 127.9000 13.8000 129.9000 ;
	    RECT 15.6000 128.1000 16.4000 129.9000 ;
	    RECT 13.4000 127.6000 14.5000 127.9000 ;
	    RECT 14.1000 127.5000 14.5000 127.6000 ;
	    RECT 15.4000 126.7000 15.8000 127.1000 ;
	    RECT 15.4000 126.4000 15.7000 126.7000 ;
	    RECT 11.0000 125.8000 12.2000 126.1000 ;
	    RECT 14.4000 126.1000 15.7000 126.4000 ;
	    RECT 16.1000 126.4000 16.4000 128.1000 ;
	    RECT 18.2000 127.9000 18.6000 129.9000 ;
	    RECT 17.4000 127.6000 18.6000 127.9000 ;
	    RECT 19.8000 128.9000 20.2000 129.9000 ;
	    RECT 17.4000 127.5000 17.8000 127.6000 ;
	    RECT 19.8000 127.2000 20.1000 128.9000 ;
	    RECT 23.0000 127.9000 23.4000 129.9000 ;
	    RECT 23.7000 128.2000 24.1000 128.6000 ;
	    RECT 19.8000 126.8000 20.2000 127.2000 ;
	    RECT 21.4000 127.1000 21.8000 127.2000 ;
	    RECT 22.2000 127.1000 22.6000 127.2000 ;
	    RECT 21.4000 126.8000 22.6000 127.1000 ;
	    RECT 16.1000 126.2000 16.6000 126.4000 ;
	    RECT 16.1000 126.1000 17.0000 126.2000 ;
	    RECT 14.4000 126.0000 14.8000 126.1000 ;
	    RECT 16.3000 125.8000 17.0000 126.1000 ;
	    RECT 11.0000 125.4000 11.4000 125.8000 ;
	    RECT 0.6000 124.8000 1.7000 125.1000 ;
	    RECT 0.6000 121.1000 1.0000 124.8000 ;
	    RECT 1.3000 124.7000 1.7000 124.8000 ;
	    RECT 2.8000 124.8000 3.8000 125.1000 ;
	    RECT 4.6000 124.8000 5.8000 125.1000 ;
	    RECT 2.8000 121.1000 3.6000 124.8000 ;
	    RECT 4.6000 124.7000 5.0000 124.8000 ;
	    RECT 5.4000 121.1000 5.8000 124.8000 ;
	    RECT 6.2000 124.8000 8.2000 125.1000 ;
	    RECT 6.2000 121.1000 6.6000 124.8000 ;
	    RECT 7.8000 121.1000 8.2000 124.8000 ;
	    RECT 8.6000 121.1000 9.0000 125.1000 ;
	    RECT 10.2000 124.7000 11.1000 125.1000 ;
	    RECT 10.7000 121.1000 11.1000 124.7000 ;
	    RECT 11.8000 121.1000 12.2000 125.8000 ;
	    RECT 15.5000 125.7000 15.9000 125.8000 ;
	    RECT 14.2000 125.4000 15.9000 125.7000 ;
	    RECT 14.2000 125.1000 14.5000 125.4000 ;
	    RECT 16.3000 125.2000 16.6000 125.8000 ;
	    RECT 19.0000 125.4000 19.4000 126.2000 ;
	    RECT 19.8000 126.1000 20.1000 126.8000 ;
	    RECT 22.2000 126.4000 22.6000 126.8000 ;
	    RECT 21.4000 126.1000 21.8000 126.2000 ;
	    RECT 23.0000 126.1000 23.3000 127.9000 ;
	    RECT 23.8000 127.8000 24.2000 128.2000 ;
	    RECT 23.8000 126.1000 24.2000 126.2000 ;
	    RECT 19.8000 125.8000 22.2000 126.1000 ;
	    RECT 23.0000 125.8000 24.2000 126.1000 ;
	    RECT 25.4000 126.1000 25.8000 129.9000 ;
	    RECT 27.0000 128.9000 27.4000 129.9000 ;
	    RECT 27.0000 128.1000 27.3000 128.9000 ;
	    RECT 26.2000 127.8000 27.3000 128.1000 ;
	    RECT 28.6000 128.0000 29.0000 129.9000 ;
	    RECT 30.2000 128.0000 30.6000 129.9000 ;
	    RECT 28.6000 127.9000 30.6000 128.0000 ;
	    RECT 31.0000 127.9000 31.4000 129.9000 ;
	    RECT 33.1000 129.2000 33.9000 129.9000 ;
	    RECT 32.6000 128.8000 33.9000 129.2000 ;
	    RECT 33.1000 127.9000 33.9000 128.8000 ;
	    RECT 26.2000 127.2000 26.5000 127.8000 ;
	    RECT 27.0000 127.2000 27.3000 127.8000 ;
	    RECT 28.7000 127.7000 30.5000 127.9000 ;
	    RECT 29.0000 127.2000 29.4000 127.4000 ;
	    RECT 31.0000 127.2000 31.3000 127.9000 ;
	    RECT 26.2000 126.8000 26.6000 127.2000 ;
	    RECT 27.0000 126.8000 27.4000 127.2000 ;
	    RECT 28.6000 126.9000 29.4000 127.2000 ;
	    RECT 28.6000 126.8000 29.0000 126.9000 ;
	    RECT 30.1000 126.8000 31.4000 127.2000 ;
	    RECT 32.6000 126.8000 33.0000 127.2000 ;
	    RECT 26.2000 126.1000 26.6000 126.2000 ;
	    RECT 25.4000 125.8000 26.6000 126.1000 ;
	    RECT 16.3000 125.1000 17.0000 125.2000 ;
	    RECT 19.8000 125.1000 20.1000 125.8000 ;
	    RECT 21.8000 125.6000 22.2000 125.8000 ;
	    RECT 23.8000 125.1000 24.1000 125.8000 ;
	    RECT 13.4000 124.8000 14.5000 125.1000 ;
	    RECT 13.4000 121.1000 13.8000 124.8000 ;
	    RECT 14.1000 124.7000 14.5000 124.8000 ;
	    RECT 15.6000 124.8000 17.0000 125.1000 ;
	    RECT 17.4000 124.8000 18.6000 125.1000 ;
	    RECT 15.6000 121.1000 16.4000 124.8000 ;
	    RECT 17.4000 124.7000 17.8000 124.8000 ;
	    RECT 18.2000 121.1000 18.6000 124.8000 ;
	    RECT 19.3000 124.7000 20.2000 125.1000 ;
	    RECT 21.4000 124.8000 23.4000 125.1000 ;
	    RECT 19.3000 121.1000 19.7000 124.7000 ;
	    RECT 21.4000 121.1000 21.8000 124.8000 ;
	    RECT 23.0000 121.1000 23.4000 124.8000 ;
	    RECT 23.8000 121.1000 24.2000 125.1000 ;
	    RECT 25.4000 121.1000 25.8000 125.8000 ;
	    RECT 26.2000 125.4000 26.6000 125.8000 ;
	    RECT 27.0000 125.1000 27.3000 126.8000 ;
	    RECT 27.8000 126.1000 28.2000 126.2000 ;
	    RECT 29.4000 126.1000 29.8000 126.6000 ;
	    RECT 27.8000 125.8000 29.8000 126.1000 ;
	    RECT 30.1000 126.2000 30.4000 126.8000 ;
	    RECT 32.7000 126.6000 33.0000 126.8000 ;
	    RECT 32.7000 126.2000 33.1000 126.6000 ;
	    RECT 33.4000 126.2000 33.7000 127.9000 ;
	    RECT 35.8000 127.8000 36.2000 128.6000 ;
	    RECT 34.2000 126.4000 34.6000 127.2000 ;
	    RECT 30.1000 125.8000 30.6000 126.2000 ;
	    RECT 30.1000 125.1000 30.4000 125.8000 ;
	    RECT 31.8000 125.4000 32.2000 126.2000 ;
	    RECT 33.4000 125.8000 33.8000 126.2000 ;
	    RECT 35.0000 126.1000 35.4000 126.2000 ;
	    RECT 34.6000 125.8000 35.4000 126.1000 ;
	    RECT 33.4000 125.7000 33.7000 125.8000 ;
	    RECT 32.7000 125.4000 33.7000 125.7000 ;
	    RECT 34.6000 125.6000 35.0000 125.8000 ;
	    RECT 31.0000 125.1000 31.4000 125.2000 ;
	    RECT 32.7000 125.1000 33.0000 125.4000 ;
	    RECT 36.6000 125.1000 37.0000 129.9000 ;
	    RECT 37.7000 128.2000 38.1000 129.9000 ;
	    RECT 37.7000 127.9000 38.6000 128.2000 ;
	    RECT 39.8000 127.9000 40.2000 129.9000 ;
	    RECT 40.6000 128.0000 41.0000 129.9000 ;
	    RECT 42.2000 128.0000 42.6000 129.9000 ;
	    RECT 40.6000 127.9000 42.6000 128.0000 ;
	    RECT 37.4000 125.1000 37.8000 125.2000 ;
	    RECT 26.5000 124.7000 27.4000 125.1000 ;
	    RECT 29.9000 124.8000 30.4000 125.1000 ;
	    RECT 30.7000 124.8000 31.4000 125.1000 ;
	    RECT 26.5000 121.1000 26.9000 124.7000 ;
	    RECT 29.9000 121.1000 30.3000 124.8000 ;
	    RECT 30.7000 124.2000 31.0000 124.8000 ;
	    RECT 30.6000 123.8000 31.0000 124.2000 ;
	    RECT 31.8000 121.4000 32.2000 125.1000 ;
	    RECT 32.6000 121.7000 33.0000 125.1000 ;
	    RECT 33.4000 124.8000 35.4000 125.1000 ;
	    RECT 33.4000 121.4000 33.8000 124.8000 ;
	    RECT 31.8000 121.1000 33.8000 121.4000 ;
	    RECT 35.0000 121.1000 35.4000 124.8000 ;
	    RECT 36.6000 124.8000 37.8000 125.1000 ;
	    RECT 36.6000 121.1000 37.0000 124.8000 ;
	    RECT 37.4000 124.4000 37.8000 124.8000 ;
	    RECT 38.2000 121.1000 38.6000 127.9000 ;
	    RECT 39.0000 126.8000 39.4000 127.6000 ;
	    RECT 39.9000 127.2000 40.2000 127.9000 ;
	    RECT 40.7000 127.7000 42.5000 127.9000 ;
	    RECT 41.8000 127.2000 42.2000 127.4000 ;
	    RECT 39.8000 126.8000 41.1000 127.2000 ;
	    RECT 41.8000 126.9000 42.6000 127.2000 ;
	    RECT 42.2000 126.8000 42.6000 126.9000 ;
	    RECT 40.8000 125.2000 41.1000 126.8000 ;
	    RECT 41.4000 126.1000 41.8000 126.6000 ;
	    RECT 43.0000 126.1000 43.4000 129.9000 ;
	    RECT 43.8000 127.8000 44.2000 128.6000 ;
	    RECT 43.8000 127.2000 44.1000 127.8000 ;
	    RECT 44.6000 127.5000 45.0000 129.9000 ;
	    RECT 46.8000 129.2000 47.2000 129.9000 ;
	    RECT 46.2000 128.9000 47.2000 129.2000 ;
	    RECT 49.0000 128.9000 49.4000 129.9000 ;
	    RECT 51.1000 129.2000 51.7000 129.9000 ;
	    RECT 51.0000 128.9000 51.7000 129.2000 ;
	    RECT 46.2000 128.5000 46.6000 128.9000 ;
	    RECT 49.0000 128.6000 49.3000 128.9000 ;
	    RECT 47.0000 128.2000 47.4000 128.6000 ;
	    RECT 47.9000 128.3000 49.3000 128.6000 ;
	    RECT 51.0000 128.5000 51.4000 128.9000 ;
	    RECT 47.9000 128.2000 48.3000 128.3000 ;
	    RECT 43.8000 126.8000 44.2000 127.2000 ;
	    RECT 45.0000 127.1000 45.8000 127.2000 ;
	    RECT 47.1000 127.1000 47.4000 128.2000 ;
	    RECT 51.9000 127.7000 52.3000 127.8000 ;
	    RECT 53.4000 127.7000 53.8000 129.9000 ;
	    RECT 54.2000 127.9000 54.6000 129.9000 ;
	    RECT 56.3000 129.1000 56.7000 129.9000 ;
	    RECT 57.4000 129.1000 57.8000 129.2000 ;
	    RECT 56.3000 128.8000 57.8000 129.1000 ;
	    RECT 56.3000 128.4000 56.7000 128.8000 ;
	    RECT 56.3000 127.9000 57.0000 128.4000 ;
	    RECT 51.9000 127.4000 53.8000 127.7000 ;
	    RECT 54.3000 127.8000 54.6000 127.9000 ;
	    RECT 54.3000 127.6000 55.2000 127.8000 ;
	    RECT 54.3000 127.5000 56.4000 127.6000 ;
	    RECT 49.9000 127.1000 50.3000 127.2000 ;
	    RECT 45.0000 126.8000 50.5000 127.1000 ;
	    RECT 46.5000 126.7000 46.9000 126.8000 ;
	    RECT 41.4000 125.8000 43.4000 126.1000 ;
	    RECT 45.7000 126.2000 46.1000 126.3000 ;
	    RECT 47.0000 126.2000 47.4000 126.3000 ;
	    RECT 50.2000 126.2000 50.5000 126.8000 ;
	    RECT 51.0000 126.4000 51.4000 126.5000 ;
	    RECT 45.7000 125.9000 48.2000 126.2000 ;
	    RECT 47.8000 125.8000 48.2000 125.9000 ;
	    RECT 50.2000 125.8000 50.6000 126.2000 ;
	    RECT 51.0000 126.1000 52.9000 126.4000 ;
	    RECT 52.5000 126.0000 52.9000 126.1000 ;
	    RECT 39.8000 125.1000 40.2000 125.2000 ;
	    RECT 39.8000 124.8000 40.5000 125.1000 ;
	    RECT 40.8000 124.8000 41.8000 125.2000 ;
	    RECT 40.2000 124.2000 40.5000 124.8000 ;
	    RECT 40.2000 123.8000 40.6000 124.2000 ;
	    RECT 40.9000 121.1000 41.3000 124.8000 ;
	    RECT 43.0000 121.1000 43.4000 125.8000 ;
	    RECT 44.6000 125.5000 47.4000 125.6000 ;
	    RECT 44.6000 125.4000 47.5000 125.5000 ;
	    RECT 44.6000 125.3000 49.5000 125.4000 ;
	    RECT 44.6000 121.1000 45.0000 125.3000 ;
	    RECT 47.1000 125.1000 49.5000 125.3000 ;
	    RECT 46.2000 124.5000 48.9000 124.8000 ;
	    RECT 46.2000 124.4000 46.6000 124.5000 ;
	    RECT 48.5000 124.4000 48.9000 124.5000 ;
	    RECT 49.2000 124.5000 49.5000 125.1000 ;
	    RECT 50.2000 125.2000 50.5000 125.8000 ;
	    RECT 51.7000 125.7000 52.1000 125.8000 ;
	    RECT 53.4000 125.7000 53.8000 127.4000 ;
	    RECT 54.9000 127.3000 56.4000 127.5000 ;
	    RECT 56.0000 127.2000 56.4000 127.3000 ;
	    RECT 54.2000 126.4000 54.6000 127.2000 ;
	    RECT 55.2000 126.9000 55.6000 127.0000 ;
	    RECT 55.1000 126.6000 55.6000 126.9000 ;
	    RECT 55.1000 126.2000 55.4000 126.6000 ;
	    RECT 55.0000 125.8000 55.4000 126.2000 ;
	    RECT 51.7000 125.4000 53.8000 125.7000 ;
	    RECT 56.0000 125.5000 56.3000 127.2000 ;
	    RECT 56.7000 126.2000 57.0000 127.9000 ;
	    RECT 59.0000 127.9000 59.4000 129.9000 ;
	    RECT 60.6000 128.9000 61.0000 129.9000 ;
	    RECT 63.0000 128.9000 63.4000 129.9000 ;
	    RECT 59.0000 126.2000 59.3000 127.9000 ;
	    RECT 60.6000 127.8000 60.9000 128.9000 ;
	    RECT 61.4000 128.1000 61.8000 128.6000 ;
	    RECT 62.2000 128.1000 62.6000 128.6000 ;
	    RECT 61.4000 127.8000 62.6000 128.1000 ;
	    RECT 63.1000 127.8000 63.4000 128.9000 ;
	    RECT 64.6000 127.9000 65.0000 129.9000 ;
	    RECT 65.4000 127.9000 65.8000 129.9000 ;
	    RECT 67.5000 129.2000 67.9000 129.9000 ;
	    RECT 67.5000 128.8000 68.2000 129.2000 ;
	    RECT 67.5000 128.4000 67.9000 128.8000 ;
	    RECT 67.5000 127.9000 68.2000 128.4000 ;
	    RECT 59.7000 127.5000 60.9000 127.8000 ;
	    RECT 63.1000 127.5000 64.3000 127.8000 ;
	    RECT 56.6000 125.8000 57.0000 126.2000 ;
	    RECT 58.2000 126.1000 58.6000 126.2000 ;
	    RECT 59.0000 126.1000 59.4000 126.2000 ;
	    RECT 58.2000 125.8000 59.4000 126.1000 ;
	    RECT 59.7000 126.0000 60.0000 127.5000 ;
	    RECT 60.5000 127.1000 61.0000 127.2000 ;
	    RECT 61.4000 127.1000 61.8000 127.2000 ;
	    RECT 60.5000 126.8000 61.8000 127.1000 ;
	    RECT 63.0000 126.8000 63.5000 127.2000 ;
	    RECT 60.4000 126.4000 60.8000 126.8000 ;
	    RECT 63.2000 126.4000 63.6000 126.8000 ;
	    RECT 64.0000 126.0000 64.3000 127.5000 ;
	    RECT 64.7000 126.2000 65.0000 127.9000 ;
	    RECT 65.5000 127.8000 65.8000 127.9000 ;
	    RECT 65.5000 127.6000 66.4000 127.8000 ;
	    RECT 65.5000 127.5000 67.6000 127.6000 ;
	    RECT 66.1000 127.3000 67.6000 127.5000 ;
	    RECT 67.2000 127.2000 67.6000 127.3000 ;
	    RECT 65.4000 126.4000 65.8000 127.2000 ;
	    RECT 66.4000 126.9000 66.8000 127.0000 ;
	    RECT 66.3000 126.6000 66.8000 126.9000 ;
	    RECT 66.3000 126.2000 66.6000 126.6000 ;
	    RECT 50.2000 124.9000 51.4000 125.2000 ;
	    RECT 49.9000 124.5000 50.3000 124.6000 ;
	    RECT 49.2000 124.2000 50.3000 124.5000 ;
	    RECT 51.1000 124.4000 51.4000 124.9000 ;
	    RECT 51.1000 124.0000 51.8000 124.4000 ;
	    RECT 47.9000 123.7000 48.3000 123.8000 ;
	    RECT 49.3000 123.7000 49.7000 123.8000 ;
	    RECT 46.2000 123.1000 46.6000 123.5000 ;
	    RECT 47.9000 123.4000 49.7000 123.7000 ;
	    RECT 49.0000 123.1000 49.3000 123.4000 ;
	    RECT 51.0000 123.1000 51.4000 123.5000 ;
	    RECT 46.2000 122.8000 47.2000 123.1000 ;
	    RECT 46.8000 121.1000 47.2000 122.8000 ;
	    RECT 49.0000 121.1000 49.4000 123.1000 ;
	    RECT 51.1000 121.1000 51.7000 123.1000 ;
	    RECT 53.4000 121.1000 53.8000 125.4000 ;
	    RECT 55.1000 125.2000 56.3000 125.5000 ;
	    RECT 55.1000 123.1000 55.4000 125.2000 ;
	    RECT 56.7000 125.1000 57.0000 125.8000 ;
	    RECT 55.0000 121.1000 55.4000 123.1000 ;
	    RECT 56.6000 121.1000 57.0000 125.1000 ;
	    RECT 59.0000 125.1000 59.3000 125.8000 ;
	    RECT 59.7000 125.7000 60.1000 126.0000 ;
	    RECT 63.9000 125.7000 64.3000 126.0000 ;
	    RECT 64.6000 125.8000 65.0000 126.2000 ;
	    RECT 66.2000 125.8000 66.6000 126.2000 ;
	    RECT 59.7000 125.6000 61.8000 125.7000 ;
	    RECT 59.8000 125.4000 61.8000 125.6000 ;
	    RECT 59.0000 124.8000 59.7000 125.1000 ;
	    RECT 59.3000 121.1000 59.7000 124.8000 ;
	    RECT 61.4000 121.1000 61.8000 125.4000 ;
	    RECT 62.2000 125.6000 64.3000 125.7000 ;
	    RECT 62.2000 125.4000 64.2000 125.6000 ;
	    RECT 62.2000 121.1000 62.6000 125.4000 ;
	    RECT 64.7000 125.1000 65.0000 125.8000 ;
	    RECT 67.2000 125.5000 67.5000 127.2000 ;
	    RECT 67.9000 126.2000 68.2000 127.9000 ;
	    RECT 67.8000 125.8000 68.2000 126.2000 ;
	    RECT 64.3000 124.8000 65.0000 125.1000 ;
	    RECT 66.3000 125.2000 67.5000 125.5000 ;
	    RECT 64.3000 121.1000 64.7000 124.8000 ;
	    RECT 66.3000 123.1000 66.6000 125.2000 ;
	    RECT 67.9000 125.1000 68.2000 125.8000 ;
	    RECT 66.2000 121.1000 66.6000 123.1000 ;
	    RECT 67.8000 121.1000 68.2000 125.1000 ;
	    RECT 68.6000 127.7000 69.0000 129.9000 ;
	    RECT 70.7000 129.2000 71.3000 129.9000 ;
	    RECT 70.7000 128.9000 71.4000 129.2000 ;
	    RECT 73.0000 128.9000 73.4000 129.9000 ;
	    RECT 75.2000 129.2000 75.6000 129.9000 ;
	    RECT 75.2000 128.9000 76.2000 129.2000 ;
	    RECT 71.0000 128.5000 71.4000 128.9000 ;
	    RECT 73.1000 128.6000 73.4000 128.9000 ;
	    RECT 73.1000 128.3000 74.5000 128.6000 ;
	    RECT 74.1000 128.2000 74.5000 128.3000 ;
	    RECT 75.0000 128.2000 75.4000 128.6000 ;
	    RECT 75.8000 128.5000 76.2000 128.9000 ;
	    RECT 70.1000 127.7000 70.5000 127.8000 ;
	    RECT 68.6000 127.4000 70.5000 127.7000 ;
	    RECT 68.6000 125.7000 69.0000 127.4000 ;
	    RECT 72.1000 127.1000 72.5000 127.2000 ;
	    RECT 75.0000 127.1000 75.3000 128.2000 ;
	    RECT 77.4000 127.5000 77.8000 129.9000 ;
	    RECT 78.3000 128.2000 78.7000 128.6000 ;
	    RECT 78.2000 127.8000 78.6000 128.2000 ;
	    RECT 79.0000 127.9000 79.4000 129.9000 ;
	    RECT 81.4000 127.9000 81.8000 129.9000 ;
	    RECT 82.2000 128.0000 82.6000 129.9000 ;
	    RECT 83.8000 128.0000 84.2000 129.9000 ;
	    RECT 82.2000 127.9000 84.2000 128.0000 ;
	    RECT 79.1000 127.2000 79.4000 127.9000 ;
	    RECT 81.5000 127.2000 81.8000 127.9000 ;
	    RECT 82.3000 127.7000 84.1000 127.9000 ;
	    RECT 85.4000 127.6000 85.8000 129.9000 ;
	    RECT 87.0000 127.6000 87.4000 129.9000 ;
	    RECT 88.6000 127.6000 89.0000 129.9000 ;
	    RECT 90.2000 127.6000 90.6000 129.9000 ;
	    RECT 92.6000 128.8000 93.0000 129.9000 ;
	    RECT 91.8000 127.8000 92.2000 128.6000 ;
	    RECT 83.4000 127.2000 83.8000 127.4000 ;
	    RECT 85.4000 127.2000 86.3000 127.6000 ;
	    RECT 87.0000 127.2000 88.1000 127.6000 ;
	    RECT 88.6000 127.2000 89.7000 127.6000 ;
	    RECT 90.2000 127.2000 91.4000 127.6000 ;
	    RECT 92.7000 127.2000 93.0000 128.8000 ;
	    RECT 95.0000 128.2000 95.4000 129.9000 ;
	    RECT 76.6000 127.1000 77.4000 127.2000 ;
	    RECT 71.9000 126.8000 77.4000 127.1000 ;
	    RECT 79.0000 126.8000 79.4000 127.2000 ;
	    RECT 71.0000 126.4000 71.4000 126.5000 ;
	    RECT 69.5000 126.1000 71.4000 126.4000 ;
	    RECT 69.5000 126.0000 69.9000 126.1000 ;
	    RECT 70.3000 125.7000 70.7000 125.8000 ;
	    RECT 68.6000 125.4000 70.7000 125.7000 ;
	    RECT 68.6000 121.1000 69.0000 125.4000 ;
	    RECT 71.9000 125.2000 72.2000 126.8000 ;
	    RECT 75.5000 126.7000 75.9000 126.8000 ;
	    RECT 75.0000 126.2000 75.4000 126.3000 ;
	    RECT 76.3000 126.2000 76.7000 126.3000 ;
	    RECT 74.2000 125.9000 76.7000 126.2000 ;
	    RECT 78.2000 126.1000 78.6000 126.2000 ;
	    RECT 79.1000 126.1000 79.4000 126.8000 ;
	    RECT 79.8000 127.1000 80.2000 127.2000 ;
	    RECT 81.4000 127.1000 82.7000 127.2000 ;
	    RECT 79.8000 126.8000 82.7000 127.1000 ;
	    RECT 83.4000 126.9000 84.2000 127.2000 ;
	    RECT 83.8000 126.8000 84.2000 126.9000 ;
	    RECT 85.9000 126.9000 86.3000 127.2000 ;
	    RECT 87.7000 126.9000 88.1000 127.2000 ;
	    RECT 89.3000 126.9000 89.7000 127.2000 ;
	    RECT 79.8000 126.4000 80.2000 126.8000 ;
	    RECT 80.6000 126.1000 81.0000 126.2000 ;
	    RECT 74.2000 125.8000 74.6000 125.9000 ;
	    RECT 78.2000 125.8000 79.4000 126.1000 ;
	    RECT 80.2000 125.8000 81.0000 126.1000 ;
	    RECT 75.0000 125.5000 77.8000 125.6000 ;
	    RECT 74.9000 125.4000 77.8000 125.5000 ;
	    RECT 71.0000 124.9000 72.2000 125.2000 ;
	    RECT 72.9000 125.3000 77.8000 125.4000 ;
	    RECT 72.9000 125.1000 75.3000 125.3000 ;
	    RECT 71.0000 124.4000 71.3000 124.9000 ;
	    RECT 70.6000 124.2000 71.3000 124.4000 ;
	    RECT 72.1000 124.5000 72.5000 124.6000 ;
	    RECT 72.9000 124.5000 73.2000 125.1000 ;
	    RECT 72.1000 124.2000 73.2000 124.5000 ;
	    RECT 73.5000 124.5000 76.2000 124.8000 ;
	    RECT 73.5000 124.4000 73.9000 124.5000 ;
	    RECT 75.8000 124.4000 76.2000 124.5000 ;
	    RECT 70.2000 124.0000 71.3000 124.2000 ;
	    RECT 70.2000 123.8000 70.9000 124.0000 ;
	    RECT 72.7000 123.7000 73.1000 123.8000 ;
	    RECT 74.1000 123.7000 74.5000 123.8000 ;
	    RECT 71.0000 123.1000 71.4000 123.5000 ;
	    RECT 72.7000 123.4000 74.5000 123.7000 ;
	    RECT 73.1000 123.1000 73.4000 123.4000 ;
	    RECT 75.8000 123.1000 76.2000 123.5000 ;
	    RECT 70.7000 121.1000 71.3000 123.1000 ;
	    RECT 73.0000 121.1000 73.4000 123.1000 ;
	    RECT 75.2000 122.8000 76.2000 123.1000 ;
	    RECT 75.2000 121.1000 75.6000 122.8000 ;
	    RECT 77.4000 121.1000 77.8000 125.3000 ;
	    RECT 78.3000 125.1000 78.6000 125.8000 ;
	    RECT 80.2000 125.6000 80.6000 125.8000 ;
	    RECT 81.4000 125.1000 81.8000 125.2000 ;
	    RECT 82.4000 125.1000 82.7000 126.8000 ;
	    RECT 83.0000 126.1000 83.4000 126.6000 ;
	    RECT 85.9000 126.5000 87.2000 126.9000 ;
	    RECT 87.7000 126.5000 88.9000 126.9000 ;
	    RECT 89.3000 126.5000 90.6000 126.9000 ;
	    RECT 84.6000 126.1000 85.0000 126.2000 ;
	    RECT 83.0000 125.8000 85.0000 126.1000 ;
	    RECT 85.9000 125.8000 86.3000 126.5000 ;
	    RECT 87.7000 125.8000 88.1000 126.5000 ;
	    RECT 89.3000 125.8000 89.7000 126.5000 ;
	    RECT 91.0000 125.8000 91.4000 127.2000 ;
	    RECT 92.6000 126.8000 93.0000 127.2000 ;
	    RECT 85.4000 125.4000 86.3000 125.8000 ;
	    RECT 87.0000 125.4000 88.1000 125.8000 ;
	    RECT 88.6000 125.4000 89.7000 125.8000 ;
	    RECT 90.2000 125.4000 91.4000 125.8000 ;
	    RECT 78.2000 121.1000 78.6000 125.1000 ;
	    RECT 79.0000 124.8000 81.0000 125.1000 ;
	    RECT 81.4000 124.8000 82.1000 125.1000 ;
	    RECT 82.4000 124.8000 82.9000 125.1000 ;
	    RECT 79.0000 121.1000 79.4000 124.8000 ;
	    RECT 80.6000 121.1000 81.0000 124.8000 ;
	    RECT 81.8000 124.2000 82.1000 124.8000 ;
	    RECT 81.4000 123.8000 82.2000 124.2000 ;
	    RECT 82.5000 121.1000 82.9000 124.8000 ;
	    RECT 85.4000 121.1000 85.8000 125.4000 ;
	    RECT 87.0000 121.1000 87.4000 125.4000 ;
	    RECT 88.6000 121.1000 89.0000 125.4000 ;
	    RECT 90.2000 121.1000 90.6000 125.4000 ;
	    RECT 92.7000 125.1000 93.0000 126.8000 ;
	    RECT 93.4000 127.8000 93.8000 128.2000 ;
	    RECT 94.9000 127.9000 95.4000 128.2000 ;
	    RECT 93.4000 127.1000 93.7000 127.8000 ;
	    RECT 94.9000 127.2000 95.2000 127.9000 ;
	    RECT 96.6000 127.6000 97.0000 129.9000 ;
	    RECT 97.4000 127.9000 97.8000 129.9000 ;
	    RECT 99.5000 128.4000 99.9000 129.9000 ;
	    RECT 99.5000 127.9000 100.2000 128.4000 ;
	    RECT 101.9000 128.2000 102.3000 129.9000 ;
	    RECT 95.7000 127.3000 97.0000 127.6000 ;
	    RECT 97.5000 127.8000 97.8000 127.9000 ;
	    RECT 97.5000 127.6000 98.4000 127.8000 ;
	    RECT 97.5000 127.5000 99.6000 127.6000 ;
	    RECT 98.1000 127.3000 99.6000 127.5000 ;
	    RECT 94.9000 127.1000 95.4000 127.2000 ;
	    RECT 93.4000 126.8000 95.4000 127.1000 ;
	    RECT 93.4000 126.2000 93.7000 126.8000 ;
	    RECT 93.4000 125.4000 93.8000 126.2000 ;
	    RECT 94.9000 125.1000 95.2000 126.8000 ;
	    RECT 95.7000 126.5000 96.0000 127.3000 ;
	    RECT 99.2000 127.2000 99.6000 127.3000 ;
	    RECT 95.5000 126.1000 96.0000 126.5000 ;
	    RECT 95.7000 125.1000 96.0000 126.1000 ;
	    RECT 96.5000 126.2000 96.9000 126.6000 ;
	    RECT 97.4000 126.4000 97.8000 127.2000 ;
	    RECT 98.2000 126.6000 98.8000 127.0000 ;
	    RECT 98.3000 126.2000 98.6000 126.6000 ;
	    RECT 96.5000 125.8000 97.0000 126.2000 ;
	    RECT 98.2000 125.8000 98.6000 126.2000 ;
	    RECT 99.2000 125.5000 99.5000 127.2000 ;
	    RECT 99.9000 126.2000 100.2000 127.9000 ;
	    RECT 101.4000 127.9000 102.3000 128.2000 ;
	    RECT 103.0000 128.0000 103.4000 129.9000 ;
	    RECT 104.6000 128.0000 105.0000 129.9000 ;
	    RECT 103.0000 127.9000 105.0000 128.0000 ;
	    RECT 105.4000 127.9000 105.8000 129.9000 ;
	    RECT 107.0000 128.9000 107.4000 129.9000 ;
	    RECT 100.6000 126.8000 101.0000 127.6000 ;
	    RECT 99.8000 125.8000 100.2000 126.2000 ;
	    RECT 98.3000 125.2000 99.5000 125.5000 ;
	    RECT 92.6000 124.7000 93.5000 125.1000 ;
	    RECT 93.1000 121.1000 93.5000 124.7000 ;
	    RECT 94.9000 124.6000 95.4000 125.1000 ;
	    RECT 95.7000 124.8000 97.0000 125.1000 ;
	    RECT 95.0000 121.1000 95.4000 124.6000 ;
	    RECT 96.6000 121.1000 97.0000 124.8000 ;
	    RECT 98.3000 123.1000 98.6000 125.2000 ;
	    RECT 99.9000 125.1000 100.2000 125.8000 ;
	    RECT 98.2000 121.1000 98.6000 123.1000 ;
	    RECT 99.8000 121.1000 100.2000 125.1000 ;
	    RECT 101.4000 121.1000 101.8000 127.9000 ;
	    RECT 103.1000 127.7000 104.9000 127.9000 ;
	    RECT 103.4000 127.2000 103.8000 127.4000 ;
	    RECT 105.4000 127.2000 105.7000 127.9000 ;
	    RECT 106.2000 127.8000 106.6000 128.6000 ;
	    RECT 107.1000 127.8000 107.4000 128.9000 ;
	    RECT 108.6000 129.1000 109.0000 129.9000 ;
	    RECT 111.3000 129.2000 111.7000 129.9000 ;
	    RECT 110.2000 129.1000 110.6000 129.2000 ;
	    RECT 108.6000 128.8000 110.6000 129.1000 ;
	    RECT 111.0000 128.8000 111.7000 129.2000 ;
	    RECT 108.6000 127.9000 109.0000 128.8000 ;
	    RECT 111.3000 128.2000 111.7000 128.8000 ;
	    RECT 111.3000 127.9000 112.2000 128.2000 ;
	    RECT 107.1000 127.5000 108.3000 127.8000 ;
	    RECT 102.2000 127.1000 102.6000 127.2000 ;
	    RECT 103.0000 127.1000 103.8000 127.2000 ;
	    RECT 102.2000 126.9000 103.8000 127.1000 ;
	    RECT 104.5000 127.1000 105.8000 127.2000 ;
	    RECT 107.0000 127.1000 107.5000 127.2000 ;
	    RECT 102.2000 126.8000 103.4000 126.9000 ;
	    RECT 104.5000 126.8000 107.5000 127.1000 ;
	    RECT 103.8000 125.8000 104.2000 126.6000 ;
	    RECT 102.2000 124.4000 102.6000 125.2000 ;
	    RECT 104.5000 125.1000 104.8000 126.8000 ;
	    RECT 107.2000 126.4000 107.6000 126.8000 ;
	    RECT 108.0000 126.0000 108.3000 127.5000 ;
	    RECT 108.7000 126.2000 109.0000 127.9000 ;
	    RECT 107.9000 125.7000 108.3000 126.0000 ;
	    RECT 108.6000 125.8000 109.0000 126.2000 ;
	    RECT 106.2000 125.6000 108.3000 125.7000 ;
	    RECT 106.2000 125.4000 108.2000 125.6000 ;
	    RECT 105.4000 125.1000 105.8000 125.2000 ;
	    RECT 104.3000 124.8000 104.8000 125.1000 ;
	    RECT 105.1000 124.8000 105.8000 125.1000 ;
	    RECT 104.3000 121.1000 104.7000 124.8000 ;
	    RECT 105.1000 124.2000 105.4000 124.8000 ;
	    RECT 105.0000 123.8000 105.4000 124.2000 ;
	    RECT 106.2000 121.1000 106.6000 125.4000 ;
	    RECT 108.7000 125.1000 109.0000 125.8000 ;
	    RECT 108.3000 124.8000 109.0000 125.1000 ;
	    RECT 108.3000 121.1000 108.7000 124.8000 ;
	    RECT 111.0000 124.4000 111.4000 125.2000 ;
	    RECT 111.8000 121.1000 112.2000 127.9000 ;
	    RECT 112.6000 126.8000 113.0000 127.6000 ;
	    RECT 115.2000 127.1000 115.6000 129.9000 ;
	    RECT 116.9000 128.4000 117.3000 129.9000 ;
	    RECT 116.6000 127.9000 117.3000 128.4000 ;
	    RECT 119.0000 127.9000 119.4000 129.9000 ;
	    RECT 115.2000 126.9000 116.1000 127.1000 ;
	    RECT 115.3000 126.8000 116.1000 126.9000 ;
	    RECT 114.2000 125.8000 115.0000 126.2000 ;
	    RECT 113.4000 124.8000 113.8000 125.6000 ;
	    RECT 115.8000 125.2000 116.1000 126.8000 ;
	    RECT 116.6000 126.2000 116.9000 127.9000 ;
	    RECT 119.0000 127.8000 119.3000 127.9000 ;
	    RECT 118.4000 127.6000 119.3000 127.8000 ;
	    RECT 117.2000 127.5000 119.3000 127.6000 ;
	    RECT 117.2000 127.3000 118.7000 127.5000 ;
	    RECT 117.2000 127.2000 117.6000 127.3000 ;
	    RECT 116.6000 125.8000 117.0000 126.2000 ;
	    RECT 115.8000 124.8000 116.2000 125.2000 ;
	    RECT 116.6000 125.1000 116.9000 125.8000 ;
	    RECT 117.3000 125.5000 117.6000 127.2000 ;
	    RECT 118.0000 126.9000 118.4000 127.0000 ;
	    RECT 118.0000 126.6000 118.5000 126.9000 ;
	    RECT 118.2000 126.2000 118.5000 126.6000 ;
	    RECT 119.0000 126.4000 119.4000 127.2000 ;
	    RECT 118.2000 125.8000 118.6000 126.2000 ;
	    RECT 119.8000 126.1000 120.2000 129.9000 ;
	    RECT 122.2000 128.9000 122.6000 129.9000 ;
	    RECT 122.2000 127.2000 122.5000 128.9000 ;
	    RECT 123.0000 127.8000 123.4000 128.6000 ;
	    RECT 123.8000 128.0000 124.2000 129.9000 ;
	    RECT 125.4000 128.0000 125.8000 129.9000 ;
	    RECT 123.8000 127.9000 125.8000 128.0000 ;
	    RECT 126.2000 128.1000 126.6000 129.9000 ;
	    RECT 127.8000 128.8000 128.2000 129.9000 ;
	    RECT 127.0000 128.1000 127.4000 128.6000 ;
	    RECT 123.9000 127.7000 125.7000 127.9000 ;
	    RECT 126.2000 127.8000 127.4000 128.1000 ;
	    RECT 126.2000 127.2000 126.5000 127.8000 ;
	    RECT 127.9000 127.2000 128.2000 128.8000 ;
	    RECT 129.4000 127.5000 129.8000 129.9000 ;
	    RECT 131.6000 129.2000 132.0000 129.9000 ;
	    RECT 131.0000 128.9000 132.0000 129.2000 ;
	    RECT 133.8000 128.9000 134.2000 129.9000 ;
	    RECT 135.9000 129.2000 136.5000 129.9000 ;
	    RECT 135.8000 128.9000 136.5000 129.2000 ;
	    RECT 131.0000 128.5000 131.4000 128.9000 ;
	    RECT 133.8000 128.6000 134.1000 128.9000 ;
	    RECT 131.8000 128.2000 132.2000 128.6000 ;
	    RECT 132.7000 128.3000 134.1000 128.6000 ;
	    RECT 135.8000 128.5000 136.2000 128.9000 ;
	    RECT 132.7000 128.2000 133.1000 128.3000 ;
	    RECT 122.2000 126.8000 122.6000 127.2000 ;
	    RECT 125.3000 126.8000 126.6000 127.2000 ;
	    RECT 127.8000 126.8000 128.2000 127.2000 ;
	    RECT 129.8000 127.1000 130.6000 127.2000 ;
	    RECT 131.9000 127.1000 132.2000 128.2000 ;
	    RECT 136.7000 127.7000 137.1000 127.8000 ;
	    RECT 138.2000 127.7000 138.6000 129.9000 ;
	    RECT 136.7000 127.4000 138.6000 127.7000 ;
	    RECT 134.7000 127.1000 135.4000 127.2000 ;
	    RECT 129.8000 126.8000 135.4000 127.1000 ;
	    RECT 121.4000 126.1000 121.8000 126.2000 ;
	    RECT 119.8000 125.8000 121.8000 126.1000 ;
	    RECT 117.3000 125.2000 118.5000 125.5000 ;
	    RECT 115.0000 123.8000 115.4000 124.6000 ;
	    RECT 115.8000 123.5000 116.1000 124.8000 ;
	    RECT 114.3000 123.2000 116.1000 123.5000 ;
	    RECT 114.2000 121.1000 114.6000 123.2000 ;
	    RECT 115.8000 123.1000 116.1000 123.2000 ;
	    RECT 115.8000 121.1000 116.2000 123.1000 ;
	    RECT 116.6000 121.1000 117.0000 125.1000 ;
	    RECT 118.2000 123.1000 118.5000 125.2000 ;
	    RECT 118.2000 121.1000 118.6000 123.1000 ;
	    RECT 119.8000 121.1000 120.2000 125.8000 ;
	    RECT 121.4000 125.4000 121.8000 125.8000 ;
	    RECT 122.2000 125.1000 122.5000 126.8000 ;
	    RECT 124.6000 125.8000 125.0000 126.6000 ;
	    RECT 125.3000 125.1000 125.6000 126.8000 ;
	    RECT 126.2000 125.1000 126.6000 125.2000 ;
	    RECT 127.9000 125.1000 128.2000 126.8000 ;
	    RECT 131.3000 126.7000 131.7000 126.8000 ;
	    RECT 130.5000 126.2000 130.9000 126.3000 ;
	    RECT 128.6000 125.4000 129.0000 126.2000 ;
	    RECT 130.5000 126.1000 133.0000 126.2000 ;
	    RECT 133.4000 126.1000 133.8000 126.2000 ;
	    RECT 130.5000 125.9000 133.8000 126.1000 ;
	    RECT 132.6000 125.8000 133.8000 125.9000 ;
	    RECT 129.4000 125.5000 132.2000 125.6000 ;
	    RECT 129.4000 125.4000 132.3000 125.5000 ;
	    RECT 129.4000 125.3000 134.3000 125.4000 ;
	    RECT 121.7000 124.7000 122.6000 125.1000 ;
	    RECT 125.1000 124.8000 125.6000 125.1000 ;
	    RECT 125.9000 124.8000 126.6000 125.1000 ;
	    RECT 121.7000 122.2000 122.1000 124.7000 ;
	    RECT 121.4000 121.8000 122.1000 122.2000 ;
	    RECT 121.7000 121.1000 122.1000 121.8000 ;
	    RECT 125.1000 121.1000 125.5000 124.8000 ;
	    RECT 125.9000 124.2000 126.2000 124.8000 ;
	    RECT 127.8000 124.7000 128.7000 125.1000 ;
	    RECT 125.8000 123.8000 126.2000 124.2000 ;
	    RECT 128.3000 121.1000 128.7000 124.7000 ;
	    RECT 129.4000 121.1000 129.8000 125.3000 ;
	    RECT 131.9000 125.1000 134.3000 125.3000 ;
	    RECT 131.0000 124.5000 133.7000 124.8000 ;
	    RECT 131.0000 124.4000 131.4000 124.5000 ;
	    RECT 133.3000 124.4000 133.7000 124.5000 ;
	    RECT 134.0000 124.5000 134.3000 125.1000 ;
	    RECT 135.0000 125.2000 135.3000 126.8000 ;
	    RECT 135.8000 126.4000 136.2000 126.5000 ;
	    RECT 135.8000 126.1000 137.7000 126.4000 ;
	    RECT 137.3000 126.0000 137.7000 126.1000 ;
	    RECT 136.5000 125.7000 136.9000 125.8000 ;
	    RECT 138.2000 125.7000 138.6000 127.4000 ;
	    RECT 140.6000 127.9000 141.0000 129.9000 ;
	    RECT 141.3000 128.2000 141.7000 128.6000 ;
	    RECT 141.4000 128.1000 141.8000 128.2000 ;
	    RECT 142.2000 128.1000 142.6000 129.9000 ;
	    RECT 139.8000 126.4000 140.2000 127.2000 ;
	    RECT 140.6000 127.1000 140.9000 127.9000 ;
	    RECT 141.4000 127.8000 142.6000 128.1000 ;
	    RECT 143.0000 128.0000 143.4000 129.9000 ;
	    RECT 144.6000 128.0000 145.0000 129.9000 ;
	    RECT 143.0000 127.9000 145.0000 128.0000 ;
	    RECT 146.2000 128.9000 146.6000 129.9000 ;
	    RECT 142.3000 127.2000 142.6000 127.8000 ;
	    RECT 143.1000 127.7000 144.9000 127.9000 ;
	    RECT 144.2000 127.2000 144.6000 127.4000 ;
	    RECT 146.2000 127.2000 146.5000 128.9000 ;
	    RECT 147.0000 127.8000 147.4000 128.6000 ;
	    RECT 149.4000 127.9000 149.8000 129.9000 ;
	    RECT 150.1000 128.2000 150.5000 128.6000 ;
	    RECT 152.3000 128.2000 152.7000 129.9000 ;
	    RECT 141.4000 127.1000 141.8000 127.2000 ;
	    RECT 140.6000 126.8000 141.8000 127.1000 ;
	    RECT 142.2000 126.8000 143.5000 127.2000 ;
	    RECT 144.2000 126.9000 145.0000 127.2000 ;
	    RECT 144.6000 126.8000 145.0000 126.9000 ;
	    RECT 145.4000 126.8000 145.8000 127.2000 ;
	    RECT 146.2000 126.8000 146.6000 127.2000 ;
	    RECT 139.0000 126.1000 139.4000 126.2000 ;
	    RECT 140.6000 126.1000 140.9000 126.8000 ;
	    RECT 141.4000 126.1000 141.8000 126.2000 ;
	    RECT 139.0000 125.8000 139.8000 126.1000 ;
	    RECT 140.6000 125.8000 141.8000 126.1000 ;
	    RECT 136.5000 125.4000 138.6000 125.7000 ;
	    RECT 139.4000 125.6000 139.8000 125.8000 ;
	    RECT 135.0000 124.9000 136.2000 125.2000 ;
	    RECT 134.7000 124.5000 135.1000 124.6000 ;
	    RECT 134.0000 124.2000 135.1000 124.5000 ;
	    RECT 135.9000 124.4000 136.2000 124.9000 ;
	    RECT 135.9000 124.0000 136.6000 124.4000 ;
	    RECT 132.7000 123.7000 133.1000 123.8000 ;
	    RECT 134.1000 123.7000 134.5000 123.8000 ;
	    RECT 131.0000 123.1000 131.4000 123.5000 ;
	    RECT 132.7000 123.4000 134.5000 123.7000 ;
	    RECT 133.8000 123.1000 134.1000 123.4000 ;
	    RECT 135.8000 123.1000 136.2000 123.5000 ;
	    RECT 131.0000 122.8000 132.0000 123.1000 ;
	    RECT 131.6000 121.1000 132.0000 122.8000 ;
	    RECT 133.8000 121.1000 134.2000 123.1000 ;
	    RECT 135.9000 121.1000 136.5000 123.1000 ;
	    RECT 138.2000 121.1000 138.6000 125.4000 ;
	    RECT 141.4000 125.1000 141.7000 125.8000 ;
	    RECT 142.2000 125.1000 142.6000 125.2000 ;
	    RECT 143.2000 125.1000 143.5000 126.8000 ;
	    RECT 143.8000 126.1000 144.2000 126.6000 ;
	    RECT 145.4000 126.2000 145.7000 126.8000 ;
	    RECT 145.4000 126.1000 145.8000 126.2000 ;
	    RECT 143.8000 125.8000 145.8000 126.1000 ;
	    RECT 145.4000 125.4000 145.8000 125.8000 ;
	    RECT 146.2000 125.1000 146.5000 126.8000 ;
	    RECT 148.6000 126.4000 149.0000 127.2000 ;
	    RECT 147.8000 126.1000 148.2000 126.2000 ;
	    RECT 149.4000 126.1000 149.7000 127.9000 ;
	    RECT 150.2000 127.8000 150.6000 128.2000 ;
	    RECT 151.8000 127.8000 152.9000 128.2000 ;
	    RECT 150.2000 127.1000 150.5000 127.8000 ;
	    RECT 151.0000 127.1000 151.4000 127.6000 ;
	    RECT 150.2000 126.8000 151.4000 127.1000 ;
	    RECT 150.2000 126.1000 150.6000 126.2000 ;
	    RECT 147.8000 125.8000 148.6000 126.1000 ;
	    RECT 149.4000 125.8000 150.6000 126.1000 ;
	    RECT 151.0000 125.8000 151.4000 126.2000 ;
	    RECT 148.2000 125.6000 148.6000 125.8000 ;
	    RECT 150.2000 125.1000 150.5000 125.8000 ;
	    RECT 151.0000 125.1000 151.3000 125.8000 ;
	    RECT 139.0000 124.8000 141.0000 125.1000 ;
	    RECT 139.0000 121.1000 139.4000 124.8000 ;
	    RECT 140.6000 121.1000 141.0000 124.8000 ;
	    RECT 141.4000 121.1000 141.8000 125.1000 ;
	    RECT 142.2000 124.8000 142.9000 125.1000 ;
	    RECT 143.2000 124.8000 143.7000 125.1000 ;
	    RECT 142.6000 124.2000 142.9000 124.8000 ;
	    RECT 142.6000 123.8000 143.0000 124.2000 ;
	    RECT 143.3000 121.1000 143.7000 124.8000 ;
	    RECT 145.7000 124.7000 146.6000 125.1000 ;
	    RECT 147.8000 124.8000 149.8000 125.1000 ;
	    RECT 145.7000 121.1000 146.1000 124.7000 ;
	    RECT 147.8000 121.1000 148.2000 124.8000 ;
	    RECT 149.4000 121.1000 149.8000 124.8000 ;
	    RECT 150.2000 124.8000 151.3000 125.1000 ;
	    RECT 150.2000 121.1000 150.6000 124.8000 ;
	    RECT 151.8000 121.1000 152.2000 127.8000 ;
	    RECT 152.6000 127.2000 152.9000 127.8000 ;
	    RECT 152.6000 126.8000 153.0000 127.2000 ;
	    RECT 152.6000 124.4000 153.0000 125.2000 ;
	    RECT 153.4000 121.1000 153.8000 129.9000 ;
	    RECT 154.2000 127.8000 154.6000 128.6000 ;
	    RECT 155.0000 128.0000 155.4000 129.9000 ;
	    RECT 156.6000 128.0000 157.0000 129.9000 ;
	    RECT 155.0000 127.9000 157.0000 128.0000 ;
	    RECT 157.4000 128.1000 157.8000 129.9000 ;
	    RECT 159.0000 128.8000 159.4000 129.9000 ;
	    RECT 155.1000 127.7000 156.9000 127.9000 ;
	    RECT 157.4000 127.8000 158.5000 128.1000 ;
	    RECT 155.4000 127.2000 155.8000 127.4000 ;
	    RECT 157.4000 127.2000 157.7000 127.8000 ;
	    RECT 158.2000 127.2000 158.5000 127.8000 ;
	    RECT 159.0000 127.2000 159.3000 128.8000 ;
	    RECT 159.8000 127.8000 160.2000 128.6000 ;
	    RECT 162.2000 127.6000 162.6000 129.9000 ;
	    RECT 163.8000 128.2000 164.2000 129.9000 ;
	    RECT 163.8000 127.9000 164.3000 128.2000 ;
	    RECT 162.2000 127.3000 163.5000 127.6000 ;
	    RECT 155.0000 126.9000 155.8000 127.2000 ;
	    RECT 155.0000 126.8000 155.4000 126.9000 ;
	    RECT 156.5000 126.8000 157.8000 127.2000 ;
	    RECT 158.2000 126.8000 158.6000 127.2000 ;
	    RECT 159.0000 126.8000 159.4000 127.2000 ;
	    RECT 154.2000 126.1000 154.6000 126.2000 ;
	    RECT 155.8000 126.1000 156.2000 126.6000 ;
	    RECT 154.2000 125.8000 156.2000 126.1000 ;
	    RECT 156.5000 125.1000 156.8000 126.8000 ;
	    RECT 158.2000 125.4000 158.6000 126.2000 ;
	    RECT 157.4000 125.1000 157.8000 125.2000 ;
	    RECT 159.0000 125.1000 159.3000 126.8000 ;
	    RECT 163.2000 126.5000 163.5000 127.3000 ;
	    RECT 164.0000 127.2000 164.3000 127.9000 ;
	    RECT 165.4000 127.5000 165.8000 129.9000 ;
	    RECT 167.6000 129.2000 168.0000 129.9000 ;
	    RECT 167.0000 128.9000 168.0000 129.2000 ;
	    RECT 169.8000 128.9000 170.2000 129.9000 ;
	    RECT 171.9000 129.2000 172.5000 129.9000 ;
	    RECT 171.8000 128.9000 172.5000 129.2000 ;
	    RECT 167.0000 128.5000 167.4000 128.9000 ;
	    RECT 169.8000 128.6000 170.1000 128.9000 ;
	    RECT 167.8000 128.2000 168.2000 128.6000 ;
	    RECT 168.7000 128.3000 170.1000 128.6000 ;
	    RECT 171.8000 128.5000 172.2000 128.9000 ;
	    RECT 168.7000 128.2000 169.1000 128.3000 ;
	    RECT 167.9000 127.2000 168.2000 128.2000 ;
	    RECT 172.7000 127.7000 173.1000 127.8000 ;
	    RECT 174.2000 127.7000 174.6000 129.9000 ;
	    RECT 175.3000 129.2000 175.7000 129.9000 ;
	    RECT 175.3000 128.8000 176.2000 129.2000 ;
	    RECT 175.3000 128.2000 175.7000 128.8000 ;
	    RECT 178.2000 128.2000 178.6000 129.9000 ;
	    RECT 175.3000 127.9000 176.2000 128.2000 ;
	    RECT 172.7000 127.4000 174.6000 127.7000 ;
	    RECT 163.8000 126.8000 164.3000 127.2000 ;
	    RECT 165.8000 127.1000 166.6000 127.2000 ;
	    RECT 167.8000 127.1000 168.2000 127.2000 ;
	    RECT 170.7000 127.1000 171.1000 127.2000 ;
	    RECT 165.8000 126.8000 171.3000 127.1000 ;
	    RECT 163.2000 126.1000 163.7000 126.5000 ;
	    RECT 163.2000 125.1000 163.5000 126.1000 ;
	    RECT 164.0000 125.1000 164.3000 126.8000 ;
	    RECT 167.3000 126.7000 167.7000 126.8000 ;
	    RECT 166.5000 126.2000 166.9000 126.3000 ;
	    RECT 166.5000 125.9000 169.0000 126.2000 ;
	    RECT 168.6000 125.8000 169.0000 125.9000 ;
	    RECT 156.3000 124.8000 156.8000 125.1000 ;
	    RECT 157.1000 124.8000 157.8000 125.1000 ;
	    RECT 156.3000 121.1000 156.7000 124.8000 ;
	    RECT 157.1000 124.2000 157.4000 124.8000 ;
	    RECT 157.0000 123.8000 157.4000 124.2000 ;
	    RECT 158.5000 124.7000 159.4000 125.1000 ;
	    RECT 162.2000 124.8000 163.5000 125.1000 ;
	    RECT 158.5000 121.1000 158.9000 124.7000 ;
	    RECT 162.2000 121.1000 162.6000 124.8000 ;
	    RECT 163.8000 124.6000 164.3000 125.1000 ;
	    RECT 165.4000 125.5000 168.2000 125.6000 ;
	    RECT 165.4000 125.4000 168.3000 125.5000 ;
	    RECT 165.4000 125.3000 170.3000 125.4000 ;
	    RECT 163.8000 121.1000 164.2000 124.6000 ;
	    RECT 165.4000 121.1000 165.8000 125.3000 ;
	    RECT 167.9000 125.1000 170.3000 125.3000 ;
	    RECT 167.0000 124.5000 169.7000 124.8000 ;
	    RECT 167.0000 124.4000 167.4000 124.5000 ;
	    RECT 169.3000 124.4000 169.7000 124.5000 ;
	    RECT 170.0000 124.5000 170.3000 125.1000 ;
	    RECT 171.0000 125.2000 171.3000 126.8000 ;
	    RECT 171.8000 126.4000 172.2000 126.5000 ;
	    RECT 171.8000 126.1000 173.7000 126.4000 ;
	    RECT 173.3000 126.0000 173.7000 126.1000 ;
	    RECT 172.5000 125.7000 172.9000 125.8000 ;
	    RECT 174.2000 125.7000 174.6000 127.4000 ;
	    RECT 172.5000 125.4000 174.6000 125.7000 ;
	    RECT 171.0000 124.9000 172.2000 125.2000 ;
	    RECT 170.7000 124.5000 171.1000 124.6000 ;
	    RECT 170.0000 124.2000 171.1000 124.5000 ;
	    RECT 171.9000 124.4000 172.2000 124.9000 ;
	    RECT 171.9000 124.0000 172.6000 124.4000 ;
	    RECT 168.7000 123.7000 169.1000 123.8000 ;
	    RECT 170.1000 123.7000 170.5000 123.8000 ;
	    RECT 167.0000 123.1000 167.4000 123.5000 ;
	    RECT 168.7000 123.4000 170.5000 123.7000 ;
	    RECT 169.8000 123.1000 170.1000 123.4000 ;
	    RECT 171.8000 123.1000 172.2000 123.5000 ;
	    RECT 167.0000 122.8000 168.0000 123.1000 ;
	    RECT 167.6000 121.1000 168.0000 122.8000 ;
	    RECT 169.8000 121.1000 170.2000 123.1000 ;
	    RECT 171.9000 121.1000 172.5000 123.1000 ;
	    RECT 174.2000 121.1000 174.6000 125.4000 ;
	    RECT 175.0000 124.4000 175.4000 125.2000 ;
	    RECT 175.8000 121.1000 176.2000 127.9000 ;
	    RECT 178.1000 127.9000 178.6000 128.2000 ;
	    RECT 176.6000 126.8000 177.0000 127.6000 ;
	    RECT 178.1000 127.2000 178.4000 127.9000 ;
	    RECT 179.8000 127.6000 180.2000 129.9000 ;
	    RECT 180.9000 129.2000 181.3000 129.9000 ;
	    RECT 180.6000 128.8000 181.3000 129.2000 ;
	    RECT 180.9000 128.2000 181.3000 128.8000 ;
	    RECT 183.8000 128.2000 184.2000 129.9000 ;
	    RECT 180.9000 127.9000 181.8000 128.2000 ;
	    RECT 178.9000 127.3000 180.2000 127.6000 ;
	    RECT 178.1000 126.8000 178.6000 127.2000 ;
	    RECT 178.1000 125.1000 178.4000 126.8000 ;
	    RECT 178.9000 126.5000 179.2000 127.3000 ;
	    RECT 178.7000 126.1000 179.2000 126.5000 ;
	    RECT 178.9000 125.1000 179.2000 126.1000 ;
	    RECT 179.7000 126.2000 180.1000 126.6000 ;
	    RECT 179.7000 125.8000 180.2000 126.2000 ;
	    RECT 178.1000 124.6000 178.6000 125.1000 ;
	    RECT 178.9000 124.8000 180.2000 125.1000 ;
	    RECT 178.2000 121.1000 178.6000 124.6000 ;
	    RECT 179.8000 121.1000 180.2000 124.8000 ;
	    RECT 180.6000 124.4000 181.0000 125.2000 ;
	    RECT 181.4000 121.1000 181.8000 127.9000 ;
	    RECT 183.7000 127.9000 184.2000 128.2000 ;
	    RECT 182.2000 126.8000 182.6000 127.6000 ;
	    RECT 183.7000 127.2000 184.0000 127.9000 ;
	    RECT 185.4000 127.6000 185.8000 129.9000 ;
	    RECT 186.5000 129.2000 186.9000 129.9000 ;
	    RECT 186.2000 128.8000 186.9000 129.2000 ;
	    RECT 186.5000 128.2000 186.9000 128.8000 ;
	    RECT 186.5000 127.9000 187.4000 128.2000 ;
	    RECT 184.5000 127.3000 185.8000 127.6000 ;
	    RECT 183.7000 126.8000 184.2000 127.2000 ;
	    RECT 183.7000 125.1000 184.0000 126.8000 ;
	    RECT 184.5000 126.5000 184.8000 127.3000 ;
	    RECT 184.3000 126.1000 184.8000 126.5000 ;
	    RECT 184.5000 125.1000 184.8000 126.1000 ;
	    RECT 185.3000 126.2000 185.7000 126.6000 ;
	    RECT 185.3000 125.8000 185.8000 126.2000 ;
	    RECT 183.7000 124.6000 184.2000 125.1000 ;
	    RECT 184.5000 124.8000 185.8000 125.1000 ;
	    RECT 183.8000 121.1000 184.2000 124.6000 ;
	    RECT 185.4000 121.1000 185.8000 124.8000 ;
	    RECT 186.2000 124.4000 186.6000 125.2000 ;
	    RECT 187.0000 121.1000 187.4000 127.9000 ;
	    RECT 187.8000 126.8000 188.2000 127.6000 ;
	    RECT 188.6000 126.8000 189.0000 127.6000 ;
	    RECT 187.8000 126.1000 188.1000 126.8000 ;
	    RECT 189.4000 126.1000 189.8000 129.9000 ;
	    RECT 190.5000 129.2000 190.9000 129.9000 ;
	    RECT 190.5000 128.8000 191.4000 129.2000 ;
	    RECT 190.5000 128.2000 190.9000 128.8000 ;
	    RECT 190.5000 127.9000 191.4000 128.2000 ;
	    RECT 187.8000 125.8000 189.8000 126.1000 ;
	    RECT 189.4000 125.1000 189.8000 125.8000 ;
	    RECT 190.2000 125.1000 190.6000 125.2000 ;
	    RECT 189.4000 124.8000 190.6000 125.1000 ;
	    RECT 189.4000 121.1000 189.8000 124.8000 ;
	    RECT 190.2000 123.8000 190.6000 124.8000 ;
	    RECT 191.0000 121.1000 191.4000 127.9000 ;
	    RECT 191.8000 126.8000 192.2000 127.6000 ;
	    RECT 193.2000 127.1000 193.6000 129.9000 ;
	    RECT 192.7000 126.9000 193.6000 127.1000 ;
	    RECT 195.8000 127.7000 196.2000 129.9000 ;
	    RECT 197.9000 129.2000 198.5000 129.9000 ;
	    RECT 197.9000 128.9000 198.6000 129.2000 ;
	    RECT 200.2000 128.9000 200.6000 129.9000 ;
	    RECT 202.4000 129.2000 202.8000 129.9000 ;
	    RECT 202.4000 128.9000 203.4000 129.2000 ;
	    RECT 198.2000 128.5000 198.6000 128.9000 ;
	    RECT 200.3000 128.6000 200.6000 128.9000 ;
	    RECT 200.3000 128.3000 201.7000 128.6000 ;
	    RECT 201.3000 128.2000 201.7000 128.3000 ;
	    RECT 202.2000 128.2000 202.6000 128.6000 ;
	    RECT 203.0000 128.5000 203.4000 128.9000 ;
	    RECT 197.3000 127.7000 197.7000 127.8000 ;
	    RECT 195.8000 127.4000 197.7000 127.7000 ;
	    RECT 192.7000 126.8000 193.5000 126.9000 ;
	    RECT 192.7000 125.2000 193.0000 126.8000 ;
	    RECT 193.8000 125.8000 194.6000 126.2000 ;
	    RECT 195.8000 125.7000 196.2000 127.4000 ;
	    RECT 199.3000 127.1000 199.7000 127.2000 ;
	    RECT 202.2000 127.1000 202.5000 128.2000 ;
	    RECT 204.6000 127.5000 205.0000 129.9000 ;
	    RECT 206.2000 128.8000 206.6000 129.9000 ;
	    RECT 205.4000 127.8000 205.8000 128.6000 ;
	    RECT 206.3000 127.2000 206.6000 128.8000 ;
	    RECT 203.8000 127.1000 204.6000 127.2000 ;
	    RECT 199.1000 126.8000 204.6000 127.1000 ;
	    RECT 206.2000 126.8000 206.6000 127.2000 ;
	    RECT 207.8000 126.8000 208.2000 127.6000 ;
	    RECT 198.2000 126.4000 198.6000 126.5000 ;
	    RECT 196.7000 126.1000 198.6000 126.4000 ;
	    RECT 199.1000 126.2000 199.4000 126.8000 ;
	    RECT 202.7000 126.7000 203.1000 126.8000 ;
	    RECT 202.2000 126.2000 202.6000 126.3000 ;
	    RECT 203.5000 126.2000 203.9000 126.3000 ;
	    RECT 196.7000 126.0000 197.1000 126.1000 ;
	    RECT 199.0000 125.8000 199.4000 126.2000 ;
	    RECT 201.4000 125.9000 203.9000 126.2000 ;
	    RECT 201.4000 125.8000 201.8000 125.9000 ;
	    RECT 197.5000 125.7000 197.9000 125.8000 ;
	    RECT 192.6000 124.8000 193.0000 125.2000 ;
	    RECT 195.0000 124.8000 195.4000 125.6000 ;
	    RECT 195.8000 125.4000 197.9000 125.7000 ;
	    RECT 192.7000 123.5000 193.0000 124.8000 ;
	    RECT 193.4000 123.8000 193.8000 124.6000 ;
	    RECT 192.7000 123.2000 194.5000 123.5000 ;
	    RECT 192.7000 123.1000 193.0000 123.2000 ;
	    RECT 192.6000 121.1000 193.0000 123.1000 ;
	    RECT 194.2000 123.1000 194.5000 123.2000 ;
	    RECT 194.2000 121.1000 194.6000 123.1000 ;
	    RECT 195.8000 121.1000 196.2000 125.4000 ;
	    RECT 199.1000 125.2000 199.4000 125.8000 ;
	    RECT 202.2000 125.5000 205.0000 125.6000 ;
	    RECT 202.1000 125.4000 205.0000 125.5000 ;
	    RECT 198.2000 124.9000 199.4000 125.2000 ;
	    RECT 200.1000 125.3000 205.0000 125.4000 ;
	    RECT 200.1000 125.1000 202.5000 125.3000 ;
	    RECT 198.2000 124.4000 198.5000 124.9000 ;
	    RECT 197.8000 124.0000 198.5000 124.4000 ;
	    RECT 199.3000 124.5000 199.7000 124.6000 ;
	    RECT 200.1000 124.5000 200.4000 125.1000 ;
	    RECT 199.3000 124.2000 200.4000 124.5000 ;
	    RECT 200.7000 124.5000 203.4000 124.8000 ;
	    RECT 200.7000 124.4000 201.1000 124.5000 ;
	    RECT 203.0000 124.4000 203.4000 124.5000 ;
	    RECT 199.9000 123.7000 200.3000 123.8000 ;
	    RECT 201.3000 123.7000 201.7000 123.8000 ;
	    RECT 198.2000 123.1000 198.6000 123.5000 ;
	    RECT 199.9000 123.4000 201.7000 123.7000 ;
	    RECT 200.3000 123.1000 200.6000 123.4000 ;
	    RECT 203.0000 123.1000 203.4000 123.5000 ;
	    RECT 197.9000 121.1000 198.5000 123.1000 ;
	    RECT 200.2000 121.1000 200.6000 123.1000 ;
	    RECT 202.4000 122.8000 203.4000 123.1000 ;
	    RECT 202.4000 121.1000 202.8000 122.8000 ;
	    RECT 204.6000 121.1000 205.0000 125.3000 ;
	    RECT 206.3000 125.1000 206.6000 126.8000 ;
	    RECT 207.0000 125.4000 207.4000 126.2000 ;
	    RECT 206.2000 124.7000 207.1000 125.1000 ;
	    RECT 206.7000 121.1000 207.1000 124.7000 ;
	    RECT 208.6000 121.1000 209.0000 129.9000 ;
	    RECT 209.4000 126.8000 209.8000 127.6000 ;
	    RECT 210.2000 126.1000 210.6000 129.9000 ;
	    RECT 213.4000 128.9000 213.8000 129.9000 ;
	    RECT 215.8000 128.9000 216.2000 129.9000 ;
	    RECT 211.0000 128.1000 211.4000 128.2000 ;
	    RECT 212.6000 128.1000 213.0000 128.6000 ;
	    RECT 211.0000 127.8000 213.0000 128.1000 ;
	    RECT 213.5000 127.2000 213.8000 128.9000 ;
	    RECT 215.0000 127.8000 215.4000 128.6000 ;
	    RECT 215.9000 127.2000 216.2000 128.9000 ;
	    RECT 217.5000 128.2000 217.9000 128.6000 ;
	    RECT 217.4000 127.8000 217.8000 128.2000 ;
	    RECT 218.2000 127.9000 218.6000 129.9000 ;
	    RECT 221.4000 128.9000 221.8000 129.9000 ;
	    RECT 223.8000 128.9000 224.2000 129.9000 ;
	    RECT 213.4000 127.1000 213.8000 127.2000 ;
	    RECT 215.0000 127.1000 215.4000 127.2000 ;
	    RECT 213.4000 126.8000 215.4000 127.1000 ;
	    RECT 215.8000 127.1000 216.2000 127.2000 ;
	    RECT 217.4000 127.1000 217.8000 127.2000 ;
	    RECT 215.8000 126.8000 217.8000 127.1000 ;
	    RECT 211.8000 126.1000 212.2000 126.2000 ;
	    RECT 210.2000 125.8000 212.2000 126.1000 ;
	    RECT 210.2000 121.1000 210.6000 125.8000 ;
	    RECT 213.5000 125.1000 213.8000 126.8000 ;
	    RECT 214.2000 125.4000 214.6000 126.2000 ;
	    RECT 215.9000 125.1000 216.2000 126.8000 ;
	    RECT 218.3000 126.2000 218.6000 127.9000 ;
	    RECT 220.6000 127.8000 221.0000 128.6000 ;
	    RECT 221.5000 127.2000 221.8000 128.9000 ;
	    RECT 223.0000 127.8000 223.4000 128.6000 ;
	    RECT 223.9000 127.2000 224.2000 128.9000 ;
	    RECT 226.7000 128.2000 227.1000 129.9000 ;
	    RECT 226.2000 127.9000 227.1000 128.2000 ;
	    RECT 219.0000 127.1000 219.4000 127.2000 ;
	    RECT 221.4000 127.1000 221.8000 127.2000 ;
	    RECT 219.0000 126.8000 221.8000 127.1000 ;
	    RECT 222.2000 127.1000 222.6000 127.2000 ;
	    RECT 223.8000 127.1000 224.2000 127.2000 ;
	    RECT 222.2000 126.8000 224.2000 127.1000 ;
	    RECT 225.4000 126.8000 225.8000 127.6000 ;
	    RECT 226.2000 127.1000 226.6000 127.9000 ;
	    RECT 227.8000 127.1000 228.2000 127.6000 ;
	    RECT 226.2000 126.8000 228.2000 127.1000 ;
	    RECT 219.0000 126.4000 219.4000 126.8000 ;
	    RECT 216.6000 125.4000 217.0000 126.2000 ;
	    RECT 217.4000 126.1000 217.8000 126.2000 ;
	    RECT 218.2000 126.1000 218.6000 126.2000 ;
	    RECT 219.8000 126.1000 220.2000 126.2000 ;
	    RECT 217.4000 125.8000 218.6000 126.1000 ;
	    RECT 219.4000 125.8000 220.2000 126.1000 ;
	    RECT 217.5000 125.1000 217.8000 125.8000 ;
	    RECT 219.4000 125.6000 219.8000 125.8000 ;
	    RECT 221.5000 125.1000 221.8000 126.8000 ;
	    RECT 222.2000 125.4000 222.6000 126.2000 ;
	    RECT 223.9000 125.1000 224.2000 126.8000 ;
	    RECT 224.6000 125.4000 225.0000 126.2000 ;
	    RECT 213.4000 124.7000 214.3000 125.1000 ;
	    RECT 215.8000 124.7000 216.7000 125.1000 ;
	    RECT 213.9000 121.1000 214.3000 124.7000 ;
	    RECT 216.3000 121.1000 216.7000 124.7000 ;
	    RECT 217.4000 121.1000 217.8000 125.1000 ;
	    RECT 218.2000 124.8000 220.2000 125.1000 ;
	    RECT 218.2000 121.1000 218.6000 124.8000 ;
	    RECT 219.8000 121.1000 220.2000 124.8000 ;
	    RECT 221.4000 124.7000 222.3000 125.1000 ;
	    RECT 223.8000 124.7000 224.7000 125.1000 ;
	    RECT 221.9000 121.1000 222.3000 124.7000 ;
	    RECT 224.3000 121.1000 224.7000 124.7000 ;
	    RECT 226.2000 121.1000 226.6000 126.8000 ;
	    RECT 227.0000 124.4000 227.4000 125.2000 ;
	    RECT 228.6000 121.1000 229.0000 129.9000 ;
	    RECT 230.2000 127.6000 230.6000 129.9000 ;
	    RECT 231.8000 127.6000 232.2000 129.9000 ;
	    RECT 234.2000 128.9000 234.6000 129.9000 ;
	    RECT 236.6000 128.9000 237.0000 129.9000 ;
	    RECT 230.2000 127.2000 232.2000 127.6000 ;
	    RECT 230.2000 125.8000 230.6000 127.2000 ;
	    RECT 232.6000 126.8000 233.0000 127.6000 ;
	    RECT 234.2000 127.2000 234.5000 128.9000 ;
	    RECT 235.0000 127.8000 235.4000 128.6000 ;
	    RECT 235.8000 127.8000 236.2000 128.6000 ;
	    RECT 236.7000 127.2000 237.0000 128.9000 ;
	    RECT 234.2000 126.8000 234.6000 127.2000 ;
	    RECT 236.6000 126.8000 237.0000 127.2000 ;
	    RECT 230.2000 125.4000 232.2000 125.8000 ;
	    RECT 233.4000 125.4000 233.8000 126.2000 ;
	    RECT 230.2000 121.1000 230.6000 125.4000 ;
	    RECT 231.8000 121.1000 232.2000 125.4000 ;
	    RECT 234.2000 125.1000 234.5000 126.8000 ;
	    RECT 236.7000 125.1000 237.0000 126.8000 ;
	    RECT 239.0000 127.1000 239.4000 129.9000 ;
	    RECT 239.8000 128.0000 240.2000 129.9000 ;
	    RECT 241.4000 128.0000 241.8000 129.9000 ;
	    RECT 239.8000 127.9000 241.8000 128.0000 ;
	    RECT 242.2000 127.9000 242.6000 129.9000 ;
	    RECT 239.9000 127.7000 241.7000 127.9000 ;
	    RECT 240.2000 127.2000 240.6000 127.4000 ;
	    RECT 242.2000 127.2000 242.5000 127.9000 ;
	    RECT 243.0000 127.8000 243.4000 128.6000 ;
	    RECT 239.8000 127.1000 240.6000 127.2000 ;
	    RECT 239.0000 126.9000 240.6000 127.1000 ;
	    RECT 239.0000 126.8000 240.2000 126.9000 ;
	    RECT 241.3000 126.8000 242.6000 127.2000 ;
	    RECT 237.4000 125.4000 237.8000 126.2000 ;
	    RECT 233.7000 124.7000 234.6000 125.1000 ;
	    RECT 236.6000 124.7000 237.5000 125.1000 ;
	    RECT 233.7000 122.2000 234.1000 124.7000 ;
	    RECT 237.1000 124.1000 237.5000 124.7000 ;
	    RECT 238.2000 124.1000 238.6000 124.2000 ;
	    RECT 237.1000 123.8000 238.6000 124.1000 ;
	    RECT 233.7000 121.8000 234.6000 122.2000 ;
	    RECT 233.7000 121.1000 234.1000 121.8000 ;
	    RECT 237.1000 121.1000 237.5000 123.8000 ;
	    RECT 239.0000 121.1000 239.4000 126.8000 ;
	    RECT 240.6000 125.8000 241.0000 126.6000 ;
	    RECT 241.3000 125.1000 241.6000 126.8000 ;
	    RECT 242.2000 125.1000 242.6000 125.2000 ;
	    RECT 243.0000 125.1000 243.4000 125.2000 ;
	    RECT 241.1000 124.8000 241.6000 125.1000 ;
	    RECT 241.9000 124.8000 243.4000 125.1000 ;
	    RECT 241.1000 123.2000 241.5000 124.8000 ;
	    RECT 241.9000 124.2000 242.2000 124.8000 ;
	    RECT 241.8000 123.8000 242.2000 124.2000 ;
	    RECT 240.6000 122.8000 241.5000 123.2000 ;
	    RECT 241.1000 121.1000 241.5000 122.8000 ;
	    RECT 243.8000 121.1000 244.2000 129.9000 ;
	    RECT 245.4000 128.8000 245.8000 129.9000 ;
	    RECT 245.4000 127.2000 245.7000 128.8000 ;
	    RECT 246.2000 128.1000 246.6000 128.6000 ;
	    RECT 247.0000 128.1000 247.4000 129.9000 ;
	    RECT 246.2000 127.8000 247.4000 128.1000 ;
	    RECT 245.4000 126.8000 245.8000 127.2000 ;
	    RECT 244.6000 125.4000 245.0000 126.2000 ;
	    RECT 245.4000 125.1000 245.7000 126.8000 ;
	    RECT 244.9000 124.7000 245.8000 125.1000 ;
	    RECT 244.9000 121.1000 245.3000 124.7000 ;
	    RECT 247.0000 121.1000 247.4000 127.8000 ;
	    RECT 249.4000 128.9000 249.8000 129.9000 ;
	    RECT 249.4000 127.2000 249.7000 128.9000 ;
	    RECT 251.0000 128.0000 251.4000 129.9000 ;
	    RECT 252.6000 128.0000 253.0000 129.9000 ;
	    RECT 251.0000 127.9000 253.0000 128.0000 ;
	    RECT 251.1000 127.7000 252.9000 127.9000 ;
	    RECT 253.4000 127.8000 253.8000 129.9000 ;
	    RECT 251.4000 127.2000 251.8000 127.4000 ;
	    RECT 253.4000 127.2000 253.7000 127.8000 ;
	    RECT 249.4000 126.8000 249.8000 127.2000 ;
	    RECT 251.0000 126.9000 251.8000 127.2000 ;
	    RECT 251.0000 126.8000 251.4000 126.9000 ;
	    RECT 252.5000 126.8000 253.8000 127.2000 ;
	    RECT 248.6000 125.4000 249.0000 126.2000 ;
	    RECT 249.4000 126.1000 249.7000 126.8000 ;
	    RECT 251.8000 126.1000 252.2000 126.6000 ;
	    RECT 249.4000 125.8000 252.2000 126.1000 ;
	    RECT 249.4000 125.1000 249.7000 125.8000 ;
	    RECT 252.5000 125.1000 252.8000 126.8000 ;
	    RECT 253.4000 125.1000 253.8000 125.2000 ;
	    RECT 254.2000 125.1000 254.6000 129.9000 ;
	    RECT 255.0000 127.8000 255.4000 128.6000 ;
	    RECT 255.9000 128.2000 256.3000 128.6000 ;
	    RECT 255.8000 127.8000 256.2000 128.2000 ;
	    RECT 256.6000 127.9000 257.0000 129.9000 ;
	    RECT 255.8000 126.1000 256.2000 126.2000 ;
	    RECT 256.7000 126.1000 257.0000 127.9000 ;
	    RECT 259.0000 127.8000 259.4000 128.6000 ;
	    RECT 257.4000 126.4000 257.8000 127.2000 ;
	    RECT 258.2000 126.1000 258.6000 126.2000 ;
	    RECT 255.8000 125.8000 257.0000 126.1000 ;
	    RECT 257.8000 125.8000 258.6000 126.1000 ;
	    RECT 259.8000 126.1000 260.2000 129.9000 ;
	    RECT 262.2000 127.9000 262.6000 129.9000 ;
	    RECT 262.9000 128.2000 263.3000 128.6000 ;
	    RECT 263.9000 128.2000 264.3000 128.6000 ;
	    RECT 261.4000 126.4000 261.8000 127.2000 ;
	    RECT 260.6000 126.1000 261.0000 126.2000 ;
	    RECT 262.2000 126.1000 262.5000 127.9000 ;
	    RECT 263.0000 127.8000 263.4000 128.2000 ;
	    RECT 263.8000 127.8000 264.2000 128.2000 ;
	    RECT 264.6000 127.9000 265.0000 129.9000 ;
	    RECT 267.3000 128.2000 267.7000 129.9000 ;
	    RECT 267.3000 127.9000 268.2000 128.2000 ;
	    RECT 263.0000 127.1000 263.3000 127.8000 ;
	    RECT 264.7000 127.1000 265.0000 127.9000 ;
	    RECT 263.0000 126.8000 265.0000 127.1000 ;
	    RECT 263.0000 126.1000 263.4000 126.2000 ;
	    RECT 259.8000 125.8000 261.4000 126.1000 ;
	    RECT 262.2000 125.8000 263.4000 126.1000 ;
	    RECT 263.8000 126.1000 264.2000 126.2000 ;
	    RECT 264.7000 126.1000 265.0000 126.8000 ;
	    RECT 265.4000 127.1000 265.8000 127.2000 ;
	    RECT 267.0000 127.1000 267.4000 127.2000 ;
	    RECT 265.4000 126.8000 267.4000 127.1000 ;
	    RECT 265.4000 126.4000 265.8000 126.8000 ;
	    RECT 266.2000 126.1000 266.6000 126.2000 ;
	    RECT 267.8000 126.1000 268.2000 127.9000 ;
	    RECT 263.8000 125.8000 265.0000 126.1000 ;
	    RECT 265.8000 125.8000 268.2000 126.1000 ;
	    RECT 255.9000 125.1000 256.2000 125.8000 ;
	    RECT 257.8000 125.6000 258.2000 125.8000 ;
	    RECT 248.9000 124.7000 249.8000 125.1000 ;
	    RECT 252.3000 124.8000 252.8000 125.1000 ;
	    RECT 253.1000 124.8000 254.6000 125.1000 ;
	    RECT 248.9000 121.1000 249.3000 124.7000 ;
	    RECT 252.3000 121.1000 252.7000 124.8000 ;
	    RECT 253.1000 124.2000 253.4000 124.8000 ;
	    RECT 253.0000 123.8000 253.4000 124.2000 ;
	    RECT 254.2000 121.1000 254.6000 124.8000 ;
	    RECT 255.8000 121.1000 256.2000 125.1000 ;
	    RECT 256.6000 124.8000 258.6000 125.1000 ;
	    RECT 256.6000 121.1000 257.0000 124.8000 ;
	    RECT 258.2000 121.1000 258.6000 124.8000 ;
	    RECT 259.8000 121.1000 260.2000 125.8000 ;
	    RECT 261.0000 125.6000 261.4000 125.8000 ;
	    RECT 263.0000 125.1000 263.3000 125.8000 ;
	    RECT 263.9000 125.1000 264.2000 125.8000 ;
	    RECT 265.8000 125.6000 266.2000 125.8000 ;
	    RECT 260.6000 124.8000 262.6000 125.1000 ;
	    RECT 260.6000 121.1000 261.0000 124.8000 ;
	    RECT 262.2000 121.1000 262.6000 124.8000 ;
	    RECT 263.0000 121.1000 263.4000 125.1000 ;
	    RECT 263.8000 121.1000 264.2000 125.1000 ;
	    RECT 264.6000 124.8000 266.6000 125.1000 ;
	    RECT 264.6000 121.1000 265.0000 124.8000 ;
	    RECT 266.2000 121.1000 266.6000 124.8000 ;
	    RECT 267.0000 124.4000 267.4000 125.2000 ;
	    RECT 267.8000 121.1000 268.2000 125.8000 ;
	    RECT 1.4000 115.1000 1.8000 119.9000 ;
	    RECT 2.5000 116.3000 2.9000 119.9000 ;
	    RECT 2.5000 115.9000 3.4000 116.3000 ;
	    RECT 4.6000 116.2000 5.0000 119.9000 ;
	    RECT 6.2000 116.2000 6.6000 119.9000 ;
	    RECT 4.6000 115.9000 6.6000 116.2000 ;
	    RECT 7.0000 115.9000 7.4000 119.9000 ;
	    RECT 9.1000 116.3000 9.5000 119.9000 ;
	    RECT 8.6000 115.9000 9.5000 116.3000 ;
	    RECT 2.2000 115.1000 2.6000 115.6000 ;
	    RECT 1.4000 114.8000 2.6000 115.1000 ;
	    RECT 3.0000 115.1000 3.3000 115.9000 ;
	    RECT 5.0000 115.2000 5.4000 115.4000 ;
	    RECT 7.0000 115.2000 7.3000 115.9000 ;
	    RECT 4.6000 115.1000 5.4000 115.2000 ;
	    RECT 3.0000 114.9000 5.4000 115.1000 ;
	    RECT 6.2000 114.9000 7.4000 115.2000 ;
	    RECT 3.0000 114.8000 5.0000 114.9000 ;
	    RECT 1.4000 111.1000 1.8000 114.8000 ;
	    RECT 3.0000 114.2000 3.3000 114.8000 ;
	    RECT 3.0000 113.8000 3.4000 114.2000 ;
	    RECT 5.4000 113.8000 5.8000 114.6000 ;
	    RECT 3.0000 112.1000 3.3000 113.8000 ;
	    RECT 6.2000 113.1000 6.5000 114.9000 ;
	    RECT 7.0000 114.8000 7.4000 114.9000 ;
	    RECT 8.7000 114.2000 9.0000 115.9000 ;
	    RECT 9.4000 115.1000 9.8000 115.6000 ;
	    RECT 10.2000 115.1000 10.6000 119.9000 ;
	    RECT 11.8000 116.2000 12.2000 119.9000 ;
	    RECT 12.6000 116.2000 13.0000 116.3000 ;
	    RECT 14.0000 116.2000 14.8000 119.9000 ;
	    RECT 11.8000 115.9000 13.0000 116.2000 ;
	    RECT 13.8000 115.9000 14.8000 116.2000 ;
	    RECT 15.9000 116.2000 16.3000 116.3000 ;
	    RECT 16.6000 116.2000 17.0000 119.9000 ;
	    RECT 18.7000 119.2000 19.1000 119.9000 ;
	    RECT 18.2000 118.8000 19.1000 119.2000 ;
	    RECT 15.9000 115.9000 17.0000 116.2000 ;
	    RECT 18.7000 116.2000 19.1000 118.8000 ;
	    RECT 19.4000 116.8000 19.8000 117.2000 ;
	    RECT 19.5000 116.2000 19.8000 116.8000 ;
	    RECT 18.7000 115.9000 19.2000 116.2000 ;
	    RECT 19.5000 115.9000 20.2000 116.2000 ;
	    RECT 13.8000 115.2000 14.1000 115.9000 ;
	    RECT 15.9000 115.6000 16.2000 115.9000 ;
	    RECT 14.5000 115.3000 16.2000 115.6000 ;
	    RECT 14.5000 115.2000 14.9000 115.3000 ;
	    RECT 9.4000 114.8000 10.6000 115.1000 ;
	    RECT 11.0000 115.1000 11.4000 115.2000 ;
	    RECT 13.4000 115.1000 14.1000 115.2000 ;
	    RECT 11.0000 114.9000 14.1000 115.1000 ;
	    RECT 15.6000 114.9000 16.0000 115.0000 ;
	    RECT 11.0000 114.8000 14.3000 114.9000 ;
	    RECT 8.6000 114.1000 9.0000 114.2000 ;
	    RECT 7.0000 113.8000 9.0000 114.1000 ;
	    RECT 7.0000 113.2000 7.3000 113.8000 ;
	    RECT 3.0000 111.1000 3.4000 112.1000 ;
	    RECT 6.2000 111.1000 6.6000 113.1000 ;
	    RECT 7.0000 112.8000 7.4000 113.2000 ;
	    RECT 6.9000 112.4000 7.3000 112.8000 ;
	    RECT 8.7000 112.1000 9.0000 113.8000 ;
	    RECT 8.6000 111.1000 9.0000 112.1000 ;
	    RECT 10.2000 111.1000 10.6000 114.8000 ;
	    RECT 13.8000 114.6000 14.3000 114.8000 ;
	    RECT 12.6000 113.4000 13.0000 113.5000 ;
	    RECT 11.8000 113.1000 13.0000 113.4000 ;
	    RECT 11.8000 111.1000 12.2000 113.1000 ;
	    RECT 14.0000 112.9000 14.3000 114.6000 ;
	    RECT 14.7000 114.6000 16.0000 114.9000 ;
	    RECT 14.7000 114.3000 15.0000 114.6000 ;
	    RECT 18.2000 114.4000 18.6000 115.2000 ;
	    RECT 14.6000 113.9000 15.0000 114.3000 ;
	    RECT 18.9000 114.2000 19.2000 115.9000 ;
	    RECT 19.8000 115.8000 20.2000 115.9000 ;
	    RECT 17.4000 114.1000 17.8000 114.2000 ;
	    RECT 17.4000 113.8000 18.2000 114.1000 ;
	    RECT 18.9000 113.8000 20.2000 114.2000 ;
	    RECT 17.8000 113.6000 18.2000 113.8000 ;
	    RECT 15.9000 113.4000 16.3000 113.5000 ;
	    RECT 15.9000 113.1000 17.0000 113.4000 ;
	    RECT 17.5000 113.1000 19.3000 113.3000 ;
	    RECT 19.8000 113.1000 20.1000 113.8000 ;
	    RECT 20.6000 113.4000 21.0000 114.2000 ;
	    RECT 21.4000 113.1000 21.8000 119.9000 ;
	    RECT 23.8000 117.9000 24.2000 119.9000 ;
	    RECT 22.2000 115.8000 22.6000 116.6000 ;
	    RECT 23.9000 115.8000 24.2000 117.9000 ;
	    RECT 25.4000 115.9000 25.8000 119.9000 ;
	    RECT 27.5000 119.2000 27.9000 119.9000 ;
	    RECT 27.0000 118.8000 27.9000 119.2000 ;
	    RECT 27.5000 116.2000 27.9000 118.8000 ;
	    RECT 30.7000 117.2000 31.1000 119.9000 ;
	    RECT 32.6000 119.6000 34.6000 119.9000 ;
	    RECT 28.2000 116.8000 28.6000 117.2000 ;
	    RECT 30.2000 116.8000 31.1000 117.2000 ;
	    RECT 31.4000 116.8000 31.8000 117.2000 ;
	    RECT 28.3000 116.2000 28.6000 116.8000 ;
	    RECT 30.7000 116.2000 31.1000 116.8000 ;
	    RECT 31.5000 116.2000 31.8000 116.8000 ;
	    RECT 27.5000 115.9000 28.0000 116.2000 ;
	    RECT 28.3000 115.9000 29.0000 116.2000 ;
	    RECT 30.7000 115.9000 31.2000 116.2000 ;
	    RECT 31.5000 115.9000 32.2000 116.2000 ;
	    RECT 32.6000 115.9000 33.0000 119.6000 ;
	    RECT 33.4000 115.9000 33.8000 119.3000 ;
	    RECT 34.2000 116.2000 34.6000 119.6000 ;
	    RECT 35.8000 116.2000 36.2000 119.9000 ;
	    RECT 34.2000 115.9000 36.2000 116.2000 ;
	    RECT 23.9000 115.5000 25.1000 115.8000 ;
	    RECT 23.8000 114.8000 24.2000 115.2000 ;
	    RECT 22.2000 114.1000 22.6000 114.2000 ;
	    RECT 23.0000 114.1000 23.4000 114.6000 ;
	    RECT 23.9000 114.4000 24.2000 114.8000 ;
	    RECT 23.9000 114.1000 24.4000 114.4000 ;
	    RECT 22.2000 113.8000 23.4000 114.1000 ;
	    RECT 24.0000 114.0000 24.4000 114.1000 ;
	    RECT 24.8000 113.8000 25.1000 115.5000 ;
	    RECT 25.5000 115.2000 25.8000 115.9000 ;
	    RECT 25.4000 114.8000 25.8000 115.2000 ;
	    RECT 24.8000 113.7000 25.2000 113.8000 ;
	    RECT 23.7000 113.5000 25.2000 113.7000 ;
	    RECT 23.1000 113.4000 25.2000 113.5000 ;
	    RECT 23.1000 113.2000 24.0000 113.4000 ;
	    RECT 23.1000 113.1000 23.4000 113.2000 ;
	    RECT 25.5000 113.1000 25.8000 114.8000 ;
	    RECT 27.0000 114.4000 27.4000 115.2000 ;
	    RECT 27.7000 114.2000 28.0000 115.9000 ;
	    RECT 28.6000 115.8000 29.0000 115.9000 ;
	    RECT 30.2000 114.4000 30.6000 115.2000 ;
	    RECT 30.9000 114.2000 31.2000 115.9000 ;
	    RECT 31.8000 115.8000 32.2000 115.9000 ;
	    RECT 33.5000 115.6000 33.8000 115.9000 ;
	    RECT 36.6000 115.7000 37.0000 119.9000 ;
	    RECT 38.8000 118.2000 39.2000 119.9000 ;
	    RECT 38.2000 117.9000 39.2000 118.2000 ;
	    RECT 41.0000 117.9000 41.4000 119.9000 ;
	    RECT 43.1000 117.9000 43.7000 119.9000 ;
	    RECT 38.2000 117.5000 38.6000 117.9000 ;
	    RECT 41.0000 117.6000 41.3000 117.9000 ;
	    RECT 39.9000 117.3000 41.7000 117.6000 ;
	    RECT 43.0000 117.5000 43.4000 117.9000 ;
	    RECT 39.9000 117.2000 40.3000 117.3000 ;
	    RECT 41.3000 117.2000 41.7000 117.3000 ;
	    RECT 45.4000 117.1000 45.8000 119.9000 ;
	    RECT 46.2000 117.1000 46.6000 117.2000 ;
	    RECT 38.2000 116.5000 38.6000 116.6000 ;
	    RECT 40.5000 116.5000 40.9000 116.6000 ;
	    RECT 38.2000 116.2000 40.9000 116.5000 ;
	    RECT 41.2000 116.5000 42.3000 116.8000 ;
	    RECT 41.2000 115.9000 41.5000 116.5000 ;
	    RECT 41.9000 116.4000 42.3000 116.5000 ;
	    RECT 43.1000 116.6000 43.8000 117.0000 ;
	    RECT 45.4000 116.8000 46.6000 117.1000 ;
	    RECT 43.1000 116.1000 43.4000 116.6000 ;
	    RECT 39.1000 115.7000 41.5000 115.9000 ;
	    RECT 36.6000 115.6000 41.5000 115.7000 ;
	    RECT 42.2000 115.8000 43.4000 116.1000 ;
	    RECT 31.8000 115.1000 32.2000 115.2000 ;
	    RECT 32.6000 115.1000 33.0000 115.6000 ;
	    RECT 33.5000 115.3000 34.5000 115.6000 ;
	    RECT 36.6000 115.5000 39.5000 115.6000 ;
	    RECT 36.6000 115.4000 39.4000 115.5000 ;
	    RECT 31.8000 114.8000 33.0000 115.1000 ;
	    RECT 34.2000 115.2000 34.5000 115.3000 ;
	    RECT 35.4000 115.2000 35.8000 115.4000 ;
	    RECT 42.2000 115.2000 42.5000 115.8000 ;
	    RECT 45.4000 115.6000 45.8000 116.8000 ;
	    RECT 43.7000 115.3000 45.8000 115.6000 ;
	    RECT 43.7000 115.2000 44.1000 115.3000 ;
	    RECT 34.2000 114.8000 34.6000 115.2000 ;
	    RECT 35.4000 114.9000 36.2000 115.2000 ;
	    RECT 39.8000 115.1000 40.2000 115.2000 ;
	    RECT 35.8000 114.8000 36.2000 114.9000 ;
	    RECT 37.7000 114.8000 40.2000 115.1000 ;
	    RECT 42.2000 114.8000 42.6000 115.2000 ;
	    RECT 44.5000 114.9000 44.9000 115.0000 ;
	    RECT 33.5000 114.4000 33.9000 114.8000 ;
	    RECT 33.5000 114.2000 33.8000 114.4000 ;
	    RECT 26.2000 114.1000 26.6000 114.2000 ;
	    RECT 26.2000 113.8000 27.0000 114.1000 ;
	    RECT 27.7000 113.8000 29.0000 114.2000 ;
	    RECT 29.4000 114.1000 29.8000 114.2000 ;
	    RECT 29.4000 113.8000 30.2000 114.1000 ;
	    RECT 30.9000 113.8000 32.2000 114.2000 ;
	    RECT 33.4000 113.8000 33.8000 114.2000 ;
	    RECT 26.6000 113.6000 27.0000 113.8000 ;
	    RECT 26.3000 113.1000 28.1000 113.3000 ;
	    RECT 28.6000 113.1000 28.9000 113.8000 ;
	    RECT 29.8000 113.6000 30.2000 113.8000 ;
	    RECT 29.5000 113.1000 31.3000 113.3000 ;
	    RECT 31.8000 113.1000 32.1000 113.8000 ;
	    RECT 34.2000 113.1000 34.5000 114.8000 ;
	    RECT 37.7000 114.7000 38.1000 114.8000 ;
	    RECT 39.0000 114.7000 39.4000 114.8000 ;
	    RECT 35.0000 113.8000 35.4000 114.6000 ;
	    RECT 38.5000 114.2000 38.9000 114.3000 ;
	    RECT 42.2000 114.2000 42.5000 114.8000 ;
	    RECT 43.0000 114.6000 44.9000 114.9000 ;
	    RECT 43.0000 114.5000 43.4000 114.6000 ;
	    RECT 37.0000 113.9000 42.5000 114.2000 ;
	    RECT 37.0000 113.8000 37.8000 113.9000 ;
	    RECT 14.0000 111.1000 14.8000 112.9000 ;
	    RECT 16.6000 111.1000 17.0000 113.1000 ;
	    RECT 17.4000 113.0000 19.4000 113.1000 ;
	    RECT 17.4000 111.1000 17.8000 113.0000 ;
	    RECT 19.0000 111.1000 19.4000 113.0000 ;
	    RECT 19.8000 111.1000 20.2000 113.1000 ;
	    RECT 21.4000 112.8000 22.3000 113.1000 ;
	    RECT 21.9000 111.1000 22.3000 112.8000 ;
	    RECT 23.0000 111.1000 23.4000 113.1000 ;
	    RECT 25.1000 112.6000 25.8000 113.1000 ;
	    RECT 26.2000 113.0000 28.2000 113.1000 ;
	    RECT 25.1000 112.2000 25.5000 112.6000 ;
	    RECT 25.1000 111.8000 25.8000 112.2000 ;
	    RECT 25.1000 111.1000 25.5000 111.8000 ;
	    RECT 26.2000 111.1000 26.6000 113.0000 ;
	    RECT 27.8000 111.1000 28.2000 113.0000 ;
	    RECT 28.6000 111.1000 29.0000 113.1000 ;
	    RECT 29.4000 113.0000 31.4000 113.1000 ;
	    RECT 29.4000 111.1000 29.8000 113.0000 ;
	    RECT 31.0000 111.1000 31.4000 113.0000 ;
	    RECT 31.8000 111.1000 32.2000 113.1000 ;
	    RECT 33.9000 111.1000 34.7000 113.1000 ;
	    RECT 36.6000 111.1000 37.0000 113.5000 ;
	    RECT 39.1000 112.8000 39.4000 113.9000 ;
	    RECT 41.9000 113.8000 42.3000 113.9000 ;
	    RECT 45.4000 113.6000 45.8000 115.3000 ;
	    RECT 43.9000 113.3000 45.8000 113.6000 ;
	    RECT 46.2000 113.4000 46.6000 114.2000 ;
	    RECT 47.0000 114.1000 47.4000 119.9000 ;
	    RECT 47.8000 116.1000 48.2000 116.6000 ;
	    RECT 48.6000 116.1000 49.0000 119.9000 ;
	    RECT 47.8000 115.8000 49.0000 116.1000 ;
	    RECT 47.8000 114.1000 48.2000 114.2000 ;
	    RECT 47.0000 113.8000 48.2000 114.1000 ;
	    RECT 43.9000 113.2000 44.3000 113.3000 ;
	    RECT 38.2000 112.1000 38.6000 112.5000 ;
	    RECT 39.0000 112.4000 39.4000 112.8000 ;
	    RECT 39.9000 112.7000 40.3000 112.8000 ;
	    RECT 39.9000 112.4000 41.3000 112.7000 ;
	    RECT 41.0000 112.1000 41.3000 112.4000 ;
	    RECT 43.0000 112.1000 43.4000 112.5000 ;
	    RECT 38.2000 111.8000 39.2000 112.1000 ;
	    RECT 38.8000 111.1000 39.2000 111.8000 ;
	    RECT 41.0000 111.1000 41.4000 112.1000 ;
	    RECT 43.0000 111.8000 43.7000 112.1000 ;
	    RECT 43.1000 111.1000 43.7000 111.8000 ;
	    RECT 45.4000 111.1000 45.8000 113.3000 ;
	    RECT 47.0000 113.1000 47.4000 113.8000 ;
	    RECT 47.0000 112.8000 47.9000 113.1000 ;
	    RECT 47.5000 111.1000 47.9000 112.8000 ;
	    RECT 48.6000 111.1000 49.0000 115.8000 ;
	    RECT 50.2000 115.7000 50.6000 119.9000 ;
	    RECT 52.4000 118.2000 52.8000 119.9000 ;
	    RECT 51.8000 117.9000 52.8000 118.2000 ;
	    RECT 54.6000 117.9000 55.0000 119.9000 ;
	    RECT 56.7000 117.9000 57.3000 119.9000 ;
	    RECT 51.8000 117.5000 52.2000 117.9000 ;
	    RECT 54.6000 117.6000 54.9000 117.9000 ;
	    RECT 53.5000 117.3000 55.3000 117.6000 ;
	    RECT 56.6000 117.5000 57.0000 117.9000 ;
	    RECT 53.5000 117.2000 53.9000 117.3000 ;
	    RECT 54.9000 117.2000 55.3000 117.3000 ;
	    RECT 51.8000 116.5000 52.2000 116.6000 ;
	    RECT 54.1000 116.5000 54.5000 116.6000 ;
	    RECT 51.8000 116.2000 54.5000 116.5000 ;
	    RECT 54.8000 116.5000 55.9000 116.8000 ;
	    RECT 54.8000 115.9000 55.1000 116.5000 ;
	    RECT 55.5000 116.4000 55.9000 116.5000 ;
	    RECT 56.7000 116.6000 57.4000 117.0000 ;
	    RECT 56.7000 116.1000 57.0000 116.6000 ;
	    RECT 52.7000 115.7000 55.1000 115.9000 ;
	    RECT 50.2000 115.6000 55.1000 115.7000 ;
	    RECT 55.8000 115.8000 57.0000 116.1000 ;
	    RECT 50.2000 115.5000 53.1000 115.6000 ;
	    RECT 50.2000 115.4000 53.0000 115.5000 ;
	    RECT 55.8000 115.2000 56.1000 115.8000 ;
	    RECT 59.0000 115.6000 59.4000 119.9000 ;
	    RECT 61.7000 116.2000 62.1000 119.9000 ;
	    RECT 57.3000 115.3000 59.4000 115.6000 ;
	    RECT 57.3000 115.2000 57.7000 115.3000 ;
	    RECT 53.4000 115.1000 53.8000 115.2000 ;
	    RECT 51.3000 114.8000 53.8000 115.1000 ;
	    RECT 55.8000 114.8000 56.2000 115.2000 ;
	    RECT 58.1000 114.9000 58.5000 115.0000 ;
	    RECT 51.3000 114.7000 51.7000 114.8000 ;
	    RECT 52.1000 114.2000 52.5000 114.3000 ;
	    RECT 55.8000 114.2000 56.1000 114.8000 ;
	    RECT 56.6000 114.6000 58.5000 114.9000 ;
	    RECT 56.6000 114.5000 57.0000 114.6000 ;
	    RECT 50.6000 113.9000 56.1000 114.2000 ;
	    RECT 50.6000 113.8000 51.4000 113.9000 ;
	    RECT 49.4000 112.4000 49.8000 113.2000 ;
	    RECT 50.2000 111.1000 50.6000 113.5000 ;
	    RECT 52.7000 112.8000 53.0000 113.9000 ;
	    RECT 55.5000 113.8000 55.9000 113.9000 ;
	    RECT 59.0000 113.6000 59.4000 115.3000 ;
	    RECT 61.4000 115.9000 62.1000 116.2000 ;
	    RECT 61.4000 115.2000 61.7000 115.9000 ;
	    RECT 63.8000 115.6000 64.2000 119.9000 ;
	    RECT 62.2000 115.4000 64.2000 115.6000 ;
	    RECT 64.6000 115.7000 65.0000 119.9000 ;
	    RECT 66.8000 118.2000 67.2000 119.9000 ;
	    RECT 66.2000 117.9000 67.2000 118.2000 ;
	    RECT 69.0000 117.9000 69.4000 119.9000 ;
	    RECT 71.1000 117.9000 71.7000 119.9000 ;
	    RECT 66.2000 117.5000 66.6000 117.9000 ;
	    RECT 69.0000 117.6000 69.3000 117.9000 ;
	    RECT 67.9000 117.3000 69.7000 117.6000 ;
	    RECT 71.0000 117.5000 71.4000 117.9000 ;
	    RECT 67.9000 117.2000 68.3000 117.3000 ;
	    RECT 69.3000 117.2000 69.7000 117.3000 ;
	    RECT 73.4000 117.1000 73.8000 119.9000 ;
	    RECT 75.0000 117.9000 75.4000 119.9000 ;
	    RECT 75.1000 117.8000 75.4000 117.9000 ;
	    RECT 76.6000 117.9000 77.0000 119.9000 ;
	    RECT 76.6000 117.8000 76.9000 117.9000 ;
	    RECT 75.1000 117.5000 76.9000 117.8000 ;
	    RECT 66.2000 116.5000 66.6000 116.6000 ;
	    RECT 68.5000 116.5000 68.9000 116.6000 ;
	    RECT 66.2000 116.2000 68.9000 116.5000 ;
	    RECT 69.2000 116.5000 70.3000 116.8000 ;
	    RECT 69.2000 115.9000 69.5000 116.5000 ;
	    RECT 69.9000 116.4000 70.3000 116.5000 ;
	    RECT 71.1000 116.6000 71.8000 117.0000 ;
	    RECT 73.4000 116.8000 74.5000 117.1000 ;
	    RECT 71.1000 116.1000 71.4000 116.6000 ;
	    RECT 67.1000 115.7000 69.5000 115.9000 ;
	    RECT 64.6000 115.6000 69.5000 115.7000 ;
	    RECT 70.2000 115.8000 71.4000 116.1000 ;
	    RECT 64.6000 115.5000 67.5000 115.6000 ;
	    RECT 64.6000 115.4000 67.4000 115.5000 ;
	    RECT 62.1000 115.3000 64.2000 115.4000 ;
	    RECT 60.6000 115.1000 61.0000 115.2000 ;
	    RECT 61.4000 115.1000 61.8000 115.2000 ;
	    RECT 60.6000 114.8000 61.8000 115.1000 ;
	    RECT 62.1000 115.0000 62.5000 115.3000 ;
	    RECT 70.2000 115.2000 70.5000 115.8000 ;
	    RECT 73.4000 115.6000 73.8000 116.8000 ;
	    RECT 71.7000 115.3000 73.8000 115.6000 ;
	    RECT 74.2000 116.2000 74.5000 116.8000 ;
	    RECT 75.8000 116.4000 76.2000 117.2000 ;
	    RECT 76.6000 116.2000 76.9000 117.5000 ;
	    RECT 74.2000 115.4000 74.6000 116.2000 ;
	    RECT 76.6000 115.8000 77.0000 116.2000 ;
	    RECT 71.7000 115.2000 72.1000 115.3000 ;
	    RECT 67.8000 115.1000 68.2000 115.2000 ;
	    RECT 57.5000 113.3000 59.4000 113.6000 ;
	    RECT 57.5000 113.2000 57.9000 113.3000 ;
	    RECT 51.8000 112.1000 52.2000 112.5000 ;
	    RECT 52.6000 112.4000 53.0000 112.8000 ;
	    RECT 53.5000 112.7000 53.9000 112.8000 ;
	    RECT 53.5000 112.4000 54.9000 112.7000 ;
	    RECT 54.6000 112.1000 54.9000 112.4000 ;
	    RECT 56.6000 112.1000 57.0000 112.5000 ;
	    RECT 51.8000 111.8000 52.8000 112.1000 ;
	    RECT 52.4000 111.1000 52.8000 111.8000 ;
	    RECT 54.6000 111.1000 55.0000 112.1000 ;
	    RECT 56.6000 111.8000 57.3000 112.1000 ;
	    RECT 56.7000 111.1000 57.3000 111.8000 ;
	    RECT 59.0000 111.1000 59.4000 113.3000 ;
	    RECT 61.4000 113.1000 61.7000 114.8000 ;
	    RECT 62.1000 113.5000 62.4000 115.0000 ;
	    RECT 65.7000 114.8000 68.2000 115.1000 ;
	    RECT 70.2000 114.8000 70.6000 115.2000 ;
	    RECT 72.5000 114.9000 72.9000 115.0000 ;
	    RECT 65.7000 114.7000 66.1000 114.8000 ;
	    RECT 62.8000 114.2000 63.2000 114.6000 ;
	    RECT 66.5000 114.2000 66.9000 114.3000 ;
	    RECT 70.2000 114.2000 70.5000 114.8000 ;
	    RECT 71.0000 114.6000 72.9000 114.9000 ;
	    RECT 71.0000 114.5000 71.4000 114.6000 ;
	    RECT 62.9000 113.8000 63.4000 114.2000 ;
	    RECT 65.0000 113.9000 70.5000 114.2000 ;
	    RECT 65.0000 113.8000 65.8000 113.9000 ;
	    RECT 62.1000 113.2000 63.3000 113.5000 ;
	    RECT 61.4000 111.1000 61.8000 113.1000 ;
	    RECT 63.0000 112.1000 63.3000 113.2000 ;
	    RECT 63.8000 112.4000 64.2000 113.2000 ;
	    RECT 63.0000 111.1000 63.4000 112.1000 ;
	    RECT 64.6000 111.1000 65.0000 113.5000 ;
	    RECT 67.1000 112.8000 67.4000 113.9000 ;
	    RECT 69.9000 113.8000 70.3000 113.9000 ;
	    RECT 73.4000 113.6000 73.8000 115.3000 ;
	    RECT 75.0000 114.8000 75.8000 115.2000 ;
	    RECT 76.6000 114.2000 76.9000 115.8000 ;
	    RECT 76.1000 114.1000 76.9000 114.2000 ;
	    RECT 71.9000 113.3000 73.8000 113.6000 ;
	    RECT 71.9000 113.2000 72.3000 113.3000 ;
	    RECT 66.2000 112.1000 66.6000 112.5000 ;
	    RECT 67.0000 112.4000 67.4000 112.8000 ;
	    RECT 67.9000 112.7000 68.3000 112.8000 ;
	    RECT 67.9000 112.4000 69.3000 112.7000 ;
	    RECT 69.0000 112.1000 69.3000 112.4000 ;
	    RECT 71.0000 112.1000 71.4000 112.5000 ;
	    RECT 66.2000 111.8000 67.2000 112.1000 ;
	    RECT 66.8000 111.1000 67.2000 111.8000 ;
	    RECT 69.0000 111.1000 69.4000 112.1000 ;
	    RECT 71.0000 111.8000 71.7000 112.1000 ;
	    RECT 71.1000 111.1000 71.7000 111.8000 ;
	    RECT 73.4000 111.1000 73.8000 113.3000 ;
	    RECT 76.0000 113.9000 76.9000 114.1000 ;
	    RECT 77.4000 115.6000 77.8000 119.9000 ;
	    RECT 79.5000 117.9000 80.1000 119.9000 ;
	    RECT 81.8000 117.9000 82.2000 119.9000 ;
	    RECT 84.0000 118.2000 84.4000 119.9000 ;
	    RECT 84.0000 117.9000 85.0000 118.2000 ;
	    RECT 79.8000 117.5000 80.2000 117.9000 ;
	    RECT 81.9000 117.6000 82.2000 117.9000 ;
	    RECT 81.5000 117.3000 83.3000 117.6000 ;
	    RECT 84.6000 117.5000 85.0000 117.9000 ;
	    RECT 81.5000 117.2000 81.9000 117.3000 ;
	    RECT 82.9000 117.2000 83.3000 117.3000 ;
	    RECT 79.4000 116.6000 80.1000 117.0000 ;
	    RECT 79.8000 116.1000 80.1000 116.6000 ;
	    RECT 80.9000 116.5000 82.0000 116.8000 ;
	    RECT 80.9000 116.4000 81.3000 116.5000 ;
	    RECT 79.8000 115.8000 81.0000 116.1000 ;
	    RECT 77.4000 115.3000 79.5000 115.6000 ;
	    RECT 76.0000 111.1000 76.4000 113.9000 ;
	    RECT 77.4000 113.6000 77.8000 115.3000 ;
	    RECT 79.1000 115.2000 79.5000 115.3000 ;
	    RECT 78.3000 114.9000 78.7000 115.0000 ;
	    RECT 78.3000 114.6000 80.2000 114.9000 ;
	    RECT 79.8000 114.5000 80.2000 114.6000 ;
	    RECT 80.7000 114.2000 81.0000 115.8000 ;
	    RECT 81.7000 115.9000 82.0000 116.5000 ;
	    RECT 82.3000 116.5000 82.7000 116.6000 ;
	    RECT 84.6000 116.5000 85.0000 116.6000 ;
	    RECT 82.3000 116.2000 85.0000 116.5000 ;
	    RECT 81.7000 115.7000 84.1000 115.9000 ;
	    RECT 86.2000 115.7000 86.6000 119.9000 ;
	    RECT 87.3000 116.3000 87.7000 119.9000 ;
	    RECT 87.3000 115.9000 88.2000 116.3000 ;
	    RECT 81.7000 115.6000 86.6000 115.7000 ;
	    RECT 83.7000 115.5000 86.6000 115.6000 ;
	    RECT 83.8000 115.4000 86.6000 115.5000 ;
	    RECT 83.0000 115.1000 83.4000 115.2000 ;
	    RECT 83.0000 114.8000 85.5000 115.1000 ;
	    RECT 87.0000 114.8000 87.4000 115.6000 ;
	    RECT 87.8000 115.1000 88.1000 115.9000 ;
	    RECT 89.4000 115.7000 89.8000 119.9000 ;
	    RECT 91.6000 118.2000 92.0000 119.9000 ;
	    RECT 91.0000 117.9000 92.0000 118.2000 ;
	    RECT 93.8000 117.9000 94.2000 119.9000 ;
	    RECT 95.9000 117.9000 96.5000 119.9000 ;
	    RECT 91.0000 117.5000 91.4000 117.9000 ;
	    RECT 93.8000 117.6000 94.1000 117.9000 ;
	    RECT 92.7000 117.3000 94.5000 117.6000 ;
	    RECT 95.8000 117.5000 96.2000 117.9000 ;
	    RECT 92.7000 117.2000 93.1000 117.3000 ;
	    RECT 94.1000 117.2000 94.5000 117.3000 ;
	    RECT 91.0000 116.5000 91.4000 116.6000 ;
	    RECT 93.3000 116.5000 93.7000 116.6000 ;
	    RECT 91.0000 116.2000 93.7000 116.5000 ;
	    RECT 94.0000 116.5000 95.1000 116.8000 ;
	    RECT 94.0000 115.9000 94.3000 116.5000 ;
	    RECT 94.7000 116.4000 95.1000 116.5000 ;
	    RECT 95.9000 116.6000 96.6000 117.0000 ;
	    RECT 95.9000 116.1000 96.2000 116.6000 ;
	    RECT 91.9000 115.7000 94.3000 115.9000 ;
	    RECT 89.4000 115.6000 94.3000 115.7000 ;
	    RECT 95.0000 115.8000 96.2000 116.1000 ;
	    RECT 89.4000 115.5000 92.3000 115.6000 ;
	    RECT 89.4000 115.4000 92.2000 115.5000 ;
	    RECT 92.6000 115.1000 93.0000 115.2000 ;
	    RECT 87.8000 114.8000 88.9000 115.1000 ;
	    RECT 85.1000 114.7000 85.5000 114.8000 ;
	    RECT 84.3000 114.2000 84.7000 114.3000 ;
	    RECT 87.8000 114.2000 88.1000 114.8000 ;
	    RECT 88.6000 114.2000 88.9000 114.8000 ;
	    RECT 90.5000 114.8000 93.0000 115.1000 ;
	    RECT 90.5000 114.7000 90.9000 114.8000 ;
	    RECT 91.8000 114.7000 92.2000 114.8000 ;
	    RECT 91.3000 114.2000 91.7000 114.3000 ;
	    RECT 95.0000 114.2000 95.3000 115.8000 ;
	    RECT 98.2000 115.6000 98.6000 119.9000 ;
	    RECT 96.5000 115.3000 98.6000 115.6000 ;
	    RECT 96.5000 115.2000 96.9000 115.3000 ;
	    RECT 97.3000 114.9000 97.7000 115.0000 ;
	    RECT 95.8000 114.6000 97.7000 114.9000 ;
	    RECT 95.8000 114.5000 96.2000 114.6000 ;
	    RECT 80.7000 113.9000 86.2000 114.2000 ;
	    RECT 80.9000 113.8000 81.3000 113.9000 ;
	    RECT 77.4000 113.3000 79.3000 113.6000 ;
	    RECT 77.4000 111.1000 77.8000 113.3000 ;
	    RECT 78.9000 113.2000 79.3000 113.3000 ;
	    RECT 83.8000 112.8000 84.1000 113.9000 ;
	    RECT 85.4000 113.8000 86.2000 113.9000 ;
	    RECT 87.8000 113.8000 88.2000 114.2000 ;
	    RECT 88.6000 113.8000 89.0000 114.2000 ;
	    RECT 89.8000 113.9000 95.3000 114.2000 ;
	    RECT 89.8000 113.8000 90.6000 113.9000 ;
	    RECT 82.9000 112.7000 83.3000 112.8000 ;
	    RECT 79.8000 112.1000 80.2000 112.5000 ;
	    RECT 81.9000 112.4000 83.3000 112.7000 ;
	    RECT 83.8000 112.4000 84.2000 112.8000 ;
	    RECT 81.9000 112.1000 82.2000 112.4000 ;
	    RECT 84.6000 112.1000 85.0000 112.5000 ;
	    RECT 79.5000 111.8000 80.2000 112.1000 ;
	    RECT 79.5000 111.1000 80.1000 111.8000 ;
	    RECT 81.8000 111.1000 82.2000 112.1000 ;
	    RECT 84.0000 111.8000 85.0000 112.1000 ;
	    RECT 84.0000 111.1000 84.4000 111.8000 ;
	    RECT 86.2000 111.1000 86.6000 113.5000 ;
	    RECT 87.8000 112.1000 88.1000 113.8000 ;
	    RECT 88.6000 112.4000 89.0000 113.2000 ;
	    RECT 87.8000 111.1000 88.2000 112.1000 ;
	    RECT 89.4000 111.1000 89.8000 113.5000 ;
	    RECT 91.9000 112.8000 92.2000 113.9000 ;
	    RECT 94.7000 113.8000 95.1000 113.9000 ;
	    RECT 98.2000 113.6000 98.6000 115.3000 ;
	    RECT 96.7000 113.3000 98.6000 113.6000 ;
	    RECT 96.7000 113.2000 97.1000 113.3000 ;
	    RECT 91.0000 112.1000 91.4000 112.5000 ;
	    RECT 91.8000 112.4000 92.2000 112.8000 ;
	    RECT 92.7000 112.7000 93.1000 112.8000 ;
	    RECT 92.7000 112.4000 94.1000 112.7000 ;
	    RECT 93.8000 112.1000 94.1000 112.4000 ;
	    RECT 95.8000 112.1000 96.2000 112.5000 ;
	    RECT 91.0000 111.8000 92.0000 112.1000 ;
	    RECT 91.6000 111.1000 92.0000 111.8000 ;
	    RECT 93.8000 111.1000 94.2000 112.1000 ;
	    RECT 95.8000 111.8000 96.5000 112.1000 ;
	    RECT 95.9000 111.1000 96.5000 111.8000 ;
	    RECT 98.2000 111.1000 98.6000 113.3000 ;
	    RECT 99.0000 111.1000 99.4000 119.9000 ;
	    RECT 101.4000 114.1000 101.8000 119.9000 ;
	    RECT 102.2000 119.6000 104.2000 119.9000 ;
	    RECT 102.2000 115.9000 102.6000 119.6000 ;
	    RECT 103.0000 115.9000 103.4000 119.3000 ;
	    RECT 103.8000 116.2000 104.2000 119.6000 ;
	    RECT 105.4000 116.2000 105.8000 119.9000 ;
	    RECT 103.8000 115.9000 105.8000 116.2000 ;
	    RECT 106.5000 116.3000 106.9000 119.9000 ;
	    RECT 106.5000 115.9000 107.4000 116.3000 ;
	    RECT 109.4000 116.1000 109.8000 116.2000 ;
	    RECT 110.2000 116.1000 110.6000 119.9000 ;
	    RECT 103.1000 115.6000 103.4000 115.9000 ;
	    RECT 102.2000 114.8000 102.6000 115.6000 ;
	    RECT 103.1000 115.3000 104.1000 115.6000 ;
	    RECT 103.8000 115.2000 104.1000 115.3000 ;
	    RECT 105.0000 115.2000 105.4000 115.4000 ;
	    RECT 103.8000 114.8000 104.2000 115.2000 ;
	    RECT 105.0000 115.1000 105.8000 115.2000 ;
	    RECT 106.2000 115.1000 106.6000 115.6000 ;
	    RECT 105.0000 114.9000 106.6000 115.1000 ;
	    RECT 105.4000 114.8000 106.6000 114.9000 ;
	    RECT 103.1000 114.4000 103.5000 114.8000 ;
	    RECT 103.1000 114.2000 103.4000 114.4000 ;
	    RECT 103.0000 114.1000 103.4000 114.2000 ;
	    RECT 101.4000 113.8000 103.4000 114.1000 ;
	    RECT 99.8000 112.4000 100.2000 113.2000 ;
	    RECT 100.6000 112.4000 101.0000 113.2000 ;
	    RECT 101.4000 111.1000 101.8000 113.8000 ;
	    RECT 103.8000 113.1000 104.1000 114.8000 ;
	    RECT 104.6000 113.8000 105.0000 114.6000 ;
	    RECT 107.0000 114.2000 107.3000 115.9000 ;
	    RECT 109.4000 115.8000 110.6000 116.1000 ;
	    RECT 107.0000 113.8000 107.4000 114.2000 ;
	    RECT 103.5000 112.2000 104.3000 113.1000 ;
	    RECT 103.0000 111.8000 104.3000 112.2000 ;
	    RECT 103.5000 111.1000 104.3000 111.8000 ;
	    RECT 107.0000 112.2000 107.3000 113.8000 ;
	    RECT 107.8000 112.4000 108.2000 113.2000 ;
	    RECT 107.0000 111.1000 107.4000 112.2000 ;
	    RECT 110.2000 111.1000 110.6000 115.8000 ;
	    RECT 111.0000 112.4000 111.4000 113.2000 ;
	    RECT 111.8000 111.1000 112.2000 119.9000 ;
	    RECT 113.4000 113.4000 113.8000 114.2000 ;
	    RECT 112.6000 112.4000 113.0000 113.2000 ;
	    RECT 114.2000 113.1000 114.6000 119.9000 ;
	    RECT 115.0000 116.1000 115.4000 116.6000 ;
	    RECT 115.8000 116.1000 116.2000 119.9000 ;
	    RECT 115.0000 115.8000 116.2000 116.1000 ;
	    RECT 114.2000 112.8000 115.1000 113.1000 ;
	    RECT 114.7000 112.2000 115.1000 112.8000 ;
	    RECT 114.2000 111.8000 115.1000 112.2000 ;
	    RECT 114.7000 111.1000 115.1000 111.8000 ;
	    RECT 115.8000 111.1000 116.2000 115.8000 ;
	    RECT 117.4000 113.4000 117.8000 114.2000 ;
	    RECT 116.6000 112.4000 117.0000 113.2000 ;
	    RECT 118.2000 113.1000 118.6000 119.9000 ;
	    RECT 119.0000 116.1000 119.4000 116.6000 ;
	    RECT 119.8000 116.1000 120.2000 119.9000 ;
	    RECT 119.0000 115.8000 120.2000 116.1000 ;
	    RECT 118.2000 112.8000 119.1000 113.1000 ;
	    RECT 118.7000 112.2000 119.1000 112.8000 ;
	    RECT 118.2000 111.8000 119.1000 112.2000 ;
	    RECT 118.7000 111.1000 119.1000 111.8000 ;
	    RECT 119.8000 111.1000 120.2000 115.8000 ;
	    RECT 121.4000 115.9000 121.8000 119.9000 ;
	    RECT 123.0000 116.2000 123.4000 119.9000 ;
	    RECT 125.1000 119.2000 125.5000 119.9000 ;
	    RECT 125.1000 118.8000 125.8000 119.2000 ;
	    RECT 125.1000 116.3000 125.5000 118.8000 ;
	    RECT 122.3000 115.9000 123.4000 116.2000 ;
	    RECT 124.6000 115.9000 125.5000 116.3000 ;
	    RECT 127.0000 116.1000 127.4000 119.9000 ;
	    RECT 128.6000 117.9000 129.0000 119.9000 ;
	    RECT 128.7000 117.8000 129.0000 117.9000 ;
	    RECT 130.2000 117.9000 130.6000 119.9000 ;
	    RECT 130.2000 117.8000 130.5000 117.9000 ;
	    RECT 128.7000 117.5000 130.5000 117.8000 ;
	    RECT 129.4000 116.4000 129.8000 117.2000 ;
	    RECT 130.2000 116.2000 130.5000 117.5000 ;
	    RECT 131.0000 117.1000 131.4000 119.9000 ;
	    RECT 131.8000 117.1000 132.2000 117.2000 ;
	    RECT 131.0000 116.8000 132.2000 117.1000 ;
	    RECT 133.0000 116.8000 133.4000 117.2000 ;
	    RECT 127.8000 116.1000 128.2000 116.2000 ;
	    RECT 121.4000 114.8000 121.7000 115.9000 ;
	    RECT 122.3000 115.6000 122.6000 115.9000 ;
	    RECT 122.0000 115.2000 122.6000 115.6000 ;
	    RECT 120.6000 112.4000 121.0000 113.2000 ;
	    RECT 121.4000 111.1000 121.8000 114.8000 ;
	    RECT 122.3000 113.7000 122.6000 115.2000 ;
	    RECT 124.7000 114.2000 125.0000 115.9000 ;
	    RECT 127.0000 115.8000 128.2000 116.1000 ;
	    RECT 125.4000 114.8000 125.8000 115.6000 ;
	    RECT 124.6000 113.8000 125.0000 114.2000 ;
	    RECT 122.3000 113.4000 123.4000 113.7000 ;
	    RECT 123.0000 111.1000 123.4000 113.4000 ;
	    RECT 123.8000 112.4000 124.2000 113.2000 ;
	    RECT 124.7000 112.1000 125.0000 113.8000 ;
	    RECT 126.2000 112.4000 126.6000 113.2000 ;
	    RECT 124.6000 111.1000 125.0000 112.1000 ;
	    RECT 127.0000 111.1000 127.4000 115.8000 ;
	    RECT 127.8000 115.4000 128.2000 115.8000 ;
	    RECT 130.2000 115.8000 130.6000 116.2000 ;
	    RECT 130.2000 115.2000 130.5000 115.8000 ;
	    RECT 128.6000 114.8000 129.4000 115.2000 ;
	    RECT 130.2000 114.8000 130.6000 115.2000 ;
	    RECT 130.2000 114.2000 130.5000 114.8000 ;
	    RECT 129.7000 114.1000 130.5000 114.2000 ;
	    RECT 129.6000 113.9000 130.5000 114.1000 ;
	    RECT 129.6000 111.1000 130.0000 113.9000 ;
	    RECT 131.0000 111.1000 131.4000 116.8000 ;
	    RECT 133.0000 116.2000 133.3000 116.8000 ;
	    RECT 133.7000 116.2000 134.1000 119.9000 ;
	    RECT 135.8000 116.2000 136.2000 119.9000 ;
	    RECT 137.4000 116.2000 137.8000 119.9000 ;
	    RECT 132.6000 115.9000 133.3000 116.2000 ;
	    RECT 132.6000 115.8000 133.0000 115.9000 ;
	    RECT 133.6000 115.8000 134.6000 116.2000 ;
	    RECT 135.8000 115.9000 137.8000 116.2000 ;
	    RECT 138.2000 115.9000 138.6000 119.9000 ;
	    RECT 139.4000 116.8000 139.8000 117.2000 ;
	    RECT 139.4000 116.2000 139.7000 116.8000 ;
	    RECT 140.1000 116.2000 140.5000 119.9000 ;
	    RECT 139.0000 115.9000 139.7000 116.2000 ;
	    RECT 140.0000 115.9000 140.5000 116.2000 ;
	    RECT 142.2000 115.9000 142.6000 119.9000 ;
	    RECT 143.0000 116.2000 143.4000 119.9000 ;
	    RECT 144.6000 116.2000 145.0000 119.9000 ;
	    RECT 143.0000 115.9000 145.0000 116.2000 ;
	    RECT 133.6000 114.2000 133.9000 115.8000 ;
	    RECT 136.2000 115.2000 136.6000 115.4000 ;
	    RECT 138.2000 115.2000 138.5000 115.9000 ;
	    RECT 139.0000 115.8000 139.4000 115.9000 ;
	    RECT 134.2000 114.4000 134.6000 115.2000 ;
	    RECT 135.8000 114.9000 136.6000 115.2000 ;
	    RECT 137.4000 114.9000 138.6000 115.2000 ;
	    RECT 135.8000 114.8000 136.2000 114.9000 ;
	    RECT 132.6000 113.8000 133.9000 114.2000 ;
	    RECT 135.0000 114.1000 135.4000 114.2000 ;
	    RECT 134.6000 113.8000 135.4000 114.1000 ;
	    RECT 136.6000 113.8000 137.0000 114.6000 ;
	    RECT 131.8000 112.4000 132.2000 113.2000 ;
	    RECT 132.7000 113.1000 133.0000 113.8000 ;
	    RECT 134.6000 113.6000 135.0000 113.8000 ;
	    RECT 133.5000 113.1000 135.3000 113.3000 ;
	    RECT 137.4000 113.1000 137.7000 114.9000 ;
	    RECT 138.2000 114.8000 138.6000 114.9000 ;
	    RECT 140.0000 114.2000 140.3000 115.9000 ;
	    RECT 142.3000 115.2000 142.6000 115.9000 ;
	    RECT 144.2000 115.2000 144.6000 115.4000 ;
	    RECT 140.6000 114.4000 141.0000 115.2000 ;
	    RECT 142.2000 114.9000 143.4000 115.2000 ;
	    RECT 144.2000 114.9000 145.0000 115.2000 ;
	    RECT 142.2000 114.8000 142.6000 114.9000 ;
	    RECT 139.0000 113.8000 140.3000 114.2000 ;
	    RECT 141.4000 114.1000 141.8000 114.2000 ;
	    RECT 141.0000 113.8000 141.8000 114.1000 ;
	    RECT 132.6000 111.1000 133.0000 113.1000 ;
	    RECT 133.4000 113.0000 135.4000 113.1000 ;
	    RECT 133.4000 111.1000 133.8000 113.0000 ;
	    RECT 135.0000 111.1000 135.4000 113.0000 ;
	    RECT 137.4000 111.1000 137.8000 113.1000 ;
	    RECT 138.2000 112.8000 138.6000 113.2000 ;
	    RECT 139.1000 113.1000 139.4000 113.8000 ;
	    RECT 141.0000 113.6000 141.4000 113.8000 ;
	    RECT 139.9000 113.1000 141.7000 113.3000 ;
	    RECT 138.1000 112.4000 138.5000 112.8000 ;
	    RECT 139.0000 111.1000 139.4000 113.1000 ;
	    RECT 139.8000 113.0000 141.8000 113.1000 ;
	    RECT 139.8000 111.1000 140.2000 113.0000 ;
	    RECT 141.4000 111.1000 141.8000 113.0000 ;
	    RECT 142.2000 112.8000 142.6000 113.2000 ;
	    RECT 143.1000 113.1000 143.4000 114.9000 ;
	    RECT 144.6000 114.8000 145.0000 114.9000 ;
	    RECT 143.8000 114.1000 144.2000 114.6000 ;
	    RECT 145.4000 114.1000 145.8000 119.9000 ;
	    RECT 147.0000 115.9000 147.4000 119.9000 ;
	    RECT 147.8000 116.2000 148.2000 119.9000 ;
	    RECT 149.4000 116.2000 149.8000 119.9000 ;
	    RECT 147.8000 115.9000 149.8000 116.2000 ;
	    RECT 147.1000 115.2000 147.4000 115.9000 ;
	    RECT 150.2000 115.8000 150.6000 116.2000 ;
	    RECT 149.0000 115.2000 149.4000 115.4000 ;
	    RECT 147.0000 114.9000 148.2000 115.2000 ;
	    RECT 149.0000 114.9000 149.8000 115.2000 ;
	    RECT 147.0000 114.8000 147.4000 114.9000 ;
	    RECT 143.8000 113.8000 145.8000 114.1000 ;
	    RECT 142.3000 112.4000 142.7000 112.8000 ;
	    RECT 143.0000 111.1000 143.4000 113.1000 ;
	    RECT 145.4000 111.1000 145.8000 113.8000 ;
	    RECT 147.0000 113.8000 147.4000 114.2000 ;
	    RECT 147.0000 113.2000 147.3000 113.8000 ;
	    RECT 146.2000 112.4000 146.6000 113.2000 ;
	    RECT 147.0000 112.8000 147.4000 113.2000 ;
	    RECT 147.9000 113.1000 148.2000 114.9000 ;
	    RECT 149.4000 114.8000 149.8000 114.9000 ;
	    RECT 150.2000 115.1000 150.5000 115.8000 ;
	    RECT 151.0000 115.1000 151.4000 119.9000 ;
	    RECT 151.8000 115.8000 152.2000 116.6000 ;
	    RECT 153.9000 116.2000 154.3000 119.9000 ;
	    RECT 154.6000 116.8000 155.0000 117.2000 ;
	    RECT 154.7000 116.2000 155.0000 116.8000 ;
	    RECT 156.6000 116.4000 157.0000 119.9000 ;
	    RECT 153.9000 115.9000 154.4000 116.2000 ;
	    RECT 154.7000 115.9000 155.4000 116.2000 ;
	    RECT 153.4000 115.1000 153.8000 115.2000 ;
	    RECT 150.2000 114.8000 153.8000 115.1000 ;
	    RECT 148.6000 113.8000 149.0000 114.6000 ;
	    RECT 150.2000 113.4000 150.6000 114.2000 ;
	    RECT 147.1000 112.4000 147.5000 112.8000 ;
	    RECT 147.8000 111.1000 148.2000 113.1000 ;
	    RECT 151.0000 113.1000 151.4000 114.8000 ;
	    RECT 153.4000 114.4000 153.8000 114.8000 ;
	    RECT 154.1000 114.2000 154.4000 115.9000 ;
	    RECT 155.0000 115.8000 155.4000 115.9000 ;
	    RECT 156.5000 115.9000 157.0000 116.4000 ;
	    RECT 158.2000 116.2000 158.6000 119.9000 ;
	    RECT 157.3000 115.9000 158.6000 116.2000 ;
	    RECT 155.0000 115.1000 155.3000 115.8000 ;
	    RECT 155.0000 114.8000 156.1000 115.1000 ;
	    RECT 152.6000 114.1000 153.0000 114.2000 ;
	    RECT 152.6000 113.8000 153.4000 114.1000 ;
	    RECT 154.1000 113.8000 155.4000 114.2000 ;
	    RECT 155.8000 114.1000 156.1000 114.8000 ;
	    RECT 156.5000 114.2000 156.8000 115.9000 ;
	    RECT 157.3000 114.9000 157.6000 115.9000 ;
	    RECT 160.6000 115.7000 161.0000 119.9000 ;
	    RECT 162.8000 118.2000 163.2000 119.9000 ;
	    RECT 162.2000 117.9000 163.2000 118.2000 ;
	    RECT 165.0000 117.9000 165.4000 119.9000 ;
	    RECT 167.1000 117.9000 167.7000 119.9000 ;
	    RECT 162.2000 117.5000 162.6000 117.9000 ;
	    RECT 165.0000 117.6000 165.3000 117.9000 ;
	    RECT 163.9000 117.3000 165.7000 117.6000 ;
	    RECT 167.0000 117.5000 167.4000 117.9000 ;
	    RECT 163.9000 117.2000 164.3000 117.3000 ;
	    RECT 165.3000 117.2000 165.7000 117.3000 ;
	    RECT 167.5000 117.0000 168.2000 117.2000 ;
	    RECT 167.1000 116.8000 168.2000 117.0000 ;
	    RECT 162.2000 116.5000 162.6000 116.6000 ;
	    RECT 164.5000 116.5000 164.9000 116.6000 ;
	    RECT 162.2000 116.2000 164.9000 116.5000 ;
	    RECT 165.2000 116.5000 166.3000 116.8000 ;
	    RECT 165.2000 115.9000 165.5000 116.5000 ;
	    RECT 165.9000 116.4000 166.3000 116.5000 ;
	    RECT 167.1000 116.6000 167.8000 116.8000 ;
	    RECT 167.1000 116.1000 167.4000 116.6000 ;
	    RECT 163.1000 115.7000 165.5000 115.9000 ;
	    RECT 160.6000 115.6000 165.5000 115.7000 ;
	    RECT 166.2000 115.8000 167.4000 116.1000 ;
	    RECT 160.6000 115.5000 163.5000 115.6000 ;
	    RECT 160.6000 115.4000 163.4000 115.5000 ;
	    RECT 163.8000 115.1000 164.2000 115.2000 ;
	    RECT 157.1000 114.5000 157.6000 114.9000 ;
	    RECT 161.7000 114.8000 164.2000 115.1000 ;
	    RECT 161.7000 114.7000 162.1000 114.8000 ;
	    RECT 163.0000 114.7000 163.4000 114.8000 ;
	    RECT 156.5000 114.1000 157.0000 114.2000 ;
	    RECT 155.8000 113.8000 157.0000 114.1000 ;
	    RECT 153.0000 113.6000 153.4000 113.8000 ;
	    RECT 152.7000 113.1000 154.5000 113.3000 ;
	    RECT 155.0000 113.1000 155.3000 113.8000 ;
	    RECT 156.5000 113.1000 156.8000 113.8000 ;
	    RECT 157.3000 113.7000 157.6000 114.5000 ;
	    RECT 162.5000 114.2000 162.9000 114.3000 ;
	    RECT 166.2000 114.2000 166.5000 115.8000 ;
	    RECT 169.4000 115.6000 169.8000 119.9000 ;
	    RECT 167.7000 115.3000 169.8000 115.6000 ;
	    RECT 167.7000 115.2000 168.1000 115.3000 ;
	    RECT 168.5000 114.9000 168.9000 115.0000 ;
	    RECT 167.0000 114.6000 168.9000 114.9000 ;
	    RECT 167.0000 114.5000 167.4000 114.6000 ;
	    RECT 161.0000 113.9000 166.5000 114.2000 ;
	    RECT 169.4000 114.1000 169.8000 115.3000 ;
	    RECT 170.2000 114.1000 170.6000 114.2000 ;
	    RECT 161.0000 113.8000 161.8000 113.9000 ;
	    RECT 157.3000 113.4000 158.6000 113.7000 ;
	    RECT 151.0000 112.8000 151.9000 113.1000 ;
	    RECT 151.5000 111.1000 151.9000 112.8000 ;
	    RECT 152.6000 113.0000 154.6000 113.1000 ;
	    RECT 152.6000 111.1000 153.0000 113.0000 ;
	    RECT 154.2000 111.1000 154.6000 113.0000 ;
	    RECT 155.0000 111.1000 155.4000 113.1000 ;
	    RECT 156.5000 112.8000 157.0000 113.1000 ;
	    RECT 156.6000 111.1000 157.0000 112.8000 ;
	    RECT 158.2000 111.1000 158.6000 113.4000 ;
	    RECT 160.6000 111.1000 161.0000 113.5000 ;
	    RECT 163.1000 112.8000 163.4000 113.9000 ;
	    RECT 164.6000 113.8000 165.0000 113.9000 ;
	    RECT 165.9000 113.8000 166.3000 113.9000 ;
	    RECT 169.4000 113.8000 170.6000 114.1000 ;
	    RECT 169.4000 113.6000 169.8000 113.8000 ;
	    RECT 167.9000 113.3000 169.8000 113.6000 ;
	    RECT 170.2000 113.4000 170.6000 113.8000 ;
	    RECT 171.0000 114.1000 171.4000 119.9000 ;
	    RECT 171.8000 116.9000 172.2000 119.9000 ;
	    RECT 171.9000 116.6000 172.2000 116.9000 ;
	    RECT 173.4000 119.6000 175.4000 119.9000 ;
	    RECT 173.4000 116.9000 173.8000 119.6000 ;
	    RECT 174.2000 116.9000 174.6000 119.3000 ;
	    RECT 175.0000 117.0000 175.4000 119.6000 ;
	    RECT 175.9000 119.6000 177.7000 119.9000 ;
	    RECT 175.9000 119.5000 176.2000 119.6000 ;
	    RECT 173.4000 116.6000 173.7000 116.9000 ;
	    RECT 171.9000 116.3000 173.7000 116.6000 ;
	    RECT 174.3000 116.7000 174.6000 116.9000 ;
	    RECT 175.8000 116.7000 176.2000 119.5000 ;
	    RECT 177.4000 119.5000 177.7000 119.6000 ;
	    RECT 174.3000 116.5000 176.2000 116.7000 ;
	    RECT 176.6000 116.5000 177.0000 119.3000 ;
	    RECT 177.4000 116.5000 177.8000 119.5000 ;
	    RECT 174.3000 116.4000 176.1000 116.5000 ;
	    RECT 176.6000 116.2000 176.9000 116.5000 ;
	    RECT 176.6000 116.1000 177.0000 116.2000 ;
	    RECT 175.3000 115.8000 177.0000 116.1000 ;
	    RECT 178.2000 115.9000 178.6000 119.9000 ;
	    RECT 179.8000 117.9000 180.2000 119.9000 ;
	    RECT 174.2000 114.8000 175.0000 115.2000 ;
	    RECT 173.4000 114.1000 174.2000 114.2000 ;
	    RECT 171.0000 113.8000 174.2000 114.1000 ;
	    RECT 167.9000 113.2000 168.3000 113.3000 ;
	    RECT 162.2000 112.1000 162.6000 112.5000 ;
	    RECT 163.0000 112.4000 163.4000 112.8000 ;
	    RECT 163.9000 112.7000 164.3000 112.8000 ;
	    RECT 163.9000 112.4000 165.3000 112.7000 ;
	    RECT 165.0000 112.1000 165.3000 112.4000 ;
	    RECT 167.0000 112.1000 167.4000 112.5000 ;
	    RECT 162.2000 111.8000 163.2000 112.1000 ;
	    RECT 162.8000 111.1000 163.2000 111.8000 ;
	    RECT 165.0000 111.1000 165.4000 112.1000 ;
	    RECT 167.0000 111.8000 167.7000 112.1000 ;
	    RECT 167.1000 111.1000 167.7000 111.8000 ;
	    RECT 169.4000 111.1000 169.8000 113.3000 ;
	    RECT 171.0000 111.1000 171.4000 113.8000 ;
	    RECT 172.6000 112.8000 173.8000 113.2000 ;
	    RECT 175.3000 112.5000 175.6000 115.8000 ;
	    RECT 178.2000 115.2000 178.5000 115.9000 ;
	    RECT 179.8000 115.8000 180.1000 117.9000 ;
	    RECT 178.9000 115.5000 180.1000 115.8000 ;
	    RECT 181.4000 115.7000 181.8000 119.9000 ;
	    RECT 183.6000 118.2000 184.0000 119.9000 ;
	    RECT 183.0000 117.9000 184.0000 118.2000 ;
	    RECT 185.8000 117.9000 186.2000 119.9000 ;
	    RECT 187.9000 117.9000 188.5000 119.9000 ;
	    RECT 183.0000 117.5000 183.4000 117.9000 ;
	    RECT 185.8000 117.6000 186.1000 117.9000 ;
	    RECT 184.7000 117.3000 186.5000 117.6000 ;
	    RECT 187.8000 117.5000 188.2000 117.9000 ;
	    RECT 184.7000 117.2000 185.1000 117.3000 ;
	    RECT 186.1000 117.2000 186.5000 117.3000 ;
	    RECT 183.0000 116.5000 183.4000 116.6000 ;
	    RECT 185.3000 116.5000 185.7000 116.6000 ;
	    RECT 183.0000 116.2000 185.7000 116.5000 ;
	    RECT 186.0000 116.5000 187.1000 116.8000 ;
	    RECT 186.0000 115.9000 186.3000 116.5000 ;
	    RECT 186.7000 116.4000 187.1000 116.5000 ;
	    RECT 187.9000 116.6000 188.6000 117.0000 ;
	    RECT 187.9000 116.1000 188.2000 116.6000 ;
	    RECT 183.9000 115.7000 186.3000 115.9000 ;
	    RECT 181.4000 115.6000 186.3000 115.7000 ;
	    RECT 187.0000 115.8000 188.2000 116.1000 ;
	    RECT 181.4000 115.5000 184.3000 115.6000 ;
	    RECT 178.2000 114.8000 178.6000 115.2000 ;
	    RECT 178.2000 113.1000 178.5000 114.8000 ;
	    RECT 178.9000 113.8000 179.2000 115.5000 ;
	    RECT 181.4000 115.4000 184.2000 115.5000 ;
	    RECT 179.8000 114.8000 180.2000 115.2000 ;
	    RECT 184.6000 115.1000 185.0000 115.2000 ;
	    RECT 182.5000 114.8000 185.0000 115.1000 ;
	    RECT 179.8000 114.4000 180.1000 114.8000 ;
	    RECT 182.5000 114.7000 182.9000 114.8000 ;
	    RECT 183.8000 114.7000 184.2000 114.8000 ;
	    RECT 179.6000 114.1000 180.1000 114.4000 ;
	    RECT 179.6000 114.0000 180.0000 114.1000 ;
	    RECT 180.6000 113.8000 181.0000 114.6000 ;
	    RECT 183.3000 114.2000 183.7000 114.3000 ;
	    RECT 187.0000 114.2000 187.3000 115.8000 ;
	    RECT 190.2000 115.6000 190.6000 119.9000 ;
	    RECT 188.5000 115.3000 190.6000 115.6000 ;
	    RECT 191.0000 115.7000 191.4000 119.9000 ;
	    RECT 193.2000 118.2000 193.6000 119.9000 ;
	    RECT 192.6000 117.9000 193.6000 118.2000 ;
	    RECT 195.4000 117.9000 195.8000 119.9000 ;
	    RECT 197.5000 117.9000 198.1000 119.9000 ;
	    RECT 192.6000 117.5000 193.0000 117.9000 ;
	    RECT 195.4000 117.6000 195.7000 117.9000 ;
	    RECT 194.3000 117.3000 196.1000 117.6000 ;
	    RECT 197.4000 117.5000 197.8000 117.9000 ;
	    RECT 194.3000 117.2000 194.7000 117.3000 ;
	    RECT 195.7000 117.2000 196.1000 117.3000 ;
	    RECT 197.9000 117.0000 198.6000 117.2000 ;
	    RECT 197.5000 116.8000 198.6000 117.0000 ;
	    RECT 192.6000 116.5000 193.0000 116.6000 ;
	    RECT 194.9000 116.5000 195.3000 116.6000 ;
	    RECT 192.6000 116.2000 195.3000 116.5000 ;
	    RECT 195.6000 116.5000 196.7000 116.8000 ;
	    RECT 195.6000 115.9000 195.9000 116.5000 ;
	    RECT 196.3000 116.4000 196.7000 116.5000 ;
	    RECT 197.5000 116.6000 198.2000 116.8000 ;
	    RECT 197.5000 116.1000 197.8000 116.6000 ;
	    RECT 193.5000 115.7000 195.9000 115.9000 ;
	    RECT 191.0000 115.6000 195.9000 115.7000 ;
	    RECT 196.6000 115.8000 197.8000 116.1000 ;
	    RECT 191.0000 115.5000 193.9000 115.6000 ;
	    RECT 191.0000 115.4000 193.8000 115.5000 ;
	    RECT 188.5000 115.2000 188.9000 115.3000 ;
	    RECT 189.3000 114.9000 189.7000 115.0000 ;
	    RECT 187.8000 114.6000 189.7000 114.9000 ;
	    RECT 187.8000 114.5000 188.2000 114.6000 ;
	    RECT 181.8000 113.9000 187.3000 114.2000 ;
	    RECT 181.8000 113.8000 182.6000 113.9000 ;
	    RECT 178.8000 113.7000 179.2000 113.8000 ;
	    RECT 178.8000 113.5000 180.3000 113.7000 ;
	    RECT 178.8000 113.4000 180.9000 113.5000 ;
	    RECT 180.0000 113.2000 180.9000 113.4000 ;
	    RECT 180.6000 113.1000 180.9000 113.2000 ;
	    RECT 178.2000 112.6000 178.9000 113.1000 ;
	    RECT 173.6000 112.2000 175.6000 112.5000 ;
	    RECT 173.4000 111.8000 173.9000 112.2000 ;
	    RECT 175.0000 112.1000 175.6000 112.2000 ;
	    RECT 177.4000 112.1000 177.8000 112.2000 ;
	    RECT 178.5000 112.1000 178.9000 112.6000 ;
	    RECT 173.4000 111.1000 173.8000 111.8000 ;
	    RECT 175.0000 111.1000 175.4000 112.1000 ;
	    RECT 177.4000 111.8000 178.9000 112.1000 ;
	    RECT 178.5000 111.1000 178.9000 111.8000 ;
	    RECT 180.6000 111.1000 181.0000 113.1000 ;
	    RECT 181.4000 111.1000 181.8000 113.5000 ;
	    RECT 183.9000 112.8000 184.2000 113.9000 ;
	    RECT 186.7000 113.8000 187.1000 113.9000 ;
	    RECT 190.2000 113.6000 190.6000 115.3000 ;
	    RECT 194.2000 115.1000 194.6000 115.2000 ;
	    RECT 192.1000 114.8000 194.6000 115.1000 ;
	    RECT 192.1000 114.7000 192.5000 114.8000 ;
	    RECT 193.4000 114.7000 193.8000 114.8000 ;
	    RECT 192.9000 114.2000 193.3000 114.3000 ;
	    RECT 196.6000 114.2000 196.9000 115.8000 ;
	    RECT 199.8000 115.6000 200.2000 119.9000 ;
	    RECT 198.1000 115.3000 200.2000 115.6000 ;
	    RECT 198.1000 115.2000 198.5000 115.3000 ;
	    RECT 198.9000 114.9000 199.3000 115.0000 ;
	    RECT 197.4000 114.6000 199.3000 114.9000 ;
	    RECT 197.4000 114.5000 197.8000 114.6000 ;
	    RECT 191.4000 113.9000 197.0000 114.2000 ;
	    RECT 191.4000 113.8000 192.2000 113.9000 ;
	    RECT 188.7000 113.3000 190.6000 113.6000 ;
	    RECT 188.7000 113.2000 189.1000 113.3000 ;
	    RECT 183.0000 112.1000 183.4000 112.5000 ;
	    RECT 183.8000 112.4000 184.2000 112.8000 ;
	    RECT 184.7000 112.7000 185.1000 112.8000 ;
	    RECT 184.7000 112.4000 186.1000 112.7000 ;
	    RECT 185.8000 112.1000 186.1000 112.4000 ;
	    RECT 187.8000 112.1000 188.2000 112.5000 ;
	    RECT 183.0000 111.8000 184.0000 112.1000 ;
	    RECT 183.6000 111.1000 184.0000 111.8000 ;
	    RECT 185.8000 111.1000 186.2000 112.1000 ;
	    RECT 187.8000 111.8000 188.5000 112.1000 ;
	    RECT 187.9000 111.1000 188.5000 111.8000 ;
	    RECT 190.2000 111.1000 190.6000 113.3000 ;
	    RECT 191.0000 111.1000 191.4000 113.5000 ;
	    RECT 193.5000 112.8000 193.8000 113.9000 ;
	    RECT 196.3000 113.8000 197.0000 113.9000 ;
	    RECT 199.8000 113.6000 200.2000 115.3000 ;
	    RECT 201.4000 115.6000 201.8000 119.9000 ;
	    RECT 203.0000 115.6000 203.4000 119.9000 ;
	    RECT 204.9000 116.3000 205.3000 119.9000 ;
	    RECT 204.9000 115.9000 205.8000 116.3000 ;
	    RECT 201.4000 115.2000 203.4000 115.6000 ;
	    RECT 198.3000 113.3000 200.2000 113.6000 ;
	    RECT 200.6000 113.4000 201.0000 114.2000 ;
	    RECT 203.0000 113.8000 203.4000 115.2000 ;
	    RECT 204.6000 114.8000 205.0000 115.6000 ;
	    RECT 205.4000 115.1000 205.7000 115.9000 ;
	    RECT 207.0000 115.8000 207.4000 116.6000 ;
	    RECT 207.0000 115.1000 207.3000 115.8000 ;
	    RECT 205.4000 114.8000 207.3000 115.1000 ;
	    RECT 201.4000 113.4000 203.4000 113.8000 ;
	    RECT 198.3000 113.2000 198.7000 113.3000 ;
	    RECT 192.6000 112.1000 193.0000 112.5000 ;
	    RECT 193.4000 112.4000 193.8000 112.8000 ;
	    RECT 194.3000 112.7000 194.7000 112.8000 ;
	    RECT 194.3000 112.4000 195.7000 112.7000 ;
	    RECT 195.4000 112.1000 195.7000 112.4000 ;
	    RECT 197.4000 112.1000 197.8000 112.5000 ;
	    RECT 192.6000 111.8000 193.6000 112.1000 ;
	    RECT 193.2000 111.1000 193.6000 111.8000 ;
	    RECT 195.4000 111.1000 195.8000 112.1000 ;
	    RECT 197.4000 111.8000 198.1000 112.1000 ;
	    RECT 197.5000 111.1000 198.1000 111.8000 ;
	    RECT 199.8000 111.1000 200.2000 113.3000 ;
	    RECT 201.4000 111.1000 201.8000 113.4000 ;
	    RECT 203.0000 111.1000 203.4000 113.4000 ;
	    RECT 205.4000 114.2000 205.7000 114.8000 ;
	    RECT 205.4000 113.8000 205.8000 114.2000 ;
	    RECT 205.4000 112.1000 205.7000 113.8000 ;
	    RECT 206.2000 112.4000 206.6000 113.2000 ;
	    RECT 207.8000 113.1000 208.2000 119.9000 ;
	    RECT 208.6000 114.1000 209.0000 114.2000 ;
	    RECT 209.4000 114.1000 209.8000 114.2000 ;
	    RECT 208.6000 113.8000 209.8000 114.1000 ;
	    RECT 210.2000 114.1000 210.6000 119.9000 ;
	    RECT 213.9000 119.2000 214.3000 119.9000 ;
	    RECT 213.4000 118.8000 214.3000 119.2000 ;
	    RECT 213.9000 116.2000 214.3000 118.8000 ;
	    RECT 214.6000 116.8000 215.0000 117.2000 ;
	    RECT 214.7000 116.2000 215.0000 116.8000 ;
	    RECT 213.9000 115.9000 214.4000 116.2000 ;
	    RECT 214.7000 115.9000 215.4000 116.2000 ;
	    RECT 212.6000 115.1000 213.0000 115.2000 ;
	    RECT 213.4000 115.1000 213.8000 115.2000 ;
	    RECT 212.6000 114.8000 213.8000 115.1000 ;
	    RECT 213.4000 114.4000 213.8000 114.8000 ;
	    RECT 214.1000 114.2000 214.4000 115.9000 ;
	    RECT 215.0000 115.8000 215.4000 115.9000 ;
	    RECT 216.6000 115.1000 217.0000 119.9000 ;
	    RECT 217.7000 116.3000 218.1000 119.9000 ;
	    RECT 221.1000 116.3000 221.5000 119.9000 ;
	    RECT 223.3000 119.2000 223.7000 119.9000 ;
	    RECT 223.3000 118.8000 224.2000 119.2000 ;
	    RECT 217.7000 115.9000 218.6000 116.3000 ;
	    RECT 220.6000 115.9000 221.5000 116.3000 ;
	    RECT 222.6000 116.8000 223.0000 117.2000 ;
	    RECT 222.6000 116.2000 222.9000 116.8000 ;
	    RECT 223.3000 116.2000 223.7000 118.8000 ;
	    RECT 226.2000 117.9000 226.6000 119.9000 ;
	    RECT 222.2000 115.9000 222.9000 116.2000 ;
	    RECT 223.2000 115.9000 223.7000 116.2000 ;
	    RECT 218.2000 115.8000 218.6000 115.9000 ;
	    RECT 217.4000 115.1000 217.8000 115.6000 ;
	    RECT 216.6000 114.8000 217.8000 115.1000 ;
	    RECT 212.6000 114.1000 213.0000 114.2000 ;
	    RECT 210.2000 113.8000 213.4000 114.1000 ;
	    RECT 214.1000 113.8000 215.4000 114.2000 ;
	    RECT 208.6000 113.4000 209.0000 113.8000 ;
	    RECT 207.3000 112.8000 208.2000 113.1000 ;
	    RECT 207.3000 112.2000 207.7000 112.8000 ;
	    RECT 209.4000 112.4000 209.8000 113.2000 ;
	    RECT 205.4000 111.1000 205.8000 112.1000 ;
	    RECT 207.0000 111.8000 207.7000 112.2000 ;
	    RECT 207.3000 111.1000 207.7000 111.8000 ;
	    RECT 210.2000 111.1000 210.6000 113.8000 ;
	    RECT 213.0000 113.6000 213.4000 113.8000 ;
	    RECT 212.7000 113.1000 214.5000 113.3000 ;
	    RECT 215.0000 113.1000 215.3000 113.8000 ;
	    RECT 212.6000 113.0000 214.6000 113.1000 ;
	    RECT 212.6000 111.1000 213.0000 113.0000 ;
	    RECT 214.2000 111.1000 214.6000 113.0000 ;
	    RECT 215.0000 111.1000 215.4000 113.1000 ;
	    RECT 215.8000 112.4000 216.2000 113.2000 ;
	    RECT 216.6000 111.1000 217.0000 114.8000 ;
	    RECT 218.2000 114.2000 218.5000 115.8000 ;
	    RECT 220.7000 114.2000 221.0000 115.9000 ;
	    RECT 222.2000 115.8000 222.6000 115.9000 ;
	    RECT 221.4000 114.8000 221.8000 115.6000 ;
	    RECT 223.2000 114.2000 223.5000 115.9000 ;
	    RECT 226.3000 115.8000 226.6000 117.9000 ;
	    RECT 227.8000 115.9000 228.2000 119.9000 ;
	    RECT 226.3000 115.5000 227.5000 115.8000 ;
	    RECT 223.8000 114.4000 224.2000 115.2000 ;
	    RECT 226.2000 114.8000 226.6000 115.2000 ;
	    RECT 218.2000 113.8000 218.6000 114.2000 ;
	    RECT 220.6000 113.8000 221.0000 114.2000 ;
	    RECT 222.2000 113.8000 223.5000 114.2000 ;
	    RECT 224.6000 114.1000 225.0000 114.2000 ;
	    RECT 224.2000 113.8000 225.0000 114.1000 ;
	    RECT 225.4000 113.8000 225.8000 114.6000 ;
	    RECT 226.3000 114.4000 226.6000 114.8000 ;
	    RECT 226.2000 114.0000 226.8000 114.4000 ;
	    RECT 227.2000 113.8000 227.5000 115.5000 ;
	    RECT 227.9000 115.2000 228.2000 115.9000 ;
	    RECT 227.8000 114.8000 228.2000 115.2000 ;
	    RECT 218.2000 112.1000 218.5000 113.8000 ;
	    RECT 219.0000 113.1000 219.4000 113.2000 ;
	    RECT 219.8000 113.1000 220.2000 113.2000 ;
	    RECT 220.7000 113.1000 221.0000 113.8000 ;
	    RECT 221.4000 113.1000 221.8000 113.2000 ;
	    RECT 222.3000 113.1000 222.6000 113.8000 ;
	    RECT 224.2000 113.6000 224.6000 113.8000 ;
	    RECT 227.2000 113.7000 227.6000 113.8000 ;
	    RECT 226.1000 113.5000 227.6000 113.7000 ;
	    RECT 225.5000 113.4000 227.6000 113.5000 ;
	    RECT 223.1000 113.1000 224.9000 113.3000 ;
	    RECT 225.5000 113.2000 226.4000 113.4000 ;
	    RECT 225.5000 113.1000 225.8000 113.2000 ;
	    RECT 227.9000 113.1000 228.2000 114.8000 ;
	    RECT 229.4000 115.1000 229.8000 119.9000 ;
	    RECT 230.2000 115.8000 230.6000 116.6000 ;
	    RECT 231.3000 116.3000 231.7000 119.9000 ;
	    RECT 234.7000 116.3000 235.1000 119.9000 ;
	    RECT 231.3000 115.9000 232.2000 116.3000 ;
	    RECT 234.2000 115.9000 235.1000 116.3000 ;
	    RECT 231.0000 115.1000 231.4000 115.6000 ;
	    RECT 229.4000 114.8000 231.4000 115.1000 ;
	    RECT 228.6000 113.4000 229.0000 114.2000 ;
	    RECT 219.0000 112.8000 220.2000 113.1000 ;
	    RECT 220.6000 112.8000 221.8000 113.1000 ;
	    RECT 219.0000 112.4000 219.4000 112.8000 ;
	    RECT 219.8000 112.4000 220.2000 112.8000 ;
	    RECT 220.7000 112.1000 221.0000 112.8000 ;
	    RECT 218.2000 111.1000 218.6000 112.1000 ;
	    RECT 220.6000 111.1000 221.0000 112.1000 ;
	    RECT 222.2000 111.1000 222.6000 113.1000 ;
	    RECT 223.0000 113.0000 225.0000 113.1000 ;
	    RECT 223.0000 111.1000 223.4000 113.0000 ;
	    RECT 224.6000 111.1000 225.0000 113.0000 ;
	    RECT 225.4000 111.1000 225.8000 113.1000 ;
	    RECT 227.5000 112.6000 228.2000 113.1000 ;
	    RECT 229.4000 113.1000 229.8000 114.8000 ;
	    RECT 231.8000 114.2000 232.1000 115.9000 ;
	    RECT 234.3000 114.2000 234.6000 115.9000 ;
	    RECT 235.0000 114.8000 235.4000 115.6000 ;
	    RECT 231.8000 113.8000 232.2000 114.2000 ;
	    RECT 234.2000 113.8000 234.6000 114.2000 ;
	    RECT 229.4000 112.8000 230.3000 113.1000 ;
	    RECT 227.5000 112.2000 227.9000 112.6000 ;
	    RECT 227.5000 111.8000 228.2000 112.2000 ;
	    RECT 227.5000 111.1000 227.9000 111.8000 ;
	    RECT 229.9000 111.1000 230.3000 112.8000 ;
	    RECT 231.8000 112.2000 232.1000 113.8000 ;
	    RECT 232.6000 113.1000 233.0000 113.2000 ;
	    RECT 233.4000 113.1000 233.8000 113.2000 ;
	    RECT 232.6000 112.8000 233.8000 113.1000 ;
	    RECT 232.6000 112.4000 233.0000 112.8000 ;
	    RECT 233.4000 112.4000 233.8000 112.8000 ;
	    RECT 234.3000 112.2000 234.6000 113.8000 ;
	    RECT 235.8000 113.4000 236.2000 114.2000 ;
	    RECT 236.6000 113.1000 237.0000 119.9000 ;
	    RECT 239.0000 117.9000 239.4000 119.9000 ;
	    RECT 237.4000 115.8000 237.8000 116.6000 ;
	    RECT 239.1000 115.8000 239.4000 117.9000 ;
	    RECT 240.6000 115.9000 241.0000 119.9000 ;
	    RECT 239.1000 115.5000 240.3000 115.8000 ;
	    RECT 239.0000 114.8000 239.4000 115.2000 ;
	    RECT 237.4000 114.1000 237.8000 114.2000 ;
	    RECT 238.2000 114.1000 238.6000 114.6000 ;
	    RECT 239.1000 114.4000 239.4000 114.8000 ;
	    RECT 239.1000 114.1000 239.6000 114.4000 ;
	    RECT 237.4000 113.8000 238.6000 114.1000 ;
	    RECT 239.2000 114.0000 239.6000 114.1000 ;
	    RECT 240.0000 113.8000 240.3000 115.5000 ;
	    RECT 240.7000 115.2000 241.0000 115.9000 ;
	    RECT 240.6000 114.8000 241.0000 115.2000 ;
	    RECT 240.0000 113.7000 240.4000 113.8000 ;
	    RECT 238.9000 113.5000 240.4000 113.7000 ;
	    RECT 238.3000 113.4000 240.4000 113.5000 ;
	    RECT 238.3000 113.2000 239.2000 113.4000 ;
	    RECT 238.3000 113.1000 238.6000 113.2000 ;
	    RECT 240.7000 113.1000 241.0000 114.8000 ;
	    RECT 241.4000 113.4000 241.8000 114.2000 ;
	    RECT 236.6000 112.8000 237.5000 113.1000 ;
	    RECT 237.1000 112.2000 237.5000 112.8000 ;
	    RECT 231.8000 111.1000 232.2000 112.2000 ;
	    RECT 234.2000 111.1000 234.6000 112.2000 ;
	    RECT 236.6000 111.8000 237.5000 112.2000 ;
	    RECT 237.1000 111.1000 237.5000 111.8000 ;
	    RECT 238.2000 111.1000 238.6000 113.1000 ;
	    RECT 240.3000 112.6000 241.0000 113.1000 ;
	    RECT 242.2000 113.1000 242.6000 119.9000 ;
	    RECT 243.0000 116.1000 243.4000 116.6000 ;
	    RECT 243.8000 116.1000 244.2000 116.6000 ;
	    RECT 243.0000 115.8000 244.2000 116.1000 ;
	    RECT 244.6000 113.1000 245.0000 119.9000 ;
	    RECT 247.0000 115.1000 247.4000 119.9000 ;
	    RECT 247.8000 116.1000 248.2000 116.6000 ;
	    RECT 248.6000 116.1000 249.0000 116.6000 ;
	    RECT 247.8000 115.8000 249.0000 116.1000 ;
	    RECT 247.8000 115.1000 248.2000 115.2000 ;
	    RECT 247.0000 114.8000 248.2000 115.1000 ;
	    RECT 245.4000 113.4000 245.8000 114.2000 ;
	    RECT 246.2000 113.4000 246.6000 114.2000 ;
	    RECT 242.2000 112.8000 243.1000 113.1000 ;
	    RECT 240.3000 112.2000 240.7000 112.6000 ;
	    RECT 242.7000 112.2000 243.1000 112.8000 ;
	    RECT 244.1000 112.8000 245.0000 113.1000 ;
	    RECT 247.0000 113.1000 247.4000 114.8000 ;
	    RECT 249.4000 113.1000 249.8000 119.9000 ;
	    RECT 251.3000 116.3000 251.7000 119.9000 ;
	    RECT 253.7000 116.3000 254.1000 119.9000 ;
	    RECT 256.1000 116.3000 256.5000 119.9000 ;
	    RECT 258.5000 116.3000 258.9000 119.9000 ;
	    RECT 251.3000 115.9000 252.2000 116.3000 ;
	    RECT 253.7000 115.9000 254.6000 116.3000 ;
	    RECT 256.1000 115.9000 257.0000 116.3000 ;
	    RECT 258.5000 115.9000 259.4000 116.3000 ;
	    RECT 261.9000 116.2000 262.3000 119.9000 ;
	    RECT 265.1000 119.2000 265.5000 119.9000 ;
	    RECT 264.6000 118.8000 265.5000 119.2000 ;
	    RECT 262.6000 116.8000 263.0000 117.2000 ;
	    RECT 262.7000 116.2000 263.0000 116.8000 ;
	    RECT 265.1000 116.2000 265.5000 118.8000 ;
	    RECT 265.8000 116.8000 266.2000 117.2000 ;
	    RECT 265.9000 116.2000 266.2000 116.8000 ;
	    RECT 261.9000 115.9000 262.4000 116.2000 ;
	    RECT 262.7000 115.9000 263.4000 116.2000 ;
	    RECT 265.1000 115.9000 265.6000 116.2000 ;
	    RECT 265.9000 115.9000 266.6000 116.2000 ;
	    RECT 251.0000 114.8000 251.4000 115.6000 ;
	    RECT 251.8000 114.2000 252.1000 115.9000 ;
	    RECT 253.4000 114.8000 253.8000 115.6000 ;
	    RECT 254.2000 115.2000 254.5000 115.9000 ;
	    RECT 254.2000 114.8000 254.6000 115.2000 ;
	    RECT 255.8000 114.8000 256.2000 115.6000 ;
	    RECT 254.2000 114.2000 254.5000 114.8000 ;
	    RECT 256.6000 114.2000 256.9000 115.9000 ;
	    RECT 258.2000 114.8000 258.6000 115.6000 ;
	    RECT 259.0000 115.1000 259.3000 115.9000 ;
	    RECT 261.4000 115.1000 261.8000 115.2000 ;
	    RECT 259.0000 114.8000 261.8000 115.1000 ;
	    RECT 259.0000 114.2000 259.3000 114.8000 ;
	    RECT 261.4000 114.4000 261.8000 114.8000 ;
	    RECT 262.1000 114.2000 262.4000 115.9000 ;
	    RECT 263.0000 115.8000 263.4000 115.9000 ;
	    RECT 263.0000 115.1000 263.4000 115.2000 ;
	    RECT 264.6000 115.1000 265.0000 115.2000 ;
	    RECT 263.0000 114.8000 265.0000 115.1000 ;
	    RECT 264.6000 114.4000 265.0000 114.8000 ;
	    RECT 265.3000 114.2000 265.6000 115.9000 ;
	    RECT 266.2000 115.8000 266.6000 115.9000 ;
	    RECT 267.0000 115.8000 267.4000 116.6000 ;
	    RECT 250.2000 113.4000 250.6000 114.2000 ;
	    RECT 251.8000 113.8000 252.2000 114.2000 ;
	    RECT 254.2000 113.8000 254.6000 114.2000 ;
	    RECT 256.6000 114.1000 257.0000 114.2000 ;
	    RECT 257.4000 114.1000 257.8000 114.2000 ;
	    RECT 256.6000 113.8000 257.8000 114.1000 ;
	    RECT 259.0000 113.8000 259.4000 114.2000 ;
	    RECT 260.6000 114.1000 261.0000 114.2000 ;
	    RECT 260.6000 113.8000 261.4000 114.1000 ;
	    RECT 262.1000 113.8000 263.4000 114.2000 ;
	    RECT 263.8000 114.1000 264.2000 114.2000 ;
	    RECT 263.8000 113.8000 264.6000 114.1000 ;
	    RECT 265.3000 113.8000 266.6000 114.2000 ;
	    RECT 247.0000 112.8000 247.9000 113.1000 ;
	    RECT 244.1000 112.2000 244.5000 112.8000 ;
	    RECT 240.3000 111.8000 241.0000 112.2000 ;
	    RECT 242.7000 111.8000 243.4000 112.2000 ;
	    RECT 243.8000 111.8000 244.5000 112.2000 ;
	    RECT 240.3000 111.1000 240.7000 111.8000 ;
	    RECT 242.7000 111.1000 243.1000 111.8000 ;
	    RECT 244.1000 111.1000 244.5000 111.8000 ;
	    RECT 247.5000 111.1000 247.9000 112.8000 ;
	    RECT 248.9000 112.8000 249.8000 113.1000 ;
	    RECT 248.9000 112.2000 249.3000 112.8000 ;
	    RECT 251.8000 112.2000 252.1000 113.8000 ;
	    RECT 252.6000 112.4000 253.0000 113.2000 ;
	    RECT 248.9000 111.8000 249.8000 112.2000 ;
	    RECT 248.9000 111.1000 249.3000 111.8000 ;
	    RECT 251.8000 111.1000 252.2000 112.2000 ;
	    RECT 254.2000 112.1000 254.5000 113.8000 ;
	    RECT 255.0000 112.4000 255.4000 113.2000 ;
	    RECT 256.6000 112.1000 256.9000 113.8000 ;
	    RECT 257.4000 112.4000 257.8000 113.2000 ;
	    RECT 259.0000 112.1000 259.3000 113.8000 ;
	    RECT 261.0000 113.6000 261.4000 113.8000 ;
	    RECT 260.7000 113.1000 262.5000 113.3000 ;
	    RECT 263.0000 113.1000 263.3000 113.8000 ;
	    RECT 264.2000 113.6000 264.6000 113.8000 ;
	    RECT 263.9000 113.1000 265.7000 113.3000 ;
	    RECT 266.2000 113.1000 266.5000 113.8000 ;
	    RECT 267.8000 113.1000 268.2000 119.9000 ;
	    RECT 260.6000 113.0000 262.6000 113.1000 ;
	    RECT 254.2000 111.1000 254.6000 112.1000 ;
	    RECT 256.6000 111.1000 257.0000 112.1000 ;
	    RECT 259.0000 111.1000 259.4000 112.1000 ;
	    RECT 260.6000 111.1000 261.0000 113.0000 ;
	    RECT 262.2000 111.1000 262.6000 113.0000 ;
	    RECT 263.0000 111.1000 263.4000 113.1000 ;
	    RECT 263.8000 113.0000 265.8000 113.1000 ;
	    RECT 263.8000 111.1000 264.2000 113.0000 ;
	    RECT 265.4000 111.1000 265.8000 113.0000 ;
	    RECT 266.2000 111.1000 266.6000 113.1000 ;
	    RECT 267.3000 112.8000 268.2000 113.1000 ;
	    RECT 267.3000 112.2000 267.7000 112.8000 ;
	    RECT 267.3000 111.8000 268.2000 112.2000 ;
	    RECT 267.3000 111.1000 267.7000 111.8000 ;
	    RECT 0.6000 108.0000 1.0000 109.9000 ;
	    RECT 2.2000 108.0000 2.6000 109.9000 ;
	    RECT 0.6000 107.9000 2.6000 108.0000 ;
	    RECT 3.0000 107.9000 3.4000 109.9000 ;
	    RECT 5.1000 108.2000 5.5000 109.9000 ;
	    RECT 4.6000 107.9000 5.5000 108.2000 ;
	    RECT 7.0000 108.9000 7.4000 109.9000 ;
	    RECT 0.7000 107.7000 2.5000 107.9000 ;
	    RECT 1.0000 107.2000 1.4000 107.4000 ;
	    RECT 3.0000 107.2000 3.3000 107.9000 ;
	    RECT 0.6000 106.9000 1.4000 107.2000 ;
	    RECT 0.6000 106.8000 1.0000 106.9000 ;
	    RECT 2.1000 106.8000 3.4000 107.2000 ;
	    RECT 3.8000 106.8000 4.2000 107.6000 ;
	    RECT 4.6000 107.1000 5.0000 107.9000 ;
	    RECT 7.0000 107.2000 7.3000 108.9000 ;
	    RECT 7.8000 107.8000 8.2000 108.6000 ;
	    RECT 10.2000 107.9000 10.6000 109.9000 ;
	    RECT 13.1000 109.2000 13.5000 109.9000 ;
	    RECT 13.1000 108.8000 13.8000 109.2000 ;
	    RECT 10.9000 108.2000 11.3000 108.6000 ;
	    RECT 13.1000 108.2000 13.5000 108.8000 ;
	    RECT 5.4000 107.1000 5.8000 107.2000 ;
	    RECT 4.6000 106.8000 5.8000 107.1000 ;
	    RECT 7.0000 106.8000 7.4000 107.2000 ;
	    RECT 1.4000 105.8000 1.8000 106.6000 ;
	    RECT 2.1000 105.1000 2.4000 106.8000 ;
	    RECT 4.6000 106.1000 5.0000 106.8000 ;
	    RECT 6.2000 106.1000 6.6000 106.2000 ;
	    RECT 4.6000 105.8000 6.6000 106.1000 ;
	    RECT 3.0000 105.1000 3.4000 105.2000 ;
	    RECT 1.9000 104.8000 2.4000 105.1000 ;
	    RECT 2.7000 104.8000 3.4000 105.1000 ;
	    RECT 1.9000 101.1000 2.3000 104.8000 ;
	    RECT 2.7000 104.2000 3.0000 104.8000 ;
	    RECT 2.6000 103.8000 3.0000 104.2000 ;
	    RECT 4.6000 101.1000 5.0000 105.8000 ;
	    RECT 6.2000 105.4000 6.6000 105.8000 ;
	    RECT 7.0000 106.1000 7.3000 106.8000 ;
	    RECT 9.4000 106.4000 9.8000 107.2000 ;
	    RECT 8.6000 106.1000 9.0000 106.2000 ;
	    RECT 10.2000 106.1000 10.5000 107.9000 ;
	    RECT 11.0000 107.8000 11.4000 108.2000 ;
	    RECT 12.6000 107.9000 13.5000 108.2000 ;
	    RECT 14.2000 107.9000 14.6000 109.9000 ;
	    RECT 16.4000 108.1000 17.2000 109.9000 ;
	    RECT 11.8000 106.8000 12.2000 107.6000 ;
	    RECT 11.0000 106.1000 11.4000 106.2000 ;
	    RECT 7.0000 105.8000 9.4000 106.1000 ;
	    RECT 10.2000 105.8000 11.4000 106.1000 ;
	    RECT 5.4000 104.4000 5.8000 105.2000 ;
	    RECT 7.0000 105.1000 7.3000 105.8000 ;
	    RECT 9.0000 105.6000 9.4000 105.8000 ;
	    RECT 11.0000 105.1000 11.3000 105.8000 ;
	    RECT 6.5000 104.7000 7.4000 105.1000 ;
	    RECT 8.6000 104.8000 10.6000 105.1000 ;
	    RECT 6.5000 101.1000 6.9000 104.7000 ;
	    RECT 8.6000 101.1000 9.0000 104.8000 ;
	    RECT 10.2000 101.1000 10.6000 104.8000 ;
	    RECT 11.0000 101.1000 11.4000 105.1000 ;
	    RECT 12.6000 101.1000 13.0000 107.9000 ;
	    RECT 14.2000 107.6000 15.4000 107.9000 ;
	    RECT 15.0000 107.5000 15.4000 107.6000 ;
	    RECT 16.4000 106.4000 16.7000 108.1000 ;
	    RECT 19.0000 107.9000 19.4000 109.9000 ;
	    RECT 18.3000 107.6000 19.4000 107.9000 ;
	    RECT 18.3000 107.5000 18.7000 107.6000 ;
	    RECT 17.0000 106.7000 17.4000 107.1000 ;
	    RECT 16.2000 106.2000 16.7000 106.4000 ;
	    RECT 15.8000 106.1000 16.7000 106.2000 ;
	    RECT 17.1000 106.4000 17.4000 106.7000 ;
	    RECT 17.1000 106.1000 18.4000 106.4000 ;
	    RECT 15.8000 105.8000 16.5000 106.1000 ;
	    RECT 18.0000 106.0000 18.4000 106.1000 ;
	    RECT 20.6000 106.1000 21.0000 109.9000 ;
	    RECT 22.2000 108.9000 22.6000 109.9000 ;
	    RECT 22.3000 107.2000 22.6000 108.9000 ;
	    RECT 21.4000 106.8000 21.8000 107.2000 ;
	    RECT 22.2000 106.8000 22.6000 107.2000 ;
	    RECT 21.4000 106.1000 21.7000 106.8000 ;
	    RECT 20.6000 105.8000 21.7000 106.1000 ;
	    RECT 16.2000 105.2000 16.5000 105.8000 ;
	    RECT 16.9000 105.7000 17.3000 105.8000 ;
	    RECT 16.9000 105.4000 18.6000 105.7000 ;
	    RECT 13.4000 104.4000 13.8000 105.2000 ;
	    RECT 15.8000 105.1000 16.5000 105.2000 ;
	    RECT 18.3000 105.1000 18.6000 105.4000 ;
	    RECT 14.2000 104.8000 15.4000 105.1000 ;
	    RECT 15.8000 104.8000 17.2000 105.1000 ;
	    RECT 14.2000 101.1000 14.6000 104.8000 ;
	    RECT 15.0000 104.7000 15.4000 104.8000 ;
	    RECT 16.4000 101.1000 17.2000 104.8000 ;
	    RECT 18.3000 104.8000 19.4000 105.1000 ;
	    RECT 18.3000 104.7000 18.7000 104.8000 ;
	    RECT 19.0000 101.1000 19.4000 104.8000 ;
	    RECT 20.6000 101.1000 21.0000 105.8000 ;
	    RECT 22.3000 105.1000 22.6000 106.8000 ;
	    RECT 23.8000 107.7000 24.2000 109.9000 ;
	    RECT 25.9000 109.2000 26.5000 109.9000 ;
	    RECT 25.9000 108.9000 26.6000 109.2000 ;
	    RECT 28.2000 108.9000 28.6000 109.9000 ;
	    RECT 30.4000 109.2000 30.8000 109.9000 ;
	    RECT 30.4000 108.9000 31.4000 109.2000 ;
	    RECT 26.2000 108.5000 26.6000 108.9000 ;
	    RECT 28.3000 108.6000 28.6000 108.9000 ;
	    RECT 28.3000 108.3000 29.7000 108.6000 ;
	    RECT 29.3000 108.2000 29.7000 108.3000 ;
	    RECT 30.2000 107.8000 30.6000 108.6000 ;
	    RECT 31.0000 108.5000 31.4000 108.9000 ;
	    RECT 25.3000 107.7000 25.7000 107.8000 ;
	    RECT 23.8000 107.4000 25.7000 107.7000 ;
	    RECT 23.0000 105.4000 23.4000 106.2000 ;
	    RECT 23.8000 105.7000 24.2000 107.4000 ;
	    RECT 27.3000 107.1000 27.7000 107.2000 ;
	    RECT 30.2000 107.1000 30.5000 107.8000 ;
	    RECT 32.6000 107.5000 33.0000 109.9000 ;
	    RECT 33.4000 107.8000 33.8000 108.6000 ;
	    RECT 34.2000 108.1000 34.6000 109.9000 ;
	    RECT 35.8000 108.9000 36.2000 109.9000 ;
	    RECT 39.8000 108.9000 40.2000 109.9000 ;
	    RECT 41.4000 109.2000 41.8000 109.9000 ;
	    RECT 35.0000 108.1000 35.4000 108.6000 ;
	    RECT 34.2000 107.8000 35.4000 108.1000 ;
	    RECT 31.8000 107.1000 32.6000 107.2000 ;
	    RECT 27.1000 106.8000 32.6000 107.1000 ;
	    RECT 26.2000 106.4000 26.6000 106.5000 ;
	    RECT 24.7000 106.1000 26.6000 106.4000 ;
	    RECT 24.7000 106.0000 25.1000 106.1000 ;
	    RECT 25.5000 105.7000 25.9000 105.8000 ;
	    RECT 23.8000 105.4000 25.9000 105.7000 ;
	    RECT 22.2000 104.7000 23.1000 105.1000 ;
	    RECT 22.7000 102.2000 23.1000 104.7000 ;
	    RECT 22.7000 101.8000 23.4000 102.2000 ;
	    RECT 22.7000 101.1000 23.1000 101.8000 ;
	    RECT 23.8000 101.1000 24.2000 105.4000 ;
	    RECT 27.1000 105.2000 27.4000 106.8000 ;
	    RECT 30.7000 106.7000 31.1000 106.8000 ;
	    RECT 30.2000 106.2000 30.6000 106.3000 ;
	    RECT 31.5000 106.2000 31.9000 106.3000 ;
	    RECT 29.4000 105.9000 31.9000 106.2000 ;
	    RECT 29.4000 105.8000 29.8000 105.9000 ;
	    RECT 30.2000 105.5000 33.0000 105.6000 ;
	    RECT 30.1000 105.4000 33.0000 105.5000 ;
	    RECT 26.2000 104.9000 27.4000 105.2000 ;
	    RECT 28.1000 105.3000 33.0000 105.4000 ;
	    RECT 28.1000 105.1000 30.5000 105.3000 ;
	    RECT 26.2000 104.4000 26.5000 104.9000 ;
	    RECT 25.8000 104.0000 26.5000 104.4000 ;
	    RECT 27.3000 104.5000 27.7000 104.6000 ;
	    RECT 28.1000 104.5000 28.4000 105.1000 ;
	    RECT 27.3000 104.2000 28.4000 104.5000 ;
	    RECT 28.7000 104.5000 31.4000 104.8000 ;
	    RECT 28.7000 104.4000 29.1000 104.5000 ;
	    RECT 31.0000 104.4000 31.4000 104.5000 ;
	    RECT 27.9000 103.7000 28.3000 103.8000 ;
	    RECT 29.3000 103.7000 29.7000 103.8000 ;
	    RECT 26.2000 103.1000 26.6000 103.5000 ;
	    RECT 27.9000 103.4000 29.7000 103.7000 ;
	    RECT 28.3000 103.1000 28.6000 103.4000 ;
	    RECT 31.0000 103.1000 31.4000 103.5000 ;
	    RECT 25.9000 101.1000 26.5000 103.1000 ;
	    RECT 28.2000 101.1000 28.6000 103.1000 ;
	    RECT 30.4000 102.8000 31.4000 103.1000 ;
	    RECT 30.4000 101.1000 30.8000 102.8000 ;
	    RECT 32.6000 101.1000 33.0000 105.3000 ;
	    RECT 34.2000 101.1000 34.6000 107.8000 ;
	    RECT 35.9000 107.2000 36.2000 108.9000 ;
	    RECT 35.0000 106.8000 35.4000 107.2000 ;
	    RECT 35.8000 106.8000 36.2000 107.2000 ;
	    RECT 35.0000 106.1000 35.3000 106.8000 ;
	    RECT 35.9000 106.1000 36.2000 106.8000 ;
	    RECT 39.6000 108.8000 40.2000 108.9000 ;
	    RECT 41.3000 108.8000 41.8000 109.2000 ;
	    RECT 39.6000 108.5000 41.6000 108.8000 ;
	    RECT 35.0000 105.8000 36.2000 106.1000 ;
	    RECT 35.9000 105.1000 36.2000 105.8000 ;
	    RECT 36.6000 105.4000 37.0000 106.2000 ;
	    RECT 39.6000 105.2000 39.9000 108.5000 ;
	    RECT 41.7000 107.8000 42.6000 108.2000 ;
	    RECT 41.0000 107.1000 41.8000 107.2000 ;
	    RECT 43.8000 107.1000 44.2000 109.9000 ;
	    RECT 46.2000 108.9000 46.6000 109.9000 ;
	    RECT 44.6000 107.8000 45.0000 108.6000 ;
	    RECT 45.4000 107.8000 45.8000 108.6000 ;
	    RECT 41.0000 106.8000 44.2000 107.1000 ;
	    RECT 45.4000 107.2000 45.7000 107.8000 ;
	    RECT 46.3000 107.2000 46.6000 108.9000 ;
	    RECT 47.8000 108.0000 48.2000 109.9000 ;
	    RECT 49.4000 108.0000 49.8000 109.9000 ;
	    RECT 47.8000 107.9000 49.8000 108.0000 ;
	    RECT 50.2000 107.9000 50.6000 109.9000 ;
	    RECT 51.8000 108.9000 52.2000 109.9000 ;
	    RECT 51.0000 108.1000 51.4000 108.2000 ;
	    RECT 51.8000 108.1000 52.1000 108.9000 ;
	    RECT 47.9000 107.7000 49.7000 107.9000 ;
	    RECT 48.2000 107.2000 48.6000 107.4000 ;
	    RECT 50.2000 107.2000 50.5000 107.9000 ;
	    RECT 51.0000 107.8000 52.1000 108.1000 ;
	    RECT 52.6000 107.8000 53.0000 108.6000 ;
	    RECT 53.4000 107.9000 53.8000 109.9000 ;
	    RECT 54.2000 108.0000 54.6000 109.9000 ;
	    RECT 55.8000 108.0000 56.2000 109.9000 ;
	    RECT 58.3000 108.2000 58.7000 108.6000 ;
	    RECT 54.2000 107.9000 56.2000 108.0000 ;
	    RECT 51.8000 107.2000 52.1000 107.8000 ;
	    RECT 53.5000 107.2000 53.8000 107.9000 ;
	    RECT 54.3000 107.7000 56.1000 107.9000 ;
	    RECT 58.2000 107.8000 58.6000 108.2000 ;
	    RECT 59.0000 107.9000 59.4000 109.9000 ;
	    RECT 55.4000 107.2000 55.8000 107.4000 ;
	    RECT 45.4000 106.8000 45.8000 107.2000 ;
	    RECT 46.2000 107.1000 46.6000 107.2000 ;
	    RECT 47.8000 107.1000 48.6000 107.2000 ;
	    RECT 46.2000 106.9000 48.6000 107.1000 ;
	    RECT 46.2000 106.8000 48.2000 106.9000 ;
	    RECT 49.3000 106.8000 50.6000 107.2000 ;
	    RECT 51.8000 106.8000 52.2000 107.2000 ;
	    RECT 53.4000 106.8000 54.7000 107.2000 ;
	    RECT 55.4000 106.9000 56.2000 107.2000 ;
	    RECT 55.8000 106.8000 56.2000 106.9000 ;
	    RECT 40.2000 105.8000 41.0000 106.2000 ;
	    RECT 35.8000 104.7000 36.7000 105.1000 ;
	    RECT 38.2000 104.9000 39.9000 105.2000 ;
	    RECT 38.2000 104.8000 38.6000 104.9000 ;
	    RECT 36.3000 101.1000 36.7000 104.7000 ;
	    RECT 38.3000 104.5000 38.6000 104.8000 ;
	    RECT 39.1000 104.5000 40.9000 104.6000 ;
	    RECT 37.4000 101.5000 37.8000 104.5000 ;
	    RECT 38.2000 101.7000 38.6000 104.5000 ;
	    RECT 39.0000 104.3000 40.9000 104.5000 ;
	    RECT 37.5000 101.4000 37.8000 101.5000 ;
	    RECT 39.0000 101.5000 39.4000 104.3000 ;
	    RECT 40.6000 104.1000 40.9000 104.3000 ;
	    RECT 41.5000 104.4000 43.3000 104.7000 ;
	    RECT 41.5000 104.1000 41.8000 104.4000 ;
	    RECT 39.0000 101.4000 39.3000 101.5000 ;
	    RECT 37.5000 101.1000 39.3000 101.4000 ;
	    RECT 39.8000 101.4000 40.2000 104.0000 ;
	    RECT 40.6000 101.7000 41.0000 104.1000 ;
	    RECT 41.4000 101.4000 41.8000 104.1000 ;
	    RECT 39.8000 101.1000 41.8000 101.4000 ;
	    RECT 43.0000 104.1000 43.3000 104.4000 ;
	    RECT 43.0000 101.1000 43.4000 104.1000 ;
	    RECT 43.8000 101.1000 44.2000 106.8000 ;
	    RECT 46.3000 105.1000 46.6000 106.8000 ;
	    RECT 47.0000 106.1000 47.4000 106.2000 ;
	    RECT 47.8000 106.1000 48.2000 106.2000 ;
	    RECT 47.0000 105.8000 48.2000 106.1000 ;
	    RECT 48.6000 105.8000 49.0000 106.6000 ;
	    RECT 49.3000 106.1000 49.6000 106.8000 ;
	    RECT 51.0000 106.1000 51.4000 106.2000 ;
	    RECT 49.3000 105.8000 51.4000 106.1000 ;
	    RECT 47.0000 105.4000 47.4000 105.8000 ;
	    RECT 49.3000 105.1000 49.6000 105.8000 ;
	    RECT 51.0000 105.4000 51.4000 105.8000 ;
	    RECT 50.2000 105.1000 50.6000 105.2000 ;
	    RECT 51.8000 105.1000 52.1000 106.8000 ;
	    RECT 53.4000 105.1000 53.8000 105.2000 ;
	    RECT 54.4000 105.1000 54.7000 106.8000 ;
	    RECT 55.0000 105.8000 55.4000 106.6000 ;
	    RECT 58.2000 106.1000 58.6000 106.2000 ;
	    RECT 59.1000 106.1000 59.4000 107.9000 ;
	    RECT 63.0000 107.9000 63.4000 109.9000 ;
	    RECT 63.7000 108.2000 64.1000 108.6000 ;
	    RECT 59.8000 107.1000 60.2000 107.2000 ;
	    RECT 62.2000 107.1000 62.6000 107.2000 ;
	    RECT 59.8000 106.8000 62.6000 107.1000 ;
	    RECT 59.8000 106.4000 60.2000 106.8000 ;
	    RECT 62.2000 106.4000 62.6000 106.8000 ;
	    RECT 60.6000 106.1000 61.0000 106.2000 ;
	    RECT 61.4000 106.1000 61.8000 106.2000 ;
	    RECT 63.0000 106.1000 63.3000 107.9000 ;
	    RECT 63.8000 107.8000 64.2000 108.2000 ;
	    RECT 65.2000 107.1000 65.6000 109.9000 ;
	    RECT 64.7000 106.9000 65.6000 107.1000 ;
	    RECT 67.8000 107.7000 68.2000 109.9000 ;
	    RECT 69.9000 109.2000 70.5000 109.9000 ;
	    RECT 69.9000 108.9000 70.6000 109.2000 ;
	    RECT 72.2000 108.9000 72.6000 109.9000 ;
	    RECT 74.4000 109.2000 74.8000 109.9000 ;
	    RECT 74.4000 108.9000 75.4000 109.2000 ;
	    RECT 70.2000 108.5000 70.6000 108.9000 ;
	    RECT 72.3000 108.6000 72.6000 108.9000 ;
	    RECT 72.3000 108.3000 73.7000 108.6000 ;
	    RECT 73.3000 108.2000 73.7000 108.3000 ;
	    RECT 74.2000 108.2000 74.6000 108.6000 ;
	    RECT 75.0000 108.5000 75.4000 108.9000 ;
	    RECT 69.3000 107.7000 69.7000 107.8000 ;
	    RECT 67.8000 107.4000 69.7000 107.7000 ;
	    RECT 64.7000 106.8000 65.5000 106.9000 ;
	    RECT 63.8000 106.1000 64.2000 106.2000 ;
	    RECT 58.2000 105.8000 59.4000 106.1000 ;
	    RECT 60.2000 105.8000 62.2000 106.1000 ;
	    RECT 63.0000 105.8000 64.2000 106.1000 ;
	    RECT 58.3000 105.1000 58.6000 105.8000 ;
	    RECT 60.2000 105.6000 60.6000 105.8000 ;
	    RECT 61.8000 105.6000 62.2000 105.8000 ;
	    RECT 63.8000 105.1000 64.1000 105.8000 ;
	    RECT 64.7000 105.2000 65.0000 106.8000 ;
	    RECT 65.8000 105.8000 66.6000 106.2000 ;
	    RECT 67.8000 105.7000 68.2000 107.4000 ;
	    RECT 71.3000 107.1000 71.7000 107.2000 ;
	    RECT 74.2000 107.1000 74.5000 108.2000 ;
	    RECT 76.6000 107.5000 77.0000 109.9000 ;
	    RECT 77.5000 108.2000 77.9000 108.6000 ;
	    RECT 77.4000 107.8000 77.8000 108.2000 ;
	    RECT 78.2000 107.9000 78.6000 109.9000 ;
	    RECT 80.6000 107.9000 81.0000 109.9000 ;
	    RECT 81.4000 108.0000 81.8000 109.9000 ;
	    RECT 83.0000 108.0000 83.4000 109.9000 ;
	    RECT 83.9000 108.2000 84.3000 108.6000 ;
	    RECT 81.4000 107.9000 83.4000 108.0000 ;
	    RECT 75.8000 107.1000 76.6000 107.2000 ;
	    RECT 71.1000 106.8000 76.6000 107.1000 ;
	    RECT 77.4000 106.8000 77.8000 107.2000 ;
	    RECT 70.2000 106.4000 70.6000 106.5000 ;
	    RECT 68.7000 106.1000 70.6000 106.4000 ;
	    RECT 71.1000 106.2000 71.4000 106.8000 ;
	    RECT 74.7000 106.7000 75.1000 106.8000 ;
	    RECT 74.2000 106.2000 74.6000 106.3000 ;
	    RECT 75.5000 106.2000 75.9000 106.3000 ;
	    RECT 68.7000 106.0000 69.1000 106.1000 ;
	    RECT 71.0000 105.8000 71.4000 106.2000 ;
	    RECT 73.4000 105.9000 75.9000 106.2000 ;
	    RECT 77.4000 106.2000 77.7000 106.8000 ;
	    RECT 77.4000 106.1000 77.8000 106.2000 ;
	    RECT 78.3000 106.1000 78.6000 107.9000 ;
	    RECT 80.7000 107.2000 81.0000 107.9000 ;
	    RECT 81.5000 107.7000 83.3000 107.9000 ;
	    RECT 83.8000 107.8000 84.2000 108.2000 ;
	    RECT 84.6000 107.9000 85.0000 109.9000 ;
	    RECT 87.0000 107.9000 87.4000 109.9000 ;
	    RECT 87.8000 108.0000 88.2000 109.9000 ;
	    RECT 89.4000 108.0000 89.8000 109.9000 ;
	    RECT 91.5000 108.2000 91.9000 109.9000 ;
	    RECT 87.8000 107.9000 89.8000 108.0000 ;
	    RECT 91.0000 107.9000 91.9000 108.2000 ;
	    RECT 82.6000 107.2000 83.0000 107.4000 ;
	    RECT 79.0000 107.1000 79.4000 107.2000 ;
	    RECT 80.6000 107.1000 81.9000 107.2000 ;
	    RECT 79.0000 106.8000 81.9000 107.1000 ;
	    RECT 82.6000 106.9000 83.4000 107.2000 ;
	    RECT 83.0000 106.8000 83.4000 106.9000 ;
	    RECT 79.0000 106.4000 79.4000 106.8000 ;
	    RECT 79.8000 106.1000 80.2000 106.2000 ;
	    RECT 73.4000 105.8000 73.8000 105.9000 ;
	    RECT 77.4000 105.8000 78.6000 106.1000 ;
	    RECT 79.4000 105.8000 80.2000 106.1000 ;
	    RECT 69.5000 105.7000 69.9000 105.8000 ;
	    RECT 46.2000 104.7000 47.1000 105.1000 ;
	    RECT 46.7000 102.2000 47.1000 104.7000 ;
	    RECT 49.1000 104.8000 49.6000 105.1000 ;
	    RECT 49.9000 104.8000 50.6000 105.1000 ;
	    RECT 46.7000 101.8000 47.4000 102.2000 ;
	    RECT 46.7000 101.1000 47.1000 101.8000 ;
	    RECT 49.1000 101.1000 49.5000 104.8000 ;
	    RECT 49.9000 104.2000 50.2000 104.8000 ;
	    RECT 49.8000 103.8000 50.2000 104.2000 ;
	    RECT 51.3000 104.7000 52.2000 105.1000 ;
	    RECT 53.4000 104.8000 54.1000 105.1000 ;
	    RECT 54.4000 104.8000 54.9000 105.1000 ;
	    RECT 51.3000 101.1000 51.7000 104.7000 ;
	    RECT 53.8000 104.2000 54.1000 104.8000 ;
	    RECT 53.8000 103.8000 54.2000 104.2000 ;
	    RECT 54.5000 101.1000 54.9000 104.8000 ;
	    RECT 57.4000 102.1000 57.8000 102.2000 ;
	    RECT 58.2000 102.1000 58.6000 105.1000 ;
	    RECT 57.4000 101.8000 58.6000 102.1000 ;
	    RECT 58.2000 101.1000 58.6000 101.8000 ;
	    RECT 59.0000 104.8000 61.0000 105.1000 ;
	    RECT 59.0000 101.1000 59.4000 104.8000 ;
	    RECT 60.6000 101.1000 61.0000 104.8000 ;
	    RECT 61.4000 104.8000 63.4000 105.1000 ;
	    RECT 61.4000 101.1000 61.8000 104.8000 ;
	    RECT 63.0000 101.1000 63.4000 104.8000 ;
	    RECT 63.8000 101.1000 64.2000 105.1000 ;
	    RECT 64.6000 104.8000 65.0000 105.2000 ;
	    RECT 67.0000 105.1000 67.4000 105.6000 ;
	    RECT 67.8000 105.4000 69.9000 105.7000 ;
	    RECT 67.8000 105.1000 68.2000 105.4000 ;
	    RECT 71.1000 105.2000 71.4000 105.8000 ;
	    RECT 74.2000 105.5000 77.0000 105.6000 ;
	    RECT 74.1000 105.4000 77.0000 105.5000 ;
	    RECT 67.0000 104.8000 68.2000 105.1000 ;
	    RECT 64.7000 103.5000 65.0000 104.8000 ;
	    RECT 65.4000 103.8000 65.8000 104.6000 ;
	    RECT 64.7000 103.2000 66.5000 103.5000 ;
	    RECT 64.7000 103.1000 65.0000 103.2000 ;
	    RECT 64.6000 101.1000 65.0000 103.1000 ;
	    RECT 66.2000 103.1000 66.5000 103.2000 ;
	    RECT 66.2000 101.1000 66.6000 103.1000 ;
	    RECT 67.8000 101.1000 68.2000 104.8000 ;
	    RECT 70.2000 104.9000 71.4000 105.2000 ;
	    RECT 72.1000 105.3000 77.0000 105.4000 ;
	    RECT 72.1000 105.1000 74.5000 105.3000 ;
	    RECT 70.2000 104.4000 70.5000 104.9000 ;
	    RECT 69.8000 104.0000 70.5000 104.4000 ;
	    RECT 71.3000 104.5000 71.7000 104.6000 ;
	    RECT 72.1000 104.5000 72.4000 105.1000 ;
	    RECT 71.3000 104.2000 72.4000 104.5000 ;
	    RECT 72.7000 104.5000 75.4000 104.8000 ;
	    RECT 72.7000 104.4000 73.1000 104.5000 ;
	    RECT 75.0000 104.4000 75.4000 104.5000 ;
	    RECT 71.9000 103.7000 72.3000 103.8000 ;
	    RECT 73.3000 103.7000 73.7000 103.8000 ;
	    RECT 70.2000 103.1000 70.6000 103.5000 ;
	    RECT 71.9000 103.4000 73.7000 103.7000 ;
	    RECT 72.3000 103.1000 72.6000 103.4000 ;
	    RECT 75.0000 103.1000 75.4000 103.5000 ;
	    RECT 69.9000 101.1000 70.5000 103.1000 ;
	    RECT 72.2000 101.1000 72.6000 103.1000 ;
	    RECT 74.4000 102.8000 75.4000 103.1000 ;
	    RECT 74.4000 101.1000 74.8000 102.8000 ;
	    RECT 76.6000 101.1000 77.0000 105.3000 ;
	    RECT 77.5000 105.1000 77.8000 105.8000 ;
	    RECT 79.4000 105.6000 79.8000 105.8000 ;
	    RECT 80.6000 105.1000 81.0000 105.2000 ;
	    RECT 81.6000 105.1000 81.9000 106.8000 ;
	    RECT 82.2000 105.8000 82.6000 106.6000 ;
	    RECT 83.8000 106.1000 84.2000 106.2000 ;
	    RECT 84.7000 106.1000 85.0000 107.9000 ;
	    RECT 87.1000 107.2000 87.4000 107.9000 ;
	    RECT 87.9000 107.7000 89.7000 107.9000 ;
	    RECT 89.0000 107.2000 89.4000 107.4000 ;
	    RECT 85.4000 107.1000 85.8000 107.2000 ;
	    RECT 87.0000 107.1000 88.3000 107.2000 ;
	    RECT 85.4000 106.8000 88.3000 107.1000 ;
	    RECT 89.0000 106.9000 89.8000 107.2000 ;
	    RECT 89.4000 106.8000 89.8000 106.9000 ;
	    RECT 90.2000 106.8000 90.6000 107.6000 ;
	    RECT 85.4000 106.4000 85.8000 106.8000 ;
	    RECT 86.2000 106.1000 86.6000 106.2000 ;
	    RECT 83.8000 105.8000 85.0000 106.1000 ;
	    RECT 85.8000 105.8000 86.6000 106.1000 ;
	    RECT 83.9000 105.1000 84.2000 105.8000 ;
	    RECT 85.8000 105.6000 86.2000 105.8000 ;
	    RECT 87.0000 105.1000 87.4000 105.2000 ;
	    RECT 88.0000 105.1000 88.3000 106.8000 ;
	    RECT 88.6000 106.1000 89.0000 106.6000 ;
	    RECT 89.4000 106.1000 89.8000 106.2000 ;
	    RECT 88.6000 105.8000 89.8000 106.1000 ;
	    RECT 90.2000 105.1000 90.6000 105.2000 ;
	    RECT 91.0000 105.1000 91.4000 107.9000 ;
	    RECT 77.4000 101.1000 77.8000 105.1000 ;
	    RECT 78.2000 104.8000 80.2000 105.1000 ;
	    RECT 80.6000 104.8000 81.3000 105.1000 ;
	    RECT 81.6000 104.8000 82.1000 105.1000 ;
	    RECT 78.2000 101.1000 78.6000 104.8000 ;
	    RECT 79.8000 101.1000 80.2000 104.8000 ;
	    RECT 81.0000 104.2000 81.3000 104.8000 ;
	    RECT 80.6000 103.8000 81.4000 104.2000 ;
	    RECT 81.7000 101.1000 82.1000 104.8000 ;
	    RECT 83.8000 101.1000 84.2000 105.1000 ;
	    RECT 84.6000 104.8000 86.6000 105.1000 ;
	    RECT 87.0000 104.8000 87.7000 105.1000 ;
	    RECT 88.0000 104.8000 88.5000 105.1000 ;
	    RECT 90.2000 104.8000 91.4000 105.1000 ;
	    RECT 84.6000 101.1000 85.0000 104.8000 ;
	    RECT 86.2000 101.1000 86.6000 104.8000 ;
	    RECT 87.4000 104.2000 87.7000 104.8000 ;
	    RECT 87.4000 103.8000 87.8000 104.2000 ;
	    RECT 88.1000 101.1000 88.5000 104.8000 ;
	    RECT 91.0000 101.1000 91.4000 104.8000 ;
	    RECT 91.8000 105.1000 92.2000 105.2000 ;
	    RECT 92.6000 105.1000 93.0000 109.9000 ;
	    RECT 93.4000 107.8000 93.8000 108.6000 ;
	    RECT 94.8000 107.2000 95.2000 109.9000 ;
	    RECT 98.2000 108.9000 98.6000 109.9000 ;
	    RECT 100.6000 108.9000 101.0000 109.9000 ;
	    RECT 95.8000 107.8000 96.2000 108.2000 ;
	    RECT 94.8000 107.1000 95.4000 107.2000 ;
	    RECT 95.8000 107.1000 96.1000 107.8000 ;
	    RECT 94.3000 106.8000 96.1000 107.1000 ;
	    RECT 98.2000 107.2000 98.5000 108.9000 ;
	    RECT 99.0000 107.8000 99.4000 108.6000 ;
	    RECT 99.8000 107.8000 100.2000 108.6000 ;
	    RECT 100.7000 107.8000 101.0000 108.9000 ;
	    RECT 102.2000 107.9000 102.6000 109.9000 ;
	    RECT 103.0000 108.0000 103.4000 109.9000 ;
	    RECT 104.6000 108.0000 105.0000 109.9000 ;
	    RECT 103.0000 107.9000 105.0000 108.0000 ;
	    RECT 105.4000 107.9000 105.8000 109.9000 ;
	    RECT 100.7000 107.5000 101.9000 107.8000 ;
	    RECT 98.2000 106.8000 98.6000 107.2000 ;
	    RECT 100.6000 106.8000 101.1000 107.2000 ;
	    RECT 94.3000 105.2000 94.6000 106.8000 ;
	    RECT 95.4000 105.8000 96.2000 106.2000 ;
	    RECT 91.8000 104.8000 93.0000 105.1000 ;
	    RECT 94.2000 104.8000 94.6000 105.2000 ;
	    RECT 96.6000 104.8000 97.0000 105.6000 ;
	    RECT 97.4000 105.4000 97.8000 106.2000 ;
	    RECT 98.2000 105.1000 98.5000 106.8000 ;
	    RECT 100.8000 106.4000 101.2000 106.8000 ;
	    RECT 101.6000 106.0000 101.9000 107.5000 ;
	    RECT 102.3000 106.2000 102.6000 107.9000 ;
	    RECT 103.1000 107.7000 104.9000 107.9000 ;
	    RECT 103.4000 107.2000 103.8000 107.4000 ;
	    RECT 105.4000 107.2000 105.7000 107.9000 ;
	    RECT 106.8000 107.2000 107.2000 109.9000 ;
	    RECT 112.3000 107.9000 113.1000 109.9000 ;
	    RECT 116.6000 107.9000 117.0000 109.9000 ;
	    RECT 119.0000 108.9000 119.4000 109.9000 ;
	    RECT 117.3000 108.2000 117.7000 108.6000 ;
	    RECT 119.0000 108.2000 119.3000 108.9000 ;
	    RECT 117.4000 108.1000 117.8000 108.2000 ;
	    RECT 118.2000 108.1000 118.6000 108.2000 ;
	    RECT 103.0000 106.9000 103.8000 107.2000 ;
	    RECT 103.0000 106.8000 103.4000 106.9000 ;
	    RECT 104.5000 106.8000 105.8000 107.2000 ;
	    RECT 106.2000 106.9000 107.2000 107.2000 ;
	    RECT 111.0000 107.1000 111.4000 107.2000 ;
	    RECT 111.8000 107.1000 112.2000 107.2000 ;
	    RECT 106.2000 106.8000 107.1000 106.9000 ;
	    RECT 111.0000 106.8000 112.2000 107.1000 ;
	    RECT 101.5000 105.7000 101.9000 106.0000 ;
	    RECT 102.2000 106.1000 102.6000 106.2000 ;
	    RECT 103.8000 106.1000 104.2000 106.6000 ;
	    RECT 102.2000 105.8000 104.2000 106.1000 ;
	    RECT 99.8000 105.6000 101.9000 105.7000 ;
	    RECT 99.8000 105.4000 101.8000 105.6000 ;
	    RECT 91.8000 104.4000 92.2000 104.8000 ;
	    RECT 92.6000 101.1000 93.0000 104.8000 ;
	    RECT 94.3000 103.5000 94.6000 104.8000 ;
	    RECT 97.7000 104.7000 98.6000 105.1000 ;
	    RECT 95.0000 103.8000 95.4000 104.6000 ;
	    RECT 94.3000 103.2000 96.1000 103.5000 ;
	    RECT 94.3000 103.1000 94.6000 103.2000 ;
	    RECT 94.2000 101.1000 94.6000 103.1000 ;
	    RECT 95.8000 103.1000 96.1000 103.2000 ;
	    RECT 95.8000 101.1000 96.2000 103.1000 ;
	    RECT 97.7000 102.2000 98.1000 104.7000 ;
	    RECT 97.7000 101.8000 98.6000 102.2000 ;
	    RECT 97.7000 101.1000 98.1000 101.8000 ;
	    RECT 99.8000 101.1000 100.2000 105.4000 ;
	    RECT 102.3000 105.1000 102.6000 105.8000 ;
	    RECT 104.5000 105.1000 104.8000 106.8000 ;
	    RECT 106.3000 105.2000 106.6000 106.8000 ;
	    RECT 111.9000 106.6000 112.2000 106.8000 ;
	    RECT 111.9000 106.2000 112.3000 106.6000 ;
	    RECT 112.6000 106.2000 112.9000 107.9000 ;
	    RECT 113.4000 107.1000 113.8000 107.2000 ;
	    RECT 115.8000 107.1000 116.2000 107.2000 ;
	    RECT 113.4000 106.8000 116.2000 107.1000 ;
	    RECT 113.4000 106.4000 113.8000 106.8000 ;
	    RECT 115.8000 106.4000 116.2000 106.8000 ;
	    RECT 107.4000 105.8000 108.2000 106.2000 ;
	    RECT 105.4000 105.1000 105.8000 105.2000 ;
	    RECT 101.9000 104.8000 102.6000 105.1000 ;
	    RECT 104.3000 104.8000 104.8000 105.1000 ;
	    RECT 105.1000 104.8000 105.8000 105.1000 ;
	    RECT 106.2000 104.8000 106.6000 105.2000 ;
	    RECT 108.6000 104.8000 109.0000 105.6000 ;
	    RECT 111.0000 105.4000 111.4000 106.2000 ;
	    RECT 112.6000 105.8000 113.0000 106.2000 ;
	    RECT 114.2000 106.1000 114.6000 106.2000 ;
	    RECT 115.0000 106.1000 115.4000 106.2000 ;
	    RECT 116.6000 106.1000 116.9000 107.9000 ;
	    RECT 117.4000 107.8000 118.6000 108.1000 ;
	    RECT 119.0000 107.8000 119.4000 108.2000 ;
	    RECT 119.8000 108.1000 120.2000 108.6000 ;
	    RECT 120.6000 108.1000 121.0000 109.9000 ;
	    RECT 119.8000 107.8000 121.0000 108.1000 ;
	    RECT 121.4000 108.0000 121.8000 109.9000 ;
	    RECT 123.0000 108.0000 123.4000 109.9000 ;
	    RECT 121.4000 107.9000 123.4000 108.0000 ;
	    RECT 119.0000 107.2000 119.3000 107.8000 ;
	    RECT 120.7000 107.2000 121.0000 107.8000 ;
	    RECT 121.5000 107.7000 123.3000 107.9000 ;
	    RECT 123.8000 107.7000 124.2000 109.9000 ;
	    RECT 125.9000 109.2000 126.5000 109.9000 ;
	    RECT 125.9000 108.9000 126.6000 109.2000 ;
	    RECT 128.2000 108.9000 128.6000 109.9000 ;
	    RECT 130.4000 109.2000 130.8000 109.9000 ;
	    RECT 130.4000 108.9000 131.4000 109.2000 ;
	    RECT 126.2000 108.5000 126.6000 108.9000 ;
	    RECT 128.3000 108.6000 128.6000 108.9000 ;
	    RECT 128.3000 108.3000 129.7000 108.6000 ;
	    RECT 129.3000 108.2000 129.7000 108.3000 ;
	    RECT 130.2000 108.2000 130.6000 108.6000 ;
	    RECT 131.0000 108.5000 131.4000 108.9000 ;
	    RECT 125.3000 107.7000 125.7000 107.8000 ;
	    RECT 123.8000 107.4000 125.7000 107.7000 ;
	    RECT 122.6000 107.2000 123.0000 107.4000 ;
	    RECT 119.0000 106.8000 119.4000 107.2000 ;
	    RECT 120.6000 106.8000 121.9000 107.2000 ;
	    RECT 122.6000 106.9000 123.4000 107.2000 ;
	    RECT 123.0000 106.8000 123.4000 106.9000 ;
	    RECT 117.4000 106.1000 117.8000 106.2000 ;
	    RECT 118.2000 106.1000 118.6000 106.2000 ;
	    RECT 113.8000 105.8000 115.8000 106.1000 ;
	    RECT 116.6000 105.8000 118.6000 106.1000 ;
	    RECT 112.6000 105.7000 112.9000 105.8000 ;
	    RECT 111.9000 105.4000 112.9000 105.7000 ;
	    RECT 113.8000 105.6000 114.2000 105.8000 ;
	    RECT 115.4000 105.6000 115.8000 105.8000 ;
	    RECT 111.9000 105.1000 112.2000 105.4000 ;
	    RECT 117.4000 105.1000 117.7000 105.8000 ;
	    RECT 118.2000 105.4000 118.6000 105.8000 ;
	    RECT 119.0000 105.1000 119.3000 106.8000 ;
	    RECT 120.6000 105.1000 121.0000 105.2000 ;
	    RECT 121.6000 105.1000 121.9000 106.8000 ;
	    RECT 122.2000 105.8000 122.6000 106.6000 ;
	    RECT 123.8000 105.7000 124.2000 107.4000 ;
	    RECT 127.0000 107.1000 127.7000 107.2000 ;
	    RECT 129.4000 107.1000 129.8000 107.2000 ;
	    RECT 130.2000 107.1000 130.5000 108.2000 ;
	    RECT 132.6000 107.5000 133.0000 109.9000 ;
	    RECT 133.4000 107.7000 133.8000 109.9000 ;
	    RECT 135.5000 109.2000 136.1000 109.9000 ;
	    RECT 135.5000 108.9000 136.2000 109.2000 ;
	    RECT 137.8000 108.9000 138.2000 109.9000 ;
	    RECT 140.0000 109.2000 140.4000 109.9000 ;
	    RECT 140.0000 108.9000 141.0000 109.2000 ;
	    RECT 135.8000 108.5000 136.2000 108.9000 ;
	    RECT 137.9000 108.6000 138.2000 108.9000 ;
	    RECT 137.9000 108.3000 139.3000 108.6000 ;
	    RECT 138.9000 108.2000 139.3000 108.3000 ;
	    RECT 139.8000 108.2000 140.2000 108.6000 ;
	    RECT 140.6000 108.5000 141.0000 108.9000 ;
	    RECT 134.9000 107.7000 135.3000 107.8000 ;
	    RECT 133.4000 107.4000 135.3000 107.7000 ;
	    RECT 131.8000 107.1000 132.6000 107.2000 ;
	    RECT 127.0000 106.8000 132.6000 107.1000 ;
	    RECT 126.2000 106.4000 126.6000 106.5000 ;
	    RECT 124.7000 106.1000 126.6000 106.4000 ;
	    RECT 124.7000 106.0000 125.1000 106.1000 ;
	    RECT 125.5000 105.7000 125.9000 105.8000 ;
	    RECT 123.8000 105.4000 125.9000 105.7000 ;
	    RECT 101.9000 101.1000 102.3000 104.8000 ;
	    RECT 104.3000 102.2000 104.7000 104.8000 ;
	    RECT 105.1000 104.2000 105.4000 104.8000 ;
	    RECT 105.0000 103.8000 105.4000 104.2000 ;
	    RECT 106.3000 103.5000 106.6000 104.8000 ;
	    RECT 107.0000 103.8000 107.4000 104.6000 ;
	    RECT 106.3000 103.2000 108.1000 103.5000 ;
	    RECT 106.3000 103.1000 106.6000 103.2000 ;
	    RECT 103.8000 101.8000 104.7000 102.2000 ;
	    RECT 104.3000 101.1000 104.7000 101.8000 ;
	    RECT 106.2000 101.1000 106.6000 103.1000 ;
	    RECT 107.8000 103.1000 108.1000 103.2000 ;
	    RECT 107.8000 101.1000 108.2000 103.1000 ;
	    RECT 111.0000 101.4000 111.4000 105.1000 ;
	    RECT 111.8000 101.7000 112.2000 105.1000 ;
	    RECT 112.6000 104.8000 114.6000 105.1000 ;
	    RECT 112.6000 101.4000 113.0000 104.8000 ;
	    RECT 111.0000 101.1000 113.0000 101.4000 ;
	    RECT 114.2000 101.1000 114.6000 104.8000 ;
	    RECT 115.0000 104.8000 117.0000 105.1000 ;
	    RECT 115.0000 101.1000 115.4000 104.8000 ;
	    RECT 116.6000 101.1000 117.0000 104.8000 ;
	    RECT 117.4000 101.1000 117.8000 105.1000 ;
	    RECT 118.5000 104.7000 119.4000 105.1000 ;
	    RECT 120.6000 104.8000 121.3000 105.1000 ;
	    RECT 121.6000 104.8000 122.1000 105.1000 ;
	    RECT 118.5000 101.1000 118.9000 104.7000 ;
	    RECT 121.0000 104.2000 121.3000 104.8000 ;
	    RECT 121.0000 103.8000 121.4000 104.2000 ;
	    RECT 121.7000 101.1000 122.1000 104.8000 ;
	    RECT 123.8000 101.1000 124.2000 105.4000 ;
	    RECT 127.1000 105.2000 127.4000 106.8000 ;
	    RECT 130.7000 106.7000 131.1000 106.8000 ;
	    RECT 130.2000 106.2000 130.6000 106.3000 ;
	    RECT 131.5000 106.2000 131.9000 106.3000 ;
	    RECT 129.4000 105.9000 131.9000 106.2000 ;
	    RECT 129.4000 105.8000 129.8000 105.9000 ;
	    RECT 133.4000 105.7000 133.8000 107.4000 ;
	    RECT 136.9000 107.1000 137.3000 107.2000 ;
	    RECT 139.8000 107.1000 140.1000 108.2000 ;
	    RECT 142.2000 107.5000 142.6000 109.9000 ;
	    RECT 143.8000 108.9000 144.2000 109.9000 ;
	    RECT 147.8000 108.9000 148.2000 109.9000 ;
	    RECT 149.4000 109.2000 149.8000 109.9000 ;
	    RECT 143.8000 107.2000 144.1000 108.9000 ;
	    RECT 147.6000 108.8000 148.2000 108.9000 ;
	    RECT 149.3000 108.8000 149.8000 109.2000 ;
	    RECT 152.1000 109.1000 152.5000 109.9000 ;
	    RECT 151.0000 108.8000 152.5000 109.1000 ;
	    RECT 144.6000 107.8000 145.0000 108.6000 ;
	    RECT 147.6000 108.5000 149.6000 108.8000 ;
	    RECT 141.4000 107.1000 142.2000 107.2000 ;
	    RECT 136.7000 106.8000 142.2000 107.1000 ;
	    RECT 143.8000 106.8000 144.2000 107.2000 ;
	    RECT 135.8000 106.4000 136.2000 106.5000 ;
	    RECT 134.3000 106.1000 136.2000 106.4000 ;
	    RECT 136.7000 106.2000 137.0000 106.8000 ;
	    RECT 140.3000 106.7000 140.7000 106.8000 ;
	    RECT 139.8000 106.2000 140.2000 106.3000 ;
	    RECT 141.1000 106.2000 141.5000 106.3000 ;
	    RECT 134.3000 106.0000 134.7000 106.1000 ;
	    RECT 136.6000 105.8000 137.0000 106.2000 ;
	    RECT 139.0000 105.9000 141.5000 106.2000 ;
	    RECT 139.0000 105.8000 139.4000 105.9000 ;
	    RECT 135.1000 105.7000 135.5000 105.8000 ;
	    RECT 130.2000 105.5000 133.0000 105.6000 ;
	    RECT 130.1000 105.4000 133.0000 105.5000 ;
	    RECT 126.2000 104.9000 127.4000 105.2000 ;
	    RECT 128.1000 105.3000 133.0000 105.4000 ;
	    RECT 128.1000 105.1000 130.5000 105.3000 ;
	    RECT 126.2000 104.4000 126.5000 104.9000 ;
	    RECT 125.8000 104.0000 126.5000 104.4000 ;
	    RECT 127.3000 104.5000 127.7000 104.6000 ;
	    RECT 128.1000 104.5000 128.4000 105.1000 ;
	    RECT 127.3000 104.2000 128.4000 104.5000 ;
	    RECT 128.7000 104.5000 131.4000 104.8000 ;
	    RECT 128.7000 104.4000 129.1000 104.5000 ;
	    RECT 131.0000 104.4000 131.4000 104.5000 ;
	    RECT 127.9000 103.7000 128.3000 103.8000 ;
	    RECT 129.3000 103.7000 129.7000 103.8000 ;
	    RECT 126.2000 103.1000 126.6000 103.5000 ;
	    RECT 127.9000 103.4000 129.7000 103.7000 ;
	    RECT 128.3000 103.1000 128.6000 103.4000 ;
	    RECT 131.0000 103.1000 131.4000 103.5000 ;
	    RECT 125.9000 101.1000 126.5000 103.1000 ;
	    RECT 128.2000 101.1000 128.6000 103.1000 ;
	    RECT 130.4000 102.8000 131.4000 103.1000 ;
	    RECT 130.4000 101.1000 130.8000 102.8000 ;
	    RECT 132.6000 101.1000 133.0000 105.3000 ;
	    RECT 133.4000 105.4000 135.5000 105.7000 ;
	    RECT 133.4000 101.1000 133.8000 105.4000 ;
	    RECT 136.7000 105.2000 137.0000 105.8000 ;
	    RECT 139.8000 105.5000 142.6000 105.6000 ;
	    RECT 139.7000 105.4000 142.6000 105.5000 ;
	    RECT 143.0000 105.4000 143.4000 106.2000 ;
	    RECT 143.8000 106.1000 144.1000 106.8000 ;
	    RECT 144.6000 106.1000 145.0000 106.2000 ;
	    RECT 143.8000 105.8000 145.0000 106.1000 ;
	    RECT 135.8000 104.9000 137.0000 105.2000 ;
	    RECT 137.7000 105.3000 142.6000 105.4000 ;
	    RECT 137.7000 105.1000 140.1000 105.3000 ;
	    RECT 135.8000 104.4000 136.1000 104.9000 ;
	    RECT 135.4000 104.0000 136.1000 104.4000 ;
	    RECT 136.9000 104.5000 137.3000 104.6000 ;
	    RECT 137.7000 104.5000 138.0000 105.1000 ;
	    RECT 136.9000 104.2000 138.0000 104.5000 ;
	    RECT 138.3000 104.5000 141.0000 104.8000 ;
	    RECT 138.3000 104.4000 138.7000 104.5000 ;
	    RECT 140.6000 104.4000 141.0000 104.5000 ;
	    RECT 137.5000 103.7000 137.9000 103.8000 ;
	    RECT 138.9000 103.7000 139.3000 103.8000 ;
	    RECT 135.8000 103.1000 136.2000 103.5000 ;
	    RECT 137.5000 103.4000 139.3000 103.7000 ;
	    RECT 137.9000 103.1000 138.2000 103.4000 ;
	    RECT 140.6000 103.1000 141.0000 103.5000 ;
	    RECT 135.5000 101.1000 136.1000 103.1000 ;
	    RECT 137.8000 101.1000 138.2000 103.1000 ;
	    RECT 140.0000 102.8000 141.0000 103.1000 ;
	    RECT 140.0000 101.1000 140.4000 102.8000 ;
	    RECT 142.2000 101.1000 142.6000 105.3000 ;
	    RECT 143.8000 105.1000 144.1000 105.8000 ;
	    RECT 147.6000 105.2000 147.9000 108.5000 ;
	    RECT 149.7000 108.1000 150.6000 108.2000 ;
	    RECT 151.0000 108.1000 151.3000 108.8000 ;
	    RECT 152.1000 108.4000 152.5000 108.8000 ;
	    RECT 149.7000 107.8000 151.3000 108.1000 ;
	    RECT 151.8000 107.9000 152.5000 108.4000 ;
	    RECT 154.2000 107.9000 154.6000 109.9000 ;
	    RECT 155.8000 108.9000 156.2000 109.9000 ;
	    RECT 149.0000 107.1000 149.8000 107.2000 ;
	    RECT 150.2000 107.1000 150.6000 107.2000 ;
	    RECT 149.0000 106.8000 150.6000 107.1000 ;
	    RECT 151.8000 106.2000 152.1000 107.9000 ;
	    RECT 154.2000 107.8000 154.5000 107.9000 ;
	    RECT 155.0000 107.8000 155.4000 108.6000 ;
	    RECT 155.9000 107.8000 156.2000 108.9000 ;
	    RECT 157.4000 107.9000 157.8000 109.9000 ;
	    RECT 153.6000 107.6000 154.5000 107.8000 ;
	    RECT 152.4000 107.5000 154.5000 107.6000 ;
	    RECT 155.9000 107.5000 157.1000 107.8000 ;
	    RECT 152.4000 107.3000 153.9000 107.5000 ;
	    RECT 152.4000 107.2000 152.8000 107.3000 ;
	    RECT 148.2000 105.8000 149.0000 106.2000 ;
	    RECT 151.8000 105.8000 152.2000 106.2000 ;
	    RECT 143.3000 104.7000 144.2000 105.1000 ;
	    RECT 146.2000 104.9000 147.9000 105.2000 ;
	    RECT 151.8000 105.1000 152.1000 105.8000 ;
	    RECT 152.5000 105.5000 152.8000 107.2000 ;
	    RECT 154.2000 107.1000 154.6000 107.2000 ;
	    RECT 155.0000 107.1000 155.4000 107.2000 ;
	    RECT 153.2000 106.6000 153.8000 107.0000 ;
	    RECT 154.2000 106.8000 155.4000 107.1000 ;
	    RECT 155.8000 106.8000 156.3000 107.2000 ;
	    RECT 153.4000 106.2000 153.7000 106.6000 ;
	    RECT 154.2000 106.4000 154.6000 106.8000 ;
	    RECT 156.0000 106.4000 156.4000 106.8000 ;
	    RECT 153.4000 105.8000 153.8000 106.2000 ;
	    RECT 156.8000 106.0000 157.1000 107.5000 ;
	    RECT 157.5000 107.1000 157.8000 107.9000 ;
	    RECT 159.8000 107.9000 160.2000 109.9000 ;
	    RECT 160.5000 108.2000 160.9000 108.6000 ;
	    RECT 160.6000 108.1000 161.0000 108.2000 ;
	    RECT 162.2000 108.1000 162.6000 108.2000 ;
	    RECT 159.0000 107.1000 159.4000 107.2000 ;
	    RECT 157.4000 106.8000 159.4000 107.1000 ;
	    RECT 157.5000 106.2000 157.8000 106.8000 ;
	    RECT 159.0000 106.4000 159.4000 106.8000 ;
	    RECT 156.7000 105.7000 157.1000 106.0000 ;
	    RECT 157.4000 105.8000 157.8000 106.2000 ;
	    RECT 158.2000 106.1000 158.6000 106.2000 ;
	    RECT 159.8000 106.1000 160.1000 107.9000 ;
	    RECT 160.6000 107.8000 162.6000 108.1000 ;
	    RECT 160.6000 106.1000 161.0000 106.2000 ;
	    RECT 158.2000 105.8000 159.0000 106.1000 ;
	    RECT 159.8000 105.8000 161.0000 106.1000 ;
	    RECT 155.0000 105.6000 157.1000 105.7000 ;
	    RECT 152.5000 105.2000 153.7000 105.5000 ;
	    RECT 146.2000 104.8000 146.6000 104.9000 ;
	    RECT 143.3000 101.1000 143.7000 104.7000 ;
	    RECT 146.3000 104.5000 146.6000 104.8000 ;
	    RECT 147.1000 104.5000 148.9000 104.6000 ;
	    RECT 145.4000 101.5000 145.8000 104.5000 ;
	    RECT 146.2000 101.7000 146.6000 104.5000 ;
	    RECT 147.0000 104.3000 148.9000 104.5000 ;
	    RECT 145.5000 101.4000 145.8000 101.5000 ;
	    RECT 147.0000 101.5000 147.4000 104.3000 ;
	    RECT 148.6000 104.1000 148.9000 104.3000 ;
	    RECT 149.5000 104.4000 151.3000 104.7000 ;
	    RECT 149.5000 104.1000 149.8000 104.4000 ;
	    RECT 147.0000 101.4000 147.3000 101.5000 ;
	    RECT 145.5000 101.1000 147.3000 101.4000 ;
	    RECT 147.8000 101.4000 148.2000 104.0000 ;
	    RECT 148.6000 101.7000 149.0000 104.1000 ;
	    RECT 149.4000 101.4000 149.8000 104.1000 ;
	    RECT 147.8000 101.1000 149.8000 101.4000 ;
	    RECT 151.0000 104.1000 151.3000 104.4000 ;
	    RECT 151.0000 101.1000 151.4000 104.1000 ;
	    RECT 151.8000 101.1000 152.2000 105.1000 ;
	    RECT 153.4000 103.1000 153.7000 105.2000 ;
	    RECT 155.0000 105.4000 157.0000 105.6000 ;
	    RECT 153.4000 101.1000 153.8000 103.1000 ;
	    RECT 155.0000 101.1000 155.4000 105.4000 ;
	    RECT 157.5000 105.1000 157.8000 105.8000 ;
	    RECT 158.6000 105.6000 159.0000 105.8000 ;
	    RECT 160.6000 105.1000 160.9000 105.8000 ;
	    RECT 157.1000 104.8000 157.8000 105.1000 ;
	    RECT 158.2000 104.8000 160.2000 105.1000 ;
	    RECT 157.1000 101.1000 157.5000 104.8000 ;
	    RECT 158.2000 101.1000 158.6000 104.8000 ;
	    RECT 159.8000 101.1000 160.2000 104.8000 ;
	    RECT 160.6000 101.1000 161.0000 105.1000 ;
	    RECT 163.0000 101.1000 163.4000 109.9000 ;
	    RECT 165.2000 109.2000 165.6000 109.9000 ;
	    RECT 165.2000 108.8000 165.8000 109.2000 ;
	    RECT 163.8000 107.8000 164.2000 108.6000 ;
	    RECT 165.2000 107.1000 165.6000 108.8000 ;
	    RECT 167.8000 107.9000 168.2000 109.9000 ;
	    RECT 169.9000 108.4000 170.3000 109.9000 ;
	    RECT 169.9000 107.9000 170.6000 108.4000 ;
	    RECT 167.9000 107.8000 168.2000 107.9000 ;
	    RECT 167.9000 107.6000 168.8000 107.8000 ;
	    RECT 167.9000 107.5000 170.0000 107.6000 ;
	    RECT 168.5000 107.3000 170.0000 107.5000 ;
	    RECT 169.6000 107.2000 170.0000 107.3000 ;
	    RECT 164.7000 106.9000 165.6000 107.1000 ;
	    RECT 164.7000 106.8000 165.5000 106.9000 ;
	    RECT 163.8000 105.8000 164.2000 106.2000 ;
	    RECT 163.8000 105.1000 164.1000 105.8000 ;
	    RECT 164.7000 105.2000 165.0000 106.8000 ;
	    RECT 167.8000 106.4000 168.2000 107.2000 ;
	    RECT 168.8000 106.9000 169.2000 107.0000 ;
	    RECT 168.7000 106.6000 169.2000 106.9000 ;
	    RECT 168.7000 106.2000 169.0000 106.6000 ;
	    RECT 165.8000 105.8000 166.6000 106.2000 ;
	    RECT 168.6000 105.8000 169.0000 106.2000 ;
	    RECT 164.6000 105.1000 165.0000 105.2000 ;
	    RECT 163.8000 104.8000 165.0000 105.1000 ;
	    RECT 167.0000 104.8000 167.4000 105.6000 ;
	    RECT 169.6000 105.5000 169.9000 107.2000 ;
	    RECT 170.3000 106.2000 170.6000 107.9000 ;
	    RECT 172.8000 107.1000 173.2000 109.9000 ;
	    RECT 172.8000 106.9000 173.7000 107.1000 ;
	    RECT 172.9000 106.8000 173.7000 106.9000 ;
	    RECT 174.2000 106.8000 174.6000 107.6000 ;
	    RECT 170.2000 105.8000 170.6000 106.2000 ;
	    RECT 171.8000 105.8000 172.6000 106.2000 ;
	    RECT 168.7000 105.2000 169.9000 105.5000 ;
	    RECT 164.7000 103.5000 165.0000 104.8000 ;
	    RECT 165.4000 103.8000 165.8000 104.6000 ;
	    RECT 164.7000 103.2000 166.5000 103.5000 ;
	    RECT 164.7000 103.1000 165.0000 103.2000 ;
	    RECT 164.6000 101.1000 165.0000 103.1000 ;
	    RECT 166.2000 103.1000 166.5000 103.2000 ;
	    RECT 168.7000 103.1000 169.0000 105.2000 ;
	    RECT 170.3000 105.1000 170.6000 105.8000 ;
	    RECT 166.2000 101.1000 166.6000 103.1000 ;
	    RECT 168.6000 101.1000 169.0000 103.1000 ;
	    RECT 170.2000 101.1000 170.6000 105.1000 ;
	    RECT 171.0000 104.8000 171.4000 105.6000 ;
	    RECT 173.4000 105.2000 173.7000 106.8000 ;
	    RECT 173.4000 104.8000 173.8000 105.2000 ;
	    RECT 172.6000 103.8000 173.0000 104.6000 ;
	    RECT 173.4000 103.5000 173.7000 104.8000 ;
	    RECT 171.9000 103.2000 173.7000 103.5000 ;
	    RECT 171.9000 103.1000 172.2000 103.2000 ;
	    RECT 171.8000 101.1000 172.2000 103.1000 ;
	    RECT 173.4000 103.1000 173.7000 103.2000 ;
	    RECT 173.4000 101.1000 173.8000 103.1000 ;
	    RECT 175.0000 101.1000 175.4000 109.9000 ;
	    RECT 176.4000 107.1000 176.8000 109.9000 ;
	    RECT 179.1000 108.2000 179.5000 108.6000 ;
	    RECT 179.0000 107.8000 179.4000 108.2000 ;
	    RECT 179.8000 107.9000 180.2000 109.9000 ;
	    RECT 182.2000 108.0000 182.6000 109.9000 ;
	    RECT 183.8000 108.0000 184.2000 109.9000 ;
	    RECT 182.2000 107.9000 184.2000 108.0000 ;
	    RECT 184.6000 107.9000 185.0000 109.9000 ;
	    RECT 185.4000 107.9000 185.8000 109.9000 ;
	    RECT 187.6000 108.1000 188.4000 109.9000 ;
	    RECT 175.9000 106.9000 176.8000 107.1000 ;
	    RECT 175.9000 106.8000 176.7000 106.9000 ;
	    RECT 175.9000 105.2000 176.2000 106.8000 ;
	    RECT 177.0000 105.8000 177.8000 106.2000 ;
	    RECT 179.0000 106.1000 179.4000 106.2000 ;
	    RECT 179.9000 106.1000 180.2000 107.9000 ;
	    RECT 182.3000 107.7000 184.1000 107.9000 ;
	    RECT 182.6000 107.2000 183.0000 107.4000 ;
	    RECT 184.6000 107.2000 184.9000 107.9000 ;
	    RECT 185.4000 107.6000 186.6000 107.9000 ;
	    RECT 186.2000 107.5000 186.6000 107.6000 ;
	    RECT 186.9000 107.4000 187.3000 107.8000 ;
	    RECT 186.9000 107.2000 187.2000 107.4000 ;
	    RECT 180.6000 106.4000 181.0000 107.2000 ;
	    RECT 182.2000 106.9000 183.0000 107.2000 ;
	    RECT 182.2000 106.8000 182.6000 106.9000 ;
	    RECT 183.7000 106.8000 185.0000 107.2000 ;
	    RECT 185.4000 106.8000 186.2000 107.2000 ;
	    RECT 186.8000 106.8000 187.2000 107.2000 ;
	    RECT 181.4000 106.1000 181.8000 106.2000 ;
	    RECT 179.0000 105.8000 180.2000 106.1000 ;
	    RECT 181.0000 105.8000 181.8000 106.1000 ;
	    RECT 183.0000 105.8000 183.4000 106.6000 ;
	    RECT 175.8000 104.8000 176.2000 105.2000 ;
	    RECT 178.2000 104.8000 178.6000 105.6000 ;
	    RECT 179.1000 105.1000 179.4000 105.8000 ;
	    RECT 181.0000 105.6000 181.4000 105.8000 ;
	    RECT 183.7000 105.2000 184.0000 106.8000 ;
	    RECT 185.4000 106.1000 185.7000 106.8000 ;
	    RECT 187.6000 106.4000 187.9000 108.1000 ;
	    RECT 190.2000 107.9000 190.6000 109.9000 ;
	    RECT 191.1000 108.2000 191.5000 108.6000 ;
	    RECT 188.2000 107.7000 189.0000 107.8000 ;
	    RECT 188.2000 107.4000 189.2000 107.7000 ;
	    RECT 189.5000 107.6000 190.6000 107.9000 ;
	    RECT 191.0000 107.8000 191.4000 108.2000 ;
	    RECT 191.8000 107.9000 192.2000 109.9000 ;
	    RECT 194.2000 108.0000 194.6000 109.9000 ;
	    RECT 195.8000 108.0000 196.2000 109.9000 ;
	    RECT 194.2000 107.9000 196.2000 108.0000 ;
	    RECT 196.6000 107.9000 197.0000 109.9000 ;
	    RECT 197.4000 107.9000 197.8000 109.9000 ;
	    RECT 199.6000 108.1000 200.4000 109.9000 ;
	    RECT 189.5000 107.5000 189.9000 107.6000 ;
	    RECT 188.9000 107.2000 189.2000 107.4000 ;
	    RECT 188.2000 106.7000 188.6000 107.1000 ;
	    RECT 188.9000 106.9000 190.6000 107.2000 ;
	    RECT 189.8000 106.8000 190.6000 106.9000 ;
	    RECT 187.4000 106.2000 187.9000 106.4000 ;
	    RECT 175.9000 103.5000 176.2000 104.8000 ;
	    RECT 176.6000 103.8000 177.0000 104.6000 ;
	    RECT 175.9000 103.2000 177.7000 103.5000 ;
	    RECT 175.9000 103.1000 176.2000 103.2000 ;
	    RECT 175.8000 101.1000 176.2000 103.1000 ;
	    RECT 177.4000 103.1000 177.7000 103.2000 ;
	    RECT 177.4000 101.1000 177.8000 103.1000 ;
	    RECT 179.0000 101.1000 179.4000 105.1000 ;
	    RECT 179.8000 104.8000 181.8000 105.1000 ;
	    RECT 183.0000 104.8000 184.0000 105.2000 ;
	    RECT 184.6000 105.8000 185.7000 106.1000 ;
	    RECT 187.0000 106.1000 187.9000 106.2000 ;
	    RECT 188.3000 106.4000 188.6000 106.7000 ;
	    RECT 188.3000 106.1000 189.6000 106.4000 ;
	    RECT 187.0000 105.8000 187.7000 106.1000 ;
	    RECT 189.2000 106.0000 189.6000 106.1000 ;
	    RECT 191.0000 106.1000 191.4000 106.2000 ;
	    RECT 191.9000 106.1000 192.2000 107.9000 ;
	    RECT 194.3000 107.7000 196.1000 107.9000 ;
	    RECT 194.6000 107.2000 195.0000 107.4000 ;
	    RECT 196.6000 107.2000 196.9000 107.9000 ;
	    RECT 197.4000 107.6000 198.6000 107.9000 ;
	    RECT 198.2000 107.5000 198.6000 107.6000 ;
	    RECT 198.9000 107.4000 199.3000 107.8000 ;
	    RECT 198.9000 107.2000 199.2000 107.4000 ;
	    RECT 192.6000 106.4000 193.0000 107.2000 ;
	    RECT 194.2000 106.9000 195.0000 107.2000 ;
	    RECT 194.2000 106.8000 194.6000 106.9000 ;
	    RECT 195.7000 106.8000 197.0000 107.2000 ;
	    RECT 197.4000 106.8000 198.2000 107.2000 ;
	    RECT 198.8000 106.8000 199.2000 107.2000 ;
	    RECT 193.4000 106.1000 193.8000 106.2000 ;
	    RECT 191.0000 105.8000 192.2000 106.1000 ;
	    RECT 193.0000 105.8000 193.8000 106.1000 ;
	    RECT 195.0000 105.8000 195.4000 106.6000 ;
	    RECT 184.6000 105.2000 184.9000 105.8000 ;
	    RECT 184.6000 105.1000 185.0000 105.2000 ;
	    RECT 187.4000 105.1000 187.7000 105.8000 ;
	    RECT 188.1000 105.7000 188.5000 105.8000 ;
	    RECT 188.1000 105.4000 189.8000 105.7000 ;
	    RECT 189.5000 105.1000 189.8000 105.4000 ;
	    RECT 191.1000 105.1000 191.4000 105.8000 ;
	    RECT 193.0000 105.6000 193.4000 105.8000 ;
	    RECT 195.7000 105.2000 196.0000 106.8000 ;
	    RECT 197.4000 106.1000 197.7000 106.8000 ;
	    RECT 199.6000 106.4000 199.9000 108.1000 ;
	    RECT 202.2000 107.9000 202.6000 109.9000 ;
	    RECT 204.3000 109.2000 204.7000 109.9000 ;
	    RECT 204.3000 108.8000 205.0000 109.2000 ;
	    RECT 204.3000 108.2000 204.7000 108.8000 ;
	    RECT 200.2000 107.7000 201.0000 107.8000 ;
	    RECT 200.2000 107.4000 201.2000 107.7000 ;
	    RECT 201.5000 107.6000 202.6000 107.9000 ;
	    RECT 203.8000 107.9000 204.7000 108.2000 ;
	    RECT 205.4000 108.0000 205.8000 109.9000 ;
	    RECT 207.0000 108.0000 207.4000 109.9000 ;
	    RECT 205.4000 107.9000 207.4000 108.0000 ;
	    RECT 207.8000 107.9000 208.2000 109.9000 ;
	    RECT 208.7000 108.2000 209.1000 108.6000 ;
	    RECT 201.5000 107.5000 201.9000 107.6000 ;
	    RECT 200.9000 107.2000 201.2000 107.4000 ;
	    RECT 200.2000 106.7000 200.6000 107.1000 ;
	    RECT 200.9000 106.9000 202.6000 107.2000 ;
	    RECT 201.8000 106.8000 202.6000 106.9000 ;
	    RECT 203.0000 106.8000 203.4000 107.6000 ;
	    RECT 199.4000 106.2000 199.9000 106.4000 ;
	    RECT 184.3000 104.8000 185.0000 105.1000 ;
	    RECT 185.4000 104.8000 186.6000 105.1000 ;
	    RECT 187.4000 104.8000 188.4000 105.1000 ;
	    RECT 179.8000 101.1000 180.2000 104.8000 ;
	    RECT 181.4000 101.1000 181.8000 104.8000 ;
	    RECT 183.5000 101.1000 183.9000 104.8000 ;
	    RECT 184.3000 104.2000 184.6000 104.8000 ;
	    RECT 184.2000 103.8000 184.6000 104.2000 ;
	    RECT 185.4000 101.1000 185.8000 104.8000 ;
	    RECT 186.2000 104.7000 186.6000 104.8000 ;
	    RECT 187.6000 104.2000 188.4000 104.8000 ;
	    RECT 189.5000 104.8000 190.6000 105.1000 ;
	    RECT 189.5000 104.7000 189.9000 104.8000 ;
	    RECT 187.6000 103.8000 189.0000 104.2000 ;
	    RECT 187.6000 101.1000 188.4000 103.8000 ;
	    RECT 190.2000 101.1000 190.6000 104.8000 ;
	    RECT 191.0000 101.1000 191.4000 105.1000 ;
	    RECT 191.8000 104.8000 193.8000 105.1000 ;
	    RECT 195.0000 104.8000 196.0000 105.2000 ;
	    RECT 196.6000 105.8000 197.7000 106.1000 ;
	    RECT 199.0000 106.1000 199.9000 106.2000 ;
	    RECT 200.3000 106.4000 200.6000 106.7000 ;
	    RECT 200.3000 106.1000 201.6000 106.4000 ;
	    RECT 199.0000 105.8000 199.7000 106.1000 ;
	    RECT 201.2000 106.0000 201.6000 106.1000 ;
	    RECT 196.6000 105.2000 196.9000 105.8000 ;
	    RECT 196.6000 105.1000 197.0000 105.2000 ;
	    RECT 199.4000 105.1000 199.7000 105.8000 ;
	    RECT 200.1000 105.7000 200.5000 105.8000 ;
	    RECT 200.1000 105.4000 201.8000 105.7000 ;
	    RECT 201.5000 105.1000 201.8000 105.4000 ;
	    RECT 196.3000 104.8000 197.0000 105.1000 ;
	    RECT 197.4000 104.8000 198.6000 105.1000 ;
	    RECT 199.4000 104.8000 200.4000 105.1000 ;
	    RECT 191.8000 101.1000 192.2000 104.8000 ;
	    RECT 193.4000 101.1000 193.8000 104.8000 ;
	    RECT 195.5000 101.1000 195.9000 104.8000 ;
	    RECT 196.3000 104.2000 196.6000 104.8000 ;
	    RECT 196.2000 103.8000 196.6000 104.2000 ;
	    RECT 197.4000 101.1000 197.8000 104.8000 ;
	    RECT 198.2000 104.7000 198.6000 104.8000 ;
	    RECT 199.6000 104.2000 200.4000 104.8000 ;
	    RECT 201.5000 104.8000 202.6000 105.1000 ;
	    RECT 201.5000 104.7000 201.9000 104.8000 ;
	    RECT 199.6000 103.8000 201.0000 104.2000 ;
	    RECT 199.6000 101.1000 200.4000 103.8000 ;
	    RECT 202.2000 101.1000 202.6000 104.8000 ;
	    RECT 203.8000 101.1000 204.2000 107.9000 ;
	    RECT 205.5000 107.7000 207.3000 107.9000 ;
	    RECT 205.8000 107.2000 206.2000 107.4000 ;
	    RECT 207.8000 107.2000 208.1000 107.9000 ;
	    RECT 208.6000 107.8000 209.0000 108.2000 ;
	    RECT 209.4000 107.9000 209.8000 109.9000 ;
	    RECT 213.4000 107.9000 213.8000 109.9000 ;
	    RECT 214.2000 108.0000 214.6000 109.9000 ;
	    RECT 215.8000 108.0000 216.2000 109.9000 ;
	    RECT 214.2000 107.9000 216.2000 108.0000 ;
	    RECT 216.6000 108.5000 217.0000 109.5000 ;
	    RECT 205.4000 106.9000 206.2000 107.2000 ;
	    RECT 205.4000 106.8000 205.8000 106.9000 ;
	    RECT 206.9000 106.8000 208.2000 107.2000 ;
	    RECT 206.2000 106.1000 206.6000 106.6000 ;
	    RECT 204.6000 105.8000 206.6000 106.1000 ;
	    RECT 204.6000 105.2000 204.9000 105.8000 ;
	    RECT 204.6000 104.4000 205.0000 105.2000 ;
	    RECT 206.9000 105.1000 207.2000 106.8000 ;
	    RECT 209.5000 106.2000 209.8000 107.9000 ;
	    RECT 213.5000 107.2000 213.8000 107.9000 ;
	    RECT 214.3000 107.7000 216.1000 107.9000 ;
	    RECT 216.6000 107.4000 216.9000 108.5000 ;
	    RECT 218.7000 108.2000 219.1000 109.5000 ;
	    RECT 218.2000 108.0000 219.1000 108.2000 ;
	    RECT 218.2000 107.8000 219.5000 108.0000 ;
	    RECT 218.7000 107.7000 219.5000 107.8000 ;
	    RECT 219.1000 107.5000 219.5000 107.7000 ;
	    RECT 215.4000 107.2000 215.8000 107.4000 ;
	    RECT 210.2000 106.4000 210.6000 107.2000 ;
	    RECT 213.4000 106.8000 214.7000 107.2000 ;
	    RECT 215.4000 106.9000 216.2000 107.2000 ;
	    RECT 216.6000 107.1000 218.7000 107.4000 ;
	    RECT 215.8000 106.8000 216.2000 106.9000 ;
	    RECT 218.2000 106.9000 218.7000 107.1000 ;
	    RECT 219.2000 107.2000 219.5000 107.5000 ;
	    RECT 208.6000 106.1000 209.0000 106.2000 ;
	    RECT 209.4000 106.1000 209.8000 106.2000 ;
	    RECT 211.0000 106.1000 211.4000 106.2000 ;
	    RECT 208.6000 105.8000 209.8000 106.1000 ;
	    RECT 210.6000 105.8000 211.4000 106.1000 ;
	    RECT 207.8000 105.1000 208.2000 105.2000 ;
	    RECT 208.7000 105.1000 209.0000 105.8000 ;
	    RECT 210.6000 105.6000 211.0000 105.8000 ;
	    RECT 211.8000 105.1000 212.2000 105.2000 ;
	    RECT 213.4000 105.1000 213.8000 105.2000 ;
	    RECT 214.4000 105.1000 214.7000 106.8000 ;
	    RECT 215.0000 105.8000 215.4000 106.6000 ;
	    RECT 216.6000 105.8000 217.0000 106.6000 ;
	    RECT 217.4000 105.8000 217.8000 106.6000 ;
	    RECT 218.2000 106.5000 218.9000 106.9000 ;
	    RECT 219.2000 106.8000 220.2000 107.2000 ;
	    RECT 218.2000 105.5000 218.5000 106.5000 ;
	    RECT 216.6000 105.2000 218.5000 105.5000 ;
	    RECT 206.7000 104.8000 207.2000 105.1000 ;
	    RECT 207.5000 104.8000 208.2000 105.1000 ;
	    RECT 206.7000 101.1000 207.1000 104.8000 ;
	    RECT 207.5000 104.2000 207.8000 104.8000 ;
	    RECT 207.4000 103.8000 207.8000 104.2000 ;
	    RECT 208.6000 101.1000 209.0000 105.1000 ;
	    RECT 209.4000 104.8000 211.4000 105.1000 ;
	    RECT 211.8000 104.8000 214.1000 105.1000 ;
	    RECT 214.4000 104.8000 214.9000 105.1000 ;
	    RECT 209.4000 101.1000 209.8000 104.8000 ;
	    RECT 211.0000 101.1000 211.4000 104.8000 ;
	    RECT 213.8000 104.2000 214.1000 104.8000 ;
	    RECT 213.8000 103.8000 214.2000 104.2000 ;
	    RECT 214.5000 101.1000 214.9000 104.8000 ;
	    RECT 216.6000 103.5000 216.9000 105.2000 ;
	    RECT 219.2000 104.9000 219.5000 106.8000 ;
	    RECT 219.8000 105.4000 220.2000 106.2000 ;
	    RECT 218.7000 104.6000 219.5000 104.9000 ;
	    RECT 216.6000 101.5000 217.0000 103.5000 ;
	    RECT 218.7000 101.1000 219.1000 104.6000 ;
	    RECT 221.4000 101.1000 221.8000 109.9000 ;
	    RECT 222.2000 107.8000 222.6000 108.6000 ;
	    RECT 223.0000 107.9000 223.4000 109.9000 ;
	    RECT 223.8000 108.0000 224.2000 109.9000 ;
	    RECT 225.4000 108.0000 225.8000 109.9000 ;
	    RECT 223.8000 107.9000 225.8000 108.0000 ;
	    RECT 226.2000 107.9000 226.6000 109.9000 ;
	    RECT 228.3000 109.2000 228.7000 109.9000 ;
	    RECT 228.3000 108.8000 229.0000 109.2000 ;
	    RECT 228.3000 108.4000 228.7000 108.8000 ;
	    RECT 228.3000 107.9000 229.0000 108.4000 ;
	    RECT 230.2000 108.2000 230.6000 109.9000 ;
	    RECT 223.1000 107.2000 223.4000 107.9000 ;
	    RECT 223.9000 107.7000 225.7000 107.9000 ;
	    RECT 226.3000 107.8000 226.6000 107.9000 ;
	    RECT 226.3000 107.6000 227.2000 107.8000 ;
	    RECT 226.3000 107.5000 228.4000 107.6000 ;
	    RECT 225.0000 107.2000 225.4000 107.4000 ;
	    RECT 226.9000 107.3000 228.4000 107.5000 ;
	    RECT 228.0000 107.2000 228.4000 107.3000 ;
	    RECT 223.0000 106.8000 224.3000 107.2000 ;
	    RECT 225.0000 106.9000 225.8000 107.2000 ;
	    RECT 225.4000 106.8000 225.8000 106.9000 ;
	    RECT 223.0000 105.1000 223.4000 105.2000 ;
	    RECT 224.0000 105.1000 224.3000 106.8000 ;
	    RECT 224.6000 106.1000 225.0000 106.6000 ;
	    RECT 226.2000 106.4000 226.6000 107.2000 ;
	    RECT 227.2000 106.9000 227.6000 107.0000 ;
	    RECT 227.1000 106.6000 227.6000 106.9000 ;
	    RECT 227.1000 106.2000 227.4000 106.6000 ;
	    RECT 225.4000 106.1000 225.8000 106.2000 ;
	    RECT 224.6000 105.8000 225.8000 106.1000 ;
	    RECT 227.0000 105.8000 227.4000 106.2000 ;
	    RECT 228.0000 105.5000 228.3000 107.2000 ;
	    RECT 228.7000 106.2000 229.0000 107.9000 ;
	    RECT 228.6000 105.8000 229.0000 106.2000 ;
	    RECT 227.1000 105.2000 228.3000 105.5000 ;
	    RECT 223.0000 104.8000 223.7000 105.1000 ;
	    RECT 224.0000 104.8000 224.5000 105.1000 ;
	    RECT 223.4000 104.2000 223.7000 104.8000 ;
	    RECT 223.4000 103.8000 223.8000 104.2000 ;
	    RECT 224.1000 101.1000 224.5000 104.8000 ;
	    RECT 227.1000 103.1000 227.4000 105.2000 ;
	    RECT 228.7000 105.1000 229.0000 105.8000 ;
	    RECT 227.0000 101.1000 227.4000 103.1000 ;
	    RECT 228.6000 101.1000 229.0000 105.1000 ;
	    RECT 230.1000 107.8000 230.6000 108.2000 ;
	    RECT 230.1000 107.2000 230.4000 107.8000 ;
	    RECT 231.8000 107.6000 232.2000 109.9000 ;
	    RECT 233.4000 108.9000 233.8000 109.9000 ;
	    RECT 235.8000 108.9000 236.2000 109.9000 ;
	    RECT 232.6000 107.8000 233.0000 108.6000 ;
	    RECT 230.9000 107.3000 232.2000 107.6000 ;
	    RECT 230.1000 106.8000 230.6000 107.2000 ;
	    RECT 230.1000 105.1000 230.4000 106.8000 ;
	    RECT 230.9000 106.5000 231.2000 107.3000 ;
	    RECT 233.5000 107.2000 233.8000 108.9000 ;
	    RECT 235.0000 107.8000 235.4000 108.6000 ;
	    RECT 235.9000 107.2000 236.2000 108.9000 ;
	    RECT 233.4000 106.8000 233.8000 107.2000 ;
	    RECT 235.8000 106.8000 236.2000 107.2000 ;
	    RECT 230.7000 106.1000 231.2000 106.5000 ;
	    RECT 230.9000 105.1000 231.2000 106.1000 ;
	    RECT 231.7000 106.2000 232.1000 106.6000 ;
	    RECT 231.7000 105.8000 232.2000 106.2000 ;
	    RECT 233.5000 105.2000 233.8000 106.8000 ;
	    RECT 234.2000 105.4000 234.6000 106.2000 ;
	    RECT 233.4000 105.1000 233.8000 105.2000 ;
	    RECT 235.9000 105.1000 236.2000 106.8000 ;
	    RECT 238.2000 108.9000 238.6000 109.9000 ;
	    RECT 238.2000 107.2000 238.5000 108.9000 ;
	    RECT 239.0000 107.8000 239.4000 108.6000 ;
	    RECT 239.8000 107.8000 240.2000 108.6000 ;
	    RECT 238.2000 107.1000 238.6000 107.2000 ;
	    RECT 239.8000 107.1000 240.1000 107.8000 ;
	    RECT 238.2000 106.8000 240.1000 107.1000 ;
	    RECT 236.6000 106.1000 237.0000 106.2000 ;
	    RECT 237.4000 106.1000 237.8000 106.2000 ;
	    RECT 236.6000 105.8000 237.8000 106.1000 ;
	    RECT 236.6000 105.4000 237.0000 105.8000 ;
	    RECT 237.4000 105.4000 237.8000 105.8000 ;
	    RECT 238.2000 105.1000 238.5000 106.8000 ;
	    RECT 230.1000 104.6000 230.6000 105.1000 ;
	    RECT 230.9000 104.8000 232.2000 105.1000 ;
	    RECT 230.2000 101.1000 230.6000 104.6000 ;
	    RECT 231.8000 101.1000 232.2000 104.8000 ;
	    RECT 233.4000 104.7000 234.3000 105.1000 ;
	    RECT 235.8000 104.7000 236.7000 105.1000 ;
	    RECT 233.9000 101.1000 234.3000 104.7000 ;
	    RECT 236.3000 102.2000 236.7000 104.7000 ;
	    RECT 235.8000 101.8000 236.7000 102.2000 ;
	    RECT 236.3000 101.1000 236.7000 101.8000 ;
	    RECT 237.7000 104.7000 238.6000 105.1000 ;
	    RECT 237.7000 101.1000 238.1000 104.7000 ;
	    RECT 240.6000 101.1000 241.0000 109.9000 ;
	    RECT 241.4000 107.9000 241.8000 109.9000 ;
	    RECT 243.6000 109.2000 244.4000 109.9000 ;
	    RECT 243.0000 108.8000 244.4000 109.2000 ;
	    RECT 243.6000 108.1000 244.4000 108.8000 ;
	    RECT 241.4000 107.6000 242.7000 107.9000 ;
	    RECT 242.3000 107.5000 242.7000 107.6000 ;
	    RECT 243.0000 107.4000 243.8000 107.8000 ;
	    RECT 241.4000 107.1000 242.2000 107.2000 ;
	    RECT 244.1000 107.1000 244.4000 108.1000 ;
	    RECT 246.2000 107.9000 246.6000 109.9000 ;
	    RECT 244.7000 107.4000 245.1000 107.8000 ;
	    RECT 245.4000 107.6000 246.6000 107.9000 ;
	    RECT 247.8000 108.9000 248.2000 109.9000 ;
	    RECT 245.4000 107.5000 245.8000 107.6000 ;
	    RECT 241.4000 107.0000 242.5000 107.1000 ;
	    RECT 241.4000 106.8000 243.6000 107.0000 ;
	    RECT 242.2000 106.7000 243.6000 106.8000 ;
	    RECT 243.2000 106.6000 243.6000 106.7000 ;
	    RECT 243.9000 106.8000 244.4000 107.1000 ;
	    RECT 244.8000 107.2000 245.1000 107.4000 ;
	    RECT 247.8000 107.2000 248.1000 108.9000 ;
	    RECT 248.6000 107.8000 249.0000 108.6000 ;
	    RECT 249.5000 108.2000 249.9000 108.6000 ;
	    RECT 249.4000 107.8000 249.8000 108.2000 ;
	    RECT 250.2000 107.9000 250.6000 109.9000 ;
	    RECT 252.6000 108.0000 253.0000 109.9000 ;
	    RECT 254.2000 108.0000 254.6000 109.9000 ;
	    RECT 252.6000 107.9000 254.6000 108.0000 ;
	    RECT 255.0000 107.9000 255.4000 109.9000 ;
	    RECT 255.8000 107.9000 256.2000 109.9000 ;
	    RECT 258.0000 108.1000 258.8000 109.9000 ;
	    RECT 244.8000 106.8000 245.2000 107.2000 ;
	    RECT 247.8000 107.1000 248.2000 107.2000 ;
	    RECT 249.4000 107.1000 249.7000 107.8000 ;
	    RECT 247.8000 106.8000 249.7000 107.1000 ;
	    RECT 243.9000 106.2000 244.2000 106.8000 ;
	    RECT 242.5000 106.1000 242.9000 106.2000 ;
	    RECT 242.5000 105.8000 243.3000 106.1000 ;
	    RECT 243.8000 105.8000 244.2000 106.2000 ;
	    RECT 242.9000 105.7000 243.3000 105.8000 ;
	    RECT 243.9000 105.1000 244.2000 105.8000 ;
	    RECT 247.0000 105.4000 247.4000 106.2000 ;
	    RECT 247.8000 105.2000 248.1000 106.8000 ;
	    RECT 249.4000 106.1000 249.8000 106.2000 ;
	    RECT 250.3000 106.1000 250.6000 107.9000 ;
	    RECT 252.7000 107.7000 254.5000 107.9000 ;
	    RECT 253.0000 107.2000 253.4000 107.4000 ;
	    RECT 255.0000 107.2000 255.3000 107.9000 ;
	    RECT 255.8000 107.6000 257.1000 107.9000 ;
	    RECT 256.7000 107.5000 257.1000 107.6000 ;
	    RECT 257.4000 107.4000 258.2000 107.8000 ;
	    RECT 251.0000 106.4000 251.4000 107.2000 ;
	    RECT 252.6000 106.9000 253.4000 107.2000 ;
	    RECT 252.6000 106.8000 253.0000 106.9000 ;
	    RECT 254.1000 106.8000 255.4000 107.2000 ;
	    RECT 258.5000 107.1000 258.8000 108.1000 ;
	    RECT 260.6000 107.9000 261.0000 109.9000 ;
	    RECT 261.4000 107.9000 261.8000 109.9000 ;
	    RECT 262.2000 108.0000 262.6000 109.9000 ;
	    RECT 263.8000 108.0000 264.2000 109.9000 ;
	    RECT 262.2000 107.9000 264.2000 108.0000 ;
	    RECT 264.6000 107.9000 265.0000 109.9000 ;
	    RECT 265.4000 108.0000 265.8000 109.9000 ;
	    RECT 267.0000 108.0000 267.4000 109.9000 ;
	    RECT 265.4000 107.9000 267.4000 108.0000 ;
	    RECT 259.1000 107.4000 259.5000 107.8000 ;
	    RECT 259.8000 107.6000 261.0000 107.9000 ;
	    RECT 259.8000 107.5000 260.2000 107.6000 ;
	    RECT 258.3000 106.8000 258.8000 107.1000 ;
	    RECT 259.2000 107.2000 259.5000 107.4000 ;
	    RECT 261.5000 107.2000 261.8000 107.9000 ;
	    RECT 262.3000 107.7000 264.1000 107.9000 ;
	    RECT 264.7000 107.2000 265.0000 107.9000 ;
	    RECT 265.5000 107.7000 267.3000 107.9000 ;
	    RECT 266.6000 107.2000 267.0000 107.4000 ;
	    RECT 259.2000 106.8000 259.6000 107.2000 ;
	    RECT 261.4000 106.8000 262.7000 107.2000 ;
	    RECT 264.6000 106.8000 265.9000 107.2000 ;
	    RECT 266.6000 107.1000 267.4000 107.2000 ;
	    RECT 267.8000 107.1000 268.2000 109.9000 ;
	    RECT 268.6000 107.8000 269.0000 108.6000 ;
	    RECT 266.6000 106.9000 268.2000 107.1000 ;
	    RECT 267.0000 106.8000 268.2000 106.9000 ;
	    RECT 251.8000 106.1000 252.2000 106.2000 ;
	    RECT 253.4000 106.1000 253.8000 106.6000 ;
	    RECT 249.4000 105.8000 250.6000 106.1000 ;
	    RECT 251.4000 105.8000 253.8000 106.1000 ;
	    RECT 254.1000 106.1000 254.4000 106.8000 ;
	    RECT 258.3000 106.2000 258.6000 106.8000 ;
	    RECT 255.0000 106.1000 255.4000 106.2000 ;
	    RECT 254.1000 105.8000 255.4000 106.1000 ;
	    RECT 256.9000 106.1000 257.3000 106.2000 ;
	    RECT 256.9000 105.8000 257.7000 106.1000 ;
	    RECT 258.2000 105.8000 258.6000 106.2000 ;
	    RECT 247.8000 105.1000 248.2000 105.2000 ;
	    RECT 249.5000 105.1000 249.8000 105.8000 ;
	    RECT 251.4000 105.6000 251.8000 105.8000 ;
	    RECT 254.1000 105.1000 254.4000 105.8000 ;
	    RECT 257.3000 105.7000 257.7000 105.8000 ;
	    RECT 255.0000 105.1000 255.4000 105.2000 ;
	    RECT 258.3000 105.1000 258.6000 105.8000 ;
	    RECT 261.4000 105.1000 261.8000 105.2000 ;
	    RECT 262.4000 105.1000 262.7000 106.8000 ;
	    RECT 263.0000 105.8000 263.4000 106.6000 ;
	    RECT 264.6000 105.1000 265.0000 105.2000 ;
	    RECT 265.6000 105.1000 265.9000 106.8000 ;
	    RECT 266.2000 105.8000 266.6000 106.6000 ;
	    RECT 241.4000 104.8000 242.7000 105.1000 ;
	    RECT 241.4000 101.1000 241.8000 104.8000 ;
	    RECT 242.3000 104.7000 242.7000 104.8000 ;
	    RECT 243.6000 101.1000 244.4000 105.1000 ;
	    RECT 245.4000 104.8000 246.6000 105.1000 ;
	    RECT 245.4000 104.7000 245.8000 104.8000 ;
	    RECT 246.2000 101.1000 246.6000 104.8000 ;
	    RECT 247.3000 104.7000 248.2000 105.1000 ;
	    RECT 247.3000 101.1000 247.7000 104.7000 ;
	    RECT 249.4000 101.1000 249.8000 105.1000 ;
	    RECT 250.2000 104.8000 252.2000 105.1000 ;
	    RECT 250.2000 101.1000 250.6000 104.8000 ;
	    RECT 251.8000 101.1000 252.2000 104.8000 ;
	    RECT 253.9000 104.8000 254.4000 105.1000 ;
	    RECT 254.7000 104.8000 255.4000 105.1000 ;
	    RECT 255.8000 104.8000 257.1000 105.1000 ;
	    RECT 253.9000 101.1000 254.3000 104.8000 ;
	    RECT 254.7000 104.2000 255.0000 104.8000 ;
	    RECT 254.6000 103.8000 255.0000 104.2000 ;
	    RECT 255.8000 101.1000 256.2000 104.8000 ;
	    RECT 256.7000 104.7000 257.1000 104.8000 ;
	    RECT 258.0000 102.2000 258.8000 105.1000 ;
	    RECT 259.8000 104.8000 261.0000 105.1000 ;
	    RECT 261.4000 104.8000 262.1000 105.1000 ;
	    RECT 262.4000 104.8000 262.9000 105.1000 ;
	    RECT 264.6000 104.8000 265.3000 105.1000 ;
	    RECT 265.6000 104.8000 266.1000 105.1000 ;
	    RECT 259.8000 104.7000 260.2000 104.8000 ;
	    RECT 257.4000 101.8000 258.8000 102.2000 ;
	    RECT 258.0000 101.1000 258.8000 101.8000 ;
	    RECT 260.6000 101.1000 261.0000 104.8000 ;
	    RECT 261.8000 104.2000 262.1000 104.8000 ;
	    RECT 261.8000 103.8000 262.2000 104.2000 ;
	    RECT 262.5000 101.1000 262.9000 104.8000 ;
	    RECT 265.0000 104.2000 265.3000 104.8000 ;
	    RECT 265.0000 103.8000 265.4000 104.2000 ;
	    RECT 265.7000 101.1000 266.1000 104.8000 ;
	    RECT 267.8000 101.1000 268.2000 106.8000 ;
	    RECT 0.6000 96.1000 1.0000 96.2000 ;
	    RECT 1.4000 96.1000 1.8000 99.9000 ;
	    RECT 0.6000 95.8000 1.8000 96.1000 ;
	    RECT 3.5000 95.9000 4.5000 99.9000 ;
	    RECT 1.4000 94.1000 1.8000 95.8000 ;
	    RECT 3.8000 94.2000 4.1000 95.9000 ;
	    RECT 7.0000 95.1000 7.4000 99.9000 ;
	    RECT 7.8000 99.6000 9.8000 99.9000 ;
	    RECT 7.8000 95.9000 8.2000 99.6000 ;
	    RECT 8.6000 95.9000 9.0000 99.3000 ;
	    RECT 9.4000 96.2000 9.8000 99.6000 ;
	    RECT 11.0000 96.2000 11.4000 99.9000 ;
	    RECT 9.4000 95.9000 11.4000 96.2000 ;
	    RECT 8.7000 95.6000 9.0000 95.9000 ;
	    RECT 11.8000 95.8000 12.2000 96.6000 ;
	    RECT 7.8000 95.1000 8.2000 95.6000 ;
	    RECT 8.7000 95.3000 9.7000 95.6000 ;
	    RECT 7.0000 94.8000 8.2000 95.1000 ;
	    RECT 9.4000 95.2000 9.7000 95.3000 ;
	    RECT 10.6000 95.2000 11.0000 95.4000 ;
	    RECT 9.4000 94.8000 9.8000 95.2000 ;
	    RECT 10.6000 94.9000 11.4000 95.2000 ;
	    RECT 11.0000 94.8000 11.4000 94.9000 ;
	    RECT 2.2000 94.1000 2.6000 94.2000 ;
	    RECT 3.8000 94.1000 4.2000 94.2000 ;
	    RECT 5.4000 94.1000 5.8000 94.6000 ;
	    RECT 7.0000 94.1000 7.4000 94.8000 ;
	    RECT 1.4000 93.8000 3.0000 94.1000 ;
	    RECT 3.8000 93.8000 5.0000 94.1000 ;
	    RECT 5.4000 93.8000 7.4000 94.1000 ;
	    RECT 1.4000 91.1000 1.8000 93.8000 ;
	    RECT 2.6000 93.6000 3.0000 93.8000 ;
	    RECT 2.3000 93.1000 4.1000 93.3000 ;
	    RECT 4.7000 93.1000 5.0000 93.8000 ;
	    RECT 2.2000 93.0000 4.2000 93.1000 ;
	    RECT 2.2000 91.1000 2.6000 93.0000 ;
	    RECT 3.8000 91.4000 4.2000 93.0000 ;
	    RECT 4.6000 91.7000 5.0000 93.1000 ;
	    RECT 5.4000 91.4000 5.8000 93.1000 ;
	    RECT 3.8000 91.1000 5.8000 91.4000 ;
	    RECT 7.0000 91.1000 7.4000 93.8000 ;
	    RECT 9.4000 93.1000 9.7000 94.8000 ;
	    RECT 12.6000 93.1000 13.0000 99.9000 ;
	    RECT 15.0000 97.9000 15.4000 99.9000 ;
	    RECT 15.1000 95.8000 15.4000 97.9000 ;
	    RECT 16.6000 95.9000 17.0000 99.9000 ;
	    RECT 17.4000 96.2000 17.8000 99.9000 ;
	    RECT 18.2000 96.2000 18.6000 96.3000 ;
	    RECT 17.4000 95.9000 18.6000 96.2000 ;
	    RECT 19.6000 95.9000 20.4000 99.9000 ;
	    RECT 21.3000 96.2000 21.7000 96.3000 ;
	    RECT 22.2000 96.2000 22.6000 99.9000 ;
	    RECT 24.3000 99.2000 24.7000 99.9000 ;
	    RECT 23.8000 98.8000 24.7000 99.2000 ;
	    RECT 21.3000 95.9000 22.6000 96.2000 ;
	    RECT 24.3000 96.2000 24.7000 98.8000 ;
	    RECT 25.0000 96.8000 25.4000 97.2000 ;
	    RECT 25.1000 96.2000 25.4000 96.8000 ;
	    RECT 24.3000 95.9000 24.8000 96.2000 ;
	    RECT 25.1000 95.9000 25.8000 96.2000 ;
	    RECT 15.1000 95.5000 16.3000 95.8000 ;
	    RECT 15.0000 94.8000 15.4000 95.2000 ;
	    RECT 13.4000 94.1000 13.8000 94.2000 ;
	    RECT 14.2000 94.1000 14.6000 94.6000 ;
	    RECT 15.1000 94.4000 15.4000 94.8000 ;
	    RECT 15.1000 94.1000 15.6000 94.4000 ;
	    RECT 13.4000 93.8000 14.6000 94.1000 ;
	    RECT 15.2000 94.0000 15.6000 94.1000 ;
	    RECT 16.0000 93.8000 16.3000 95.5000 ;
	    RECT 16.7000 95.2000 17.0000 95.9000 ;
	    RECT 16.6000 94.8000 17.0000 95.2000 ;
	    RECT 13.4000 93.4000 13.8000 93.8000 ;
	    RECT 16.0000 93.7000 16.4000 93.8000 ;
	    RECT 14.9000 93.5000 16.4000 93.7000 ;
	    RECT 14.3000 93.4000 16.4000 93.5000 ;
	    RECT 14.3000 93.2000 15.2000 93.4000 ;
	    RECT 14.3000 93.1000 14.6000 93.2000 ;
	    RECT 16.7000 93.1000 17.0000 94.8000 ;
	    RECT 19.8000 95.2000 20.1000 95.9000 ;
	    RECT 20.7000 95.2000 21.1000 95.3000 ;
	    RECT 19.8000 94.8000 20.2000 95.2000 ;
	    RECT 20.7000 94.9000 21.5000 95.2000 ;
	    RECT 21.1000 94.8000 21.5000 94.9000 ;
	    RECT 19.8000 94.2000 20.1000 94.8000 ;
	    RECT 23.8000 94.4000 24.2000 95.2000 ;
	    RECT 24.5000 94.2000 24.8000 95.9000 ;
	    RECT 25.4000 95.8000 25.8000 95.9000 ;
	    RECT 26.2000 95.8000 26.6000 96.6000 ;
	    RECT 18.8000 93.8000 19.2000 94.2000 ;
	    RECT 18.9000 93.6000 19.2000 93.8000 ;
	    RECT 19.6000 93.9000 20.1000 94.2000 ;
	    RECT 23.0000 94.1000 23.4000 94.2000 ;
	    RECT 18.2000 93.4000 18.6000 93.5000 ;
	    RECT 9.1000 91.1000 9.9000 93.1000 ;
	    RECT 12.1000 92.8000 13.0000 93.1000 ;
	    RECT 12.1000 91.1000 12.5000 92.8000 ;
	    RECT 14.2000 91.1000 14.6000 93.1000 ;
	    RECT 16.3000 92.6000 17.0000 93.1000 ;
	    RECT 17.4000 93.1000 18.6000 93.4000 ;
	    RECT 18.9000 93.2000 19.3000 93.6000 ;
	    RECT 16.3000 92.2000 16.7000 92.6000 ;
	    RECT 16.3000 91.8000 17.0000 92.2000 ;
	    RECT 16.3000 91.1000 16.7000 91.8000 ;
	    RECT 17.4000 91.1000 17.8000 93.1000 ;
	    RECT 19.6000 92.9000 19.9000 93.9000 ;
	    RECT 23.0000 93.8000 23.8000 94.1000 ;
	    RECT 24.5000 93.8000 25.8000 94.2000 ;
	    RECT 23.4000 93.6000 23.8000 93.8000 ;
	    RECT 20.2000 93.2000 21.0000 93.6000 ;
	    RECT 21.3000 93.4000 21.7000 93.5000 ;
	    RECT 21.3000 93.1000 22.6000 93.4000 ;
	    RECT 23.1000 93.1000 24.9000 93.3000 ;
	    RECT 25.4000 93.1000 25.7000 93.8000 ;
	    RECT 27.0000 93.1000 27.4000 99.9000 ;
	    RECT 28.6000 96.2000 29.0000 99.9000 ;
	    RECT 30.2000 96.2000 30.6000 99.9000 ;
	    RECT 28.6000 95.9000 30.6000 96.2000 ;
	    RECT 31.0000 95.9000 31.4000 99.9000 ;
	    RECT 33.1000 96.3000 33.5000 99.9000 ;
	    RECT 32.6000 95.9000 33.5000 96.3000 ;
	    RECT 29.0000 95.2000 29.4000 95.4000 ;
	    RECT 31.0000 95.2000 31.3000 95.9000 ;
	    RECT 28.6000 94.9000 29.4000 95.2000 ;
	    RECT 30.2000 94.9000 31.4000 95.2000 ;
	    RECT 28.6000 94.8000 29.0000 94.9000 ;
	    RECT 27.8000 94.1000 28.2000 94.2000 ;
	    RECT 29.4000 94.1000 29.8000 94.6000 ;
	    RECT 27.8000 93.8000 29.8000 94.1000 ;
	    RECT 27.8000 93.4000 28.2000 93.8000 ;
	    RECT 19.6000 92.2000 20.4000 92.9000 ;
	    RECT 19.6000 91.8000 21.0000 92.2000 ;
	    RECT 19.6000 91.1000 20.4000 91.8000 ;
	    RECT 22.2000 91.1000 22.6000 93.1000 ;
	    RECT 23.0000 93.0000 25.0000 93.1000 ;
	    RECT 23.0000 91.1000 23.4000 93.0000 ;
	    RECT 24.6000 91.1000 25.0000 93.0000 ;
	    RECT 25.4000 91.1000 25.8000 93.1000 ;
	    RECT 26.5000 92.8000 27.4000 93.1000 ;
	    RECT 30.2000 93.1000 30.5000 94.9000 ;
	    RECT 31.0000 94.8000 31.4000 94.9000 ;
	    RECT 32.7000 94.2000 33.0000 95.9000 ;
	    RECT 33.4000 95.1000 33.8000 95.6000 ;
	    RECT 34.2000 95.1000 34.6000 99.9000 ;
	    RECT 33.4000 94.8000 34.6000 95.1000 ;
	    RECT 32.6000 94.1000 33.0000 94.2000 ;
	    RECT 31.0000 93.8000 33.0000 94.1000 ;
	    RECT 31.0000 93.2000 31.3000 93.8000 ;
	    RECT 26.5000 92.2000 26.9000 92.8000 ;
	    RECT 26.5000 91.8000 27.4000 92.2000 ;
	    RECT 26.5000 91.1000 26.9000 91.8000 ;
	    RECT 30.2000 91.1000 30.6000 93.1000 ;
	    RECT 31.0000 92.8000 31.4000 93.2000 ;
	    RECT 30.9000 92.4000 31.3000 92.8000 ;
	    RECT 32.7000 92.1000 33.0000 93.8000 ;
	    RECT 32.6000 91.1000 33.0000 92.1000 ;
	    RECT 34.2000 91.1000 34.6000 94.8000 ;
	    RECT 35.8000 92.4000 36.2000 93.2000 ;
	    RECT 36.6000 91.1000 37.0000 99.9000 ;
	    RECT 37.4000 96.2000 37.8000 99.9000 ;
	    RECT 39.6000 97.2000 40.4000 99.9000 ;
	    RECT 39.6000 96.8000 41.0000 97.2000 ;
	    RECT 38.2000 96.2000 38.6000 96.3000 ;
	    RECT 39.6000 96.2000 40.4000 96.8000 ;
	    RECT 37.4000 95.9000 38.6000 96.2000 ;
	    RECT 39.4000 95.9000 40.4000 96.2000 ;
	    RECT 41.5000 96.2000 41.9000 96.3000 ;
	    RECT 42.2000 96.2000 42.6000 99.9000 ;
	    RECT 41.5000 95.9000 42.6000 96.2000 ;
	    RECT 43.3000 96.3000 43.7000 99.9000 ;
	    RECT 43.3000 95.9000 44.2000 96.3000 ;
	    RECT 39.4000 95.2000 39.7000 95.9000 ;
	    RECT 41.5000 95.6000 41.8000 95.9000 ;
	    RECT 40.1000 95.3000 41.8000 95.6000 ;
	    RECT 40.1000 95.2000 40.5000 95.3000 ;
	    RECT 39.0000 94.9000 39.7000 95.2000 ;
	    RECT 41.2000 94.9000 41.6000 95.0000 ;
	    RECT 39.0000 94.8000 39.9000 94.9000 ;
	    RECT 39.4000 94.6000 39.9000 94.8000 ;
	    RECT 37.4000 93.8000 38.2000 94.2000 ;
	    RECT 38.8000 93.8000 39.2000 94.2000 ;
	    RECT 38.9000 93.6000 39.2000 93.8000 ;
	    RECT 38.2000 93.4000 38.6000 93.5000 ;
	    RECT 37.4000 93.1000 38.6000 93.4000 ;
	    RECT 38.9000 93.2000 39.3000 93.6000 ;
	    RECT 37.4000 91.1000 37.8000 93.1000 ;
	    RECT 39.6000 92.9000 39.9000 94.6000 ;
	    RECT 40.3000 94.6000 41.6000 94.9000 ;
	    RECT 43.0000 94.8000 43.4000 95.6000 ;
	    RECT 40.3000 94.3000 40.6000 94.6000 ;
	    RECT 40.2000 93.9000 40.6000 94.3000 ;
	    RECT 43.8000 94.2000 44.1000 95.9000 ;
	    RECT 41.8000 94.1000 42.6000 94.2000 ;
	    RECT 40.9000 93.8000 42.6000 94.1000 ;
	    RECT 43.8000 93.8000 44.2000 94.2000 ;
	    RECT 40.9000 93.6000 41.2000 93.8000 ;
	    RECT 40.2000 93.3000 41.2000 93.6000 ;
	    RECT 41.5000 93.4000 41.9000 93.5000 ;
	    RECT 40.2000 93.2000 41.0000 93.3000 ;
	    RECT 41.5000 93.1000 42.6000 93.4000 ;
	    RECT 39.6000 91.1000 40.4000 92.9000 ;
	    RECT 42.2000 91.1000 42.6000 93.1000 ;
	    RECT 43.0000 93.1000 43.4000 93.2000 ;
	    RECT 43.8000 93.1000 44.1000 93.8000 ;
	    RECT 43.0000 92.8000 44.1000 93.1000 ;
	    RECT 43.8000 92.1000 44.1000 92.8000 ;
	    RECT 44.6000 92.4000 45.0000 93.2000 ;
	    RECT 43.8000 91.1000 44.2000 92.1000 ;
	    RECT 45.4000 91.1000 45.8000 99.9000 ;
	    RECT 47.0000 95.9000 47.4000 99.9000 ;
	    RECT 47.8000 96.2000 48.2000 99.9000 ;
	    RECT 49.4000 96.2000 49.8000 99.9000 ;
	    RECT 51.5000 96.3000 51.9000 99.9000 ;
	    RECT 47.8000 95.9000 49.8000 96.2000 ;
	    RECT 51.0000 95.9000 51.9000 96.3000 ;
	    RECT 53.0000 96.8000 53.4000 97.2000 ;
	    RECT 53.0000 96.2000 53.3000 96.8000 ;
	    RECT 53.7000 96.2000 54.1000 99.9000 ;
	    RECT 52.6000 95.9000 53.3000 96.2000 ;
	    RECT 53.6000 95.9000 54.1000 96.2000 ;
	    RECT 47.1000 95.2000 47.4000 95.9000 ;
	    RECT 49.0000 95.2000 49.4000 95.4000 ;
	    RECT 47.0000 94.9000 48.2000 95.2000 ;
	    RECT 49.0000 94.9000 49.8000 95.2000 ;
	    RECT 47.0000 94.8000 47.4000 94.9000 ;
	    RECT 46.2000 92.4000 46.6000 93.2000 ;
	    RECT 47.0000 92.8000 47.4000 93.2000 ;
	    RECT 47.9000 93.1000 48.2000 94.9000 ;
	    RECT 49.4000 94.8000 49.8000 94.9000 ;
	    RECT 50.2000 95.1000 50.6000 95.2000 ;
	    RECT 51.1000 95.1000 51.4000 95.9000 ;
	    RECT 52.6000 95.8000 53.0000 95.9000 ;
	    RECT 50.2000 94.8000 51.4000 95.1000 ;
	    RECT 51.8000 95.1000 52.2000 95.6000 ;
	    RECT 53.6000 95.1000 53.9000 95.9000 ;
	    RECT 51.8000 94.8000 53.9000 95.1000 ;
	    RECT 48.6000 93.8000 49.0000 94.6000 ;
	    RECT 51.1000 94.2000 51.4000 94.8000 ;
	    RECT 53.6000 94.2000 53.9000 94.8000 ;
	    RECT 54.2000 94.4000 54.6000 95.2000 ;
	    RECT 51.0000 93.8000 51.4000 94.2000 ;
	    RECT 52.6000 93.8000 53.9000 94.2000 ;
	    RECT 55.0000 94.1000 55.4000 94.2000 ;
	    RECT 56.6000 94.1000 57.0000 99.9000 ;
	    RECT 59.0000 95.9000 59.4000 99.9000 ;
	    RECT 59.8000 96.2000 60.2000 99.9000 ;
	    RECT 61.4000 96.2000 61.8000 99.9000 ;
	    RECT 59.8000 95.9000 61.8000 96.2000 ;
	    RECT 59.1000 95.2000 59.4000 95.9000 ;
	    RECT 62.2000 95.7000 62.6000 99.9000 ;
	    RECT 64.4000 98.2000 64.8000 99.9000 ;
	    RECT 63.8000 97.9000 64.8000 98.2000 ;
	    RECT 66.6000 97.9000 67.0000 99.9000 ;
	    RECT 68.7000 97.9000 69.3000 99.9000 ;
	    RECT 63.8000 97.5000 64.2000 97.9000 ;
	    RECT 66.6000 97.6000 66.9000 97.9000 ;
	    RECT 65.5000 97.3000 67.3000 97.6000 ;
	    RECT 68.6000 97.5000 69.0000 97.9000 ;
	    RECT 65.5000 97.2000 65.9000 97.3000 ;
	    RECT 66.9000 97.2000 67.3000 97.3000 ;
	    RECT 71.0000 97.1000 71.4000 99.9000 ;
	    RECT 72.6000 97.8000 73.0000 99.9000 ;
	    RECT 74.2000 97.9000 74.6000 99.9000 ;
	    RECT 74.2000 97.8000 74.5000 97.9000 ;
	    RECT 72.7000 97.5000 74.5000 97.8000 ;
	    RECT 63.8000 96.5000 64.2000 96.6000 ;
	    RECT 66.1000 96.5000 66.5000 96.6000 ;
	    RECT 63.8000 96.2000 66.5000 96.5000 ;
	    RECT 66.8000 96.5000 67.9000 96.8000 ;
	    RECT 66.8000 95.9000 67.1000 96.5000 ;
	    RECT 67.5000 96.4000 67.9000 96.5000 ;
	    RECT 68.7000 96.6000 69.4000 97.0000 ;
	    RECT 71.0000 96.8000 72.1000 97.1000 ;
	    RECT 68.7000 96.1000 69.0000 96.6000 ;
	    RECT 64.7000 95.7000 67.1000 95.9000 ;
	    RECT 62.2000 95.6000 67.1000 95.7000 ;
	    RECT 67.8000 95.8000 69.0000 96.1000 ;
	    RECT 62.2000 95.5000 65.1000 95.6000 ;
	    RECT 62.2000 95.4000 65.0000 95.5000 ;
	    RECT 61.0000 95.2000 61.4000 95.4000 ;
	    RECT 67.8000 95.2000 68.1000 95.8000 ;
	    RECT 71.0000 95.6000 71.4000 96.8000 ;
	    RECT 69.3000 95.3000 71.4000 95.6000 ;
	    RECT 71.8000 96.2000 72.1000 96.8000 ;
	    RECT 73.4000 96.4000 73.8000 97.2000 ;
	    RECT 74.2000 96.2000 74.5000 97.5000 ;
	    RECT 76.3000 96.3000 76.7000 99.9000 ;
	    RECT 71.8000 95.4000 72.2000 96.2000 ;
	    RECT 74.2000 95.8000 74.6000 96.2000 ;
	    RECT 75.8000 95.9000 76.7000 96.3000 ;
	    RECT 69.3000 95.2000 69.7000 95.3000 ;
	    RECT 59.0000 94.9000 60.2000 95.2000 ;
	    RECT 61.0000 94.9000 61.8000 95.2000 ;
	    RECT 65.4000 95.1000 65.8000 95.2000 ;
	    RECT 59.0000 94.8000 59.4000 94.9000 ;
	    RECT 54.6000 93.8000 57.0000 94.1000 ;
	    RECT 47.1000 92.4000 47.5000 92.8000 ;
	    RECT 47.8000 91.1000 48.2000 93.1000 ;
	    RECT 50.2000 92.4000 50.6000 93.2000 ;
	    RECT 51.1000 92.1000 51.4000 93.8000 ;
	    RECT 52.7000 93.1000 53.0000 93.8000 ;
	    RECT 54.6000 93.6000 55.0000 93.8000 ;
	    RECT 53.5000 93.1000 55.3000 93.3000 ;
	    RECT 51.0000 91.1000 51.4000 92.1000 ;
	    RECT 52.6000 91.1000 53.0000 93.1000 ;
	    RECT 53.4000 93.0000 55.4000 93.1000 ;
	    RECT 53.4000 91.1000 53.8000 93.0000 ;
	    RECT 55.0000 91.1000 55.4000 93.0000 ;
	    RECT 55.8000 92.4000 56.2000 93.2000 ;
	    RECT 56.6000 92.1000 57.0000 93.8000 ;
	    RECT 59.0000 92.8000 59.4000 93.2000 ;
	    RECT 59.9000 93.1000 60.2000 94.9000 ;
	    RECT 61.4000 94.8000 61.8000 94.9000 ;
	    RECT 63.3000 94.8000 65.8000 95.1000 ;
	    RECT 67.8000 94.8000 68.2000 95.2000 ;
	    RECT 70.1000 94.9000 70.5000 95.0000 ;
	    RECT 63.3000 94.7000 63.7000 94.8000 ;
	    RECT 64.6000 94.7000 65.0000 94.8000 ;
	    RECT 60.6000 93.8000 61.0000 94.6000 ;
	    RECT 64.1000 94.2000 64.5000 94.3000 ;
	    RECT 67.8000 94.2000 68.1000 94.8000 ;
	    RECT 68.6000 94.6000 70.5000 94.9000 ;
	    RECT 68.6000 94.5000 69.0000 94.6000 ;
	    RECT 62.6000 93.9000 68.1000 94.2000 ;
	    RECT 62.6000 93.8000 63.4000 93.9000 ;
	    RECT 59.1000 92.4000 59.5000 92.8000 ;
	    RECT 57.4000 92.1000 57.8000 92.2000 ;
	    RECT 56.6000 91.8000 57.8000 92.1000 ;
	    RECT 56.6000 91.1000 57.0000 91.8000 ;
	    RECT 59.8000 91.1000 60.2000 93.1000 ;
	    RECT 62.2000 91.1000 62.6000 93.5000 ;
	    RECT 64.7000 92.8000 65.0000 93.9000 ;
	    RECT 67.5000 93.8000 67.9000 93.9000 ;
	    RECT 71.0000 93.6000 71.4000 95.3000 ;
	    RECT 72.6000 94.8000 73.4000 95.2000 ;
	    RECT 74.2000 94.2000 74.5000 95.8000 ;
	    RECT 75.9000 94.2000 76.2000 95.9000 ;
	    RECT 77.4000 95.8000 77.8000 96.6000 ;
	    RECT 76.6000 95.1000 77.0000 95.6000 ;
	    RECT 78.2000 95.1000 78.6000 99.9000 ;
	    RECT 79.8000 97.9000 80.2000 99.9000 ;
	    RECT 79.9000 97.8000 80.2000 97.9000 ;
	    RECT 81.4000 97.9000 81.8000 99.9000 ;
	    RECT 83.0000 97.9000 83.4000 99.9000 ;
	    RECT 81.4000 97.8000 81.7000 97.9000 ;
	    RECT 79.9000 97.5000 81.7000 97.8000 ;
	    RECT 83.1000 97.8000 83.4000 97.9000 ;
	    RECT 84.6000 97.9000 85.0000 99.9000 ;
	    RECT 84.6000 97.8000 84.9000 97.9000 ;
	    RECT 83.1000 97.5000 84.9000 97.8000 ;
	    RECT 79.9000 96.2000 80.2000 97.5000 ;
	    RECT 80.6000 96.4000 81.0000 97.2000 ;
	    RECT 83.1000 96.2000 83.4000 97.5000 ;
	    RECT 83.8000 96.4000 84.2000 97.2000 ;
	    RECT 87.0000 96.4000 87.4000 99.9000 ;
	    RECT 79.8000 95.8000 80.2000 96.2000 ;
	    RECT 76.6000 94.8000 78.6000 95.1000 ;
	    RECT 73.7000 94.1000 74.5000 94.2000 ;
	    RECT 69.5000 93.3000 71.4000 93.6000 ;
	    RECT 69.5000 93.2000 69.9000 93.3000 ;
	    RECT 63.8000 92.1000 64.2000 92.5000 ;
	    RECT 64.6000 92.4000 65.0000 92.8000 ;
	    RECT 65.5000 92.7000 65.9000 92.8000 ;
	    RECT 65.5000 92.4000 66.9000 92.7000 ;
	    RECT 66.6000 92.1000 66.9000 92.4000 ;
	    RECT 68.6000 92.1000 69.0000 92.5000 ;
	    RECT 63.8000 91.8000 64.8000 92.1000 ;
	    RECT 64.4000 91.1000 64.8000 91.8000 ;
	    RECT 66.6000 91.1000 67.0000 92.1000 ;
	    RECT 68.6000 91.8000 69.3000 92.1000 ;
	    RECT 68.7000 91.1000 69.3000 91.8000 ;
	    RECT 71.0000 91.1000 71.4000 93.3000 ;
	    RECT 73.6000 93.9000 74.5000 94.1000 ;
	    RECT 73.6000 91.1000 74.0000 93.9000 ;
	    RECT 75.8000 93.8000 76.2000 94.2000 ;
	    RECT 75.0000 92.4000 75.4000 93.2000 ;
	    RECT 75.9000 92.2000 76.2000 93.8000 ;
	    RECT 78.2000 93.1000 78.6000 94.8000 ;
	    RECT 79.9000 94.2000 80.2000 95.8000 ;
	    RECT 81.0000 94.8000 81.8000 95.2000 ;
	    RECT 82.2000 94.8000 82.6000 96.2000 ;
	    RECT 83.0000 95.8000 83.4000 96.2000 ;
	    RECT 83.1000 94.2000 83.4000 95.8000 ;
	    RECT 84.2000 94.8000 85.0000 95.2000 ;
	    RECT 85.4000 95.1000 85.8000 96.2000 ;
	    RECT 86.9000 95.9000 87.4000 96.4000 ;
	    RECT 88.6000 96.2000 89.0000 99.9000 ;
	    RECT 90.2000 96.4000 90.6000 99.9000 ;
	    RECT 87.7000 95.9000 89.0000 96.2000 ;
	    RECT 90.1000 95.9000 90.6000 96.4000 ;
	    RECT 91.8000 96.2000 92.2000 99.9000 ;
	    RECT 93.4000 96.4000 93.8000 99.9000 ;
	    RECT 90.9000 95.9000 92.2000 96.2000 ;
	    RECT 93.3000 95.9000 93.8000 96.4000 ;
	    RECT 95.0000 96.2000 95.4000 99.9000 ;
	    RECT 96.2000 96.8000 96.6000 97.2000 ;
	    RECT 96.2000 96.2000 96.5000 96.8000 ;
	    RECT 96.9000 96.2000 97.3000 99.9000 ;
	    RECT 94.1000 95.9000 95.4000 96.2000 ;
	    RECT 95.8000 95.9000 96.5000 96.2000 ;
	    RECT 96.8000 95.9000 97.3000 96.2000 ;
	    RECT 99.0000 95.9000 99.4000 99.9000 ;
	    RECT 99.8000 96.2000 100.2000 99.9000 ;
	    RECT 101.4000 96.2000 101.8000 99.9000 ;
	    RECT 99.8000 95.9000 101.8000 96.2000 ;
	    RECT 86.2000 95.1000 86.6000 95.2000 ;
	    RECT 85.4000 94.8000 86.6000 95.1000 ;
	    RECT 86.9000 94.2000 87.2000 95.9000 ;
	    RECT 87.7000 94.9000 88.0000 95.9000 ;
	    RECT 87.5000 94.5000 88.0000 94.9000 ;
	    RECT 79.0000 93.4000 79.4000 94.2000 ;
	    RECT 79.9000 94.1000 80.7000 94.2000 ;
	    RECT 83.1000 94.1000 83.9000 94.2000 ;
	    RECT 79.9000 93.9000 80.8000 94.1000 ;
	    RECT 83.1000 93.9000 84.0000 94.1000 ;
	    RECT 75.8000 91.1000 76.2000 92.2000 ;
	    RECT 77.7000 92.8000 78.6000 93.1000 ;
	    RECT 77.7000 91.1000 78.1000 92.8000 ;
	    RECT 80.4000 91.1000 80.8000 93.9000 ;
	    RECT 83.6000 91.1000 84.0000 93.9000 ;
	    RECT 86.9000 93.8000 87.4000 94.2000 ;
	    RECT 86.9000 93.1000 87.2000 93.8000 ;
	    RECT 87.7000 93.7000 88.0000 94.5000 ;
	    RECT 88.5000 94.8000 89.0000 95.2000 ;
	    RECT 88.5000 94.4000 88.9000 94.8000 ;
	    RECT 90.1000 94.2000 90.4000 95.9000 ;
	    RECT 90.9000 94.9000 91.2000 95.9000 ;
	    RECT 90.7000 94.5000 91.2000 94.9000 ;
	    RECT 89.4000 94.1000 89.8000 94.2000 ;
	    RECT 90.1000 94.1000 90.6000 94.2000 ;
	    RECT 89.4000 93.8000 90.6000 94.1000 ;
	    RECT 87.7000 93.4000 89.0000 93.7000 ;
	    RECT 86.9000 92.8000 87.4000 93.1000 ;
	    RECT 87.0000 91.1000 87.4000 92.8000 ;
	    RECT 88.6000 91.1000 89.0000 93.4000 ;
	    RECT 90.1000 93.1000 90.4000 93.8000 ;
	    RECT 90.9000 93.7000 91.2000 94.5000 ;
	    RECT 91.7000 94.8000 92.2000 95.2000 ;
	    RECT 91.7000 94.4000 92.1000 94.8000 ;
	    RECT 93.3000 94.2000 93.6000 95.9000 ;
	    RECT 94.1000 94.9000 94.4000 95.9000 ;
	    RECT 95.8000 95.8000 96.2000 95.9000 ;
	    RECT 93.9000 94.5000 94.4000 94.9000 ;
	    RECT 93.3000 93.8000 93.8000 94.2000 ;
	    RECT 90.9000 93.4000 92.2000 93.7000 ;
	    RECT 90.1000 92.8000 90.6000 93.1000 ;
	    RECT 90.2000 91.1000 90.6000 92.8000 ;
	    RECT 91.8000 91.1000 92.2000 93.4000 ;
	    RECT 93.3000 93.2000 93.6000 93.8000 ;
	    RECT 94.1000 93.7000 94.4000 94.5000 ;
	    RECT 94.9000 94.8000 95.4000 95.2000 ;
	    RECT 94.9000 94.4000 95.3000 94.8000 ;
	    RECT 96.8000 94.2000 97.1000 95.9000 ;
	    RECT 99.1000 95.2000 99.4000 95.9000 ;
	    RECT 101.0000 95.2000 101.4000 95.4000 ;
	    RECT 97.4000 94.4000 97.8000 95.2000 ;
	    RECT 99.0000 94.9000 100.2000 95.2000 ;
	    RECT 101.0000 95.1000 101.8000 95.2000 ;
	    RECT 102.2000 95.1000 102.6000 99.9000 ;
	    RECT 103.8000 95.7000 104.2000 99.9000 ;
	    RECT 106.0000 98.2000 106.4000 99.9000 ;
	    RECT 105.4000 97.9000 106.4000 98.2000 ;
	    RECT 108.2000 97.9000 108.6000 99.9000 ;
	    RECT 110.3000 97.9000 110.9000 99.9000 ;
	    RECT 105.4000 97.5000 105.8000 97.9000 ;
	    RECT 108.2000 97.6000 108.5000 97.9000 ;
	    RECT 107.1000 97.3000 108.9000 97.6000 ;
	    RECT 110.2000 97.5000 110.6000 97.9000 ;
	    RECT 107.1000 97.2000 107.5000 97.3000 ;
	    RECT 108.5000 97.2000 108.9000 97.3000 ;
	    RECT 105.4000 96.5000 105.8000 96.6000 ;
	    RECT 107.7000 96.5000 108.1000 96.6000 ;
	    RECT 105.4000 96.2000 108.1000 96.5000 ;
	    RECT 108.4000 96.5000 109.5000 96.8000 ;
	    RECT 108.4000 95.9000 108.7000 96.5000 ;
	    RECT 109.1000 96.4000 109.5000 96.5000 ;
	    RECT 110.3000 96.6000 111.0000 97.0000 ;
	    RECT 110.3000 96.1000 110.6000 96.6000 ;
	    RECT 106.3000 95.7000 108.7000 95.9000 ;
	    RECT 103.8000 95.6000 108.7000 95.7000 ;
	    RECT 109.4000 95.8000 110.6000 96.1000 ;
	    RECT 103.8000 95.5000 106.7000 95.6000 ;
	    RECT 103.8000 95.4000 106.6000 95.5000 ;
	    RECT 109.4000 95.2000 109.7000 95.8000 ;
	    RECT 112.6000 95.6000 113.0000 99.9000 ;
	    RECT 110.9000 95.3000 113.0000 95.6000 ;
	    RECT 115.0000 95.7000 115.4000 99.9000 ;
	    RECT 117.2000 98.2000 117.6000 99.9000 ;
	    RECT 116.6000 97.9000 117.6000 98.2000 ;
	    RECT 119.4000 97.9000 119.8000 99.9000 ;
	    RECT 121.5000 97.9000 122.1000 99.9000 ;
	    RECT 116.6000 97.5000 117.0000 97.9000 ;
	    RECT 119.4000 97.6000 119.7000 97.9000 ;
	    RECT 118.3000 97.3000 120.1000 97.6000 ;
	    RECT 121.4000 97.5000 121.8000 97.9000 ;
	    RECT 118.3000 97.2000 118.7000 97.3000 ;
	    RECT 119.7000 97.2000 120.1000 97.3000 ;
	    RECT 116.6000 96.5000 117.0000 96.6000 ;
	    RECT 118.9000 96.5000 119.3000 96.6000 ;
	    RECT 116.6000 96.2000 119.3000 96.5000 ;
	    RECT 119.6000 96.5000 120.7000 96.8000 ;
	    RECT 119.6000 95.9000 119.9000 96.5000 ;
	    RECT 120.3000 96.4000 120.7000 96.5000 ;
	    RECT 121.5000 96.6000 122.2000 97.0000 ;
	    RECT 121.5000 96.1000 121.8000 96.6000 ;
	    RECT 117.5000 95.7000 119.9000 95.9000 ;
	    RECT 115.0000 95.6000 119.9000 95.7000 ;
	    RECT 120.6000 95.8000 121.8000 96.1000 ;
	    RECT 115.0000 95.5000 117.9000 95.6000 ;
	    RECT 115.0000 95.4000 117.8000 95.5000 ;
	    RECT 110.9000 95.2000 111.3000 95.3000 ;
	    RECT 107.0000 95.1000 107.4000 95.2000 ;
	    RECT 101.0000 94.9000 102.6000 95.1000 ;
	    RECT 99.0000 94.8000 99.4000 94.9000 ;
	    RECT 95.8000 93.8000 97.1000 94.2000 ;
	    RECT 98.2000 94.1000 98.6000 94.2000 ;
	    RECT 97.8000 93.8000 98.6000 94.1000 ;
	    RECT 99.0000 94.1000 99.4000 94.2000 ;
	    RECT 99.9000 94.1000 100.2000 94.9000 ;
	    RECT 101.4000 94.8000 102.6000 94.9000 ;
	    RECT 99.0000 93.8000 100.2000 94.1000 ;
	    RECT 100.6000 93.8000 101.0000 94.6000 ;
	    RECT 101.4000 94.2000 101.7000 94.8000 ;
	    RECT 101.4000 93.8000 101.8000 94.2000 ;
	    RECT 94.1000 93.4000 95.4000 93.7000 ;
	    RECT 93.3000 92.8000 93.8000 93.2000 ;
	    RECT 93.4000 91.1000 93.8000 92.8000 ;
	    RECT 95.0000 91.1000 95.4000 93.4000 ;
	    RECT 95.9000 93.1000 96.2000 93.8000 ;
	    RECT 97.8000 93.6000 98.2000 93.8000 ;
	    RECT 96.7000 93.1000 98.5000 93.3000 ;
	    RECT 95.8000 91.1000 96.2000 93.1000 ;
	    RECT 96.6000 93.0000 98.6000 93.1000 ;
	    RECT 96.6000 91.1000 97.0000 93.0000 ;
	    RECT 98.2000 91.1000 98.6000 93.0000 ;
	    RECT 99.0000 92.8000 99.4000 93.2000 ;
	    RECT 99.9000 93.1000 100.2000 93.8000 ;
	    RECT 99.1000 92.4000 99.5000 92.8000 ;
	    RECT 99.8000 91.1000 100.2000 93.1000 ;
	    RECT 102.2000 91.1000 102.6000 94.8000 ;
	    RECT 104.9000 94.8000 107.4000 95.1000 ;
	    RECT 109.4000 94.8000 109.8000 95.2000 ;
	    RECT 111.7000 94.9000 112.1000 95.0000 ;
	    RECT 104.9000 94.7000 105.3000 94.8000 ;
	    RECT 106.2000 94.7000 106.6000 94.8000 ;
	    RECT 105.7000 94.2000 106.1000 94.3000 ;
	    RECT 109.4000 94.2000 109.7000 94.8000 ;
	    RECT 110.2000 94.6000 112.1000 94.9000 ;
	    RECT 110.2000 94.5000 110.6000 94.6000 ;
	    RECT 104.2000 93.9000 109.7000 94.2000 ;
	    RECT 104.2000 93.8000 105.0000 93.9000 ;
	    RECT 103.0000 92.4000 103.4000 93.2000 ;
	    RECT 103.8000 91.1000 104.2000 93.5000 ;
	    RECT 106.3000 92.8000 106.6000 93.9000 ;
	    RECT 109.1000 93.8000 109.5000 93.9000 ;
	    RECT 112.6000 93.6000 113.0000 95.3000 ;
	    RECT 120.6000 95.2000 120.9000 95.8000 ;
	    RECT 122.2000 95.6000 122.6000 96.2000 ;
	    RECT 123.8000 95.6000 124.2000 99.9000 ;
	    RECT 122.1000 95.3000 124.2000 95.6000 ;
	    RECT 122.1000 95.2000 122.5000 95.3000 ;
	    RECT 118.2000 95.1000 118.6000 95.2000 ;
	    RECT 116.1000 94.8000 118.6000 95.1000 ;
	    RECT 120.6000 94.8000 121.0000 95.2000 ;
	    RECT 122.9000 94.9000 123.3000 95.0000 ;
	    RECT 116.1000 94.7000 116.5000 94.8000 ;
	    RECT 117.4000 94.7000 117.8000 94.8000 ;
	    RECT 116.9000 94.2000 117.3000 94.3000 ;
	    RECT 120.6000 94.2000 120.9000 94.8000 ;
	    RECT 121.4000 94.6000 123.3000 94.9000 ;
	    RECT 121.4000 94.5000 121.8000 94.6000 ;
	    RECT 114.2000 94.1000 114.6000 94.2000 ;
	    RECT 115.4000 94.1000 120.9000 94.2000 ;
	    RECT 114.2000 93.9000 120.9000 94.1000 ;
	    RECT 114.2000 93.8000 116.2000 93.9000 ;
	    RECT 111.1000 93.3000 113.0000 93.6000 ;
	    RECT 111.1000 93.2000 111.5000 93.3000 ;
	    RECT 105.4000 92.1000 105.8000 92.5000 ;
	    RECT 106.2000 92.4000 106.6000 92.8000 ;
	    RECT 107.1000 92.7000 107.5000 92.8000 ;
	    RECT 107.1000 92.4000 108.5000 92.7000 ;
	    RECT 108.2000 92.1000 108.5000 92.4000 ;
	    RECT 110.2000 92.1000 110.6000 92.5000 ;
	    RECT 112.6000 92.1000 113.0000 93.3000 ;
	    RECT 113.4000 92.1000 113.8000 92.2000 ;
	    RECT 105.4000 91.8000 106.4000 92.1000 ;
	    RECT 106.0000 91.1000 106.4000 91.8000 ;
	    RECT 108.2000 91.1000 108.6000 92.1000 ;
	    RECT 110.2000 91.8000 110.9000 92.1000 ;
	    RECT 110.3000 91.1000 110.9000 91.8000 ;
	    RECT 112.6000 91.8000 113.8000 92.1000 ;
	    RECT 112.6000 91.1000 113.0000 91.8000 ;
	    RECT 115.0000 91.1000 115.4000 93.5000 ;
	    RECT 117.5000 92.8000 117.8000 93.9000 ;
	    RECT 120.3000 93.8000 120.7000 93.9000 ;
	    RECT 123.8000 93.6000 124.2000 95.3000 ;
	    RECT 122.3000 93.3000 124.2000 93.6000 ;
	    RECT 122.3000 93.2000 122.7000 93.3000 ;
	    RECT 116.6000 92.1000 117.0000 92.5000 ;
	    RECT 117.4000 92.4000 117.8000 92.8000 ;
	    RECT 118.3000 92.7000 118.7000 92.8000 ;
	    RECT 118.3000 92.4000 119.7000 92.7000 ;
	    RECT 119.4000 92.1000 119.7000 92.4000 ;
	    RECT 121.4000 92.1000 121.8000 92.5000 ;
	    RECT 116.6000 91.8000 117.6000 92.1000 ;
	    RECT 117.2000 91.1000 117.6000 91.8000 ;
	    RECT 119.4000 91.1000 119.8000 92.1000 ;
	    RECT 121.4000 91.8000 122.1000 92.1000 ;
	    RECT 121.5000 91.1000 122.1000 91.8000 ;
	    RECT 123.8000 91.1000 124.2000 93.3000 ;
	    RECT 124.6000 91.1000 125.0000 99.9000 ;
	    RECT 125.4000 94.1000 125.8000 94.2000 ;
	    RECT 125.4000 93.8000 126.5000 94.1000 ;
	    RECT 125.4000 93.4000 125.8000 93.8000 ;
	    RECT 126.2000 93.2000 126.5000 93.8000 ;
	    RECT 126.2000 92.4000 126.6000 93.2000 ;
	    RECT 127.0000 91.1000 127.4000 99.9000 ;
	    RECT 127.8000 95.6000 128.2000 99.9000 ;
	    RECT 129.9000 97.9000 130.5000 99.9000 ;
	    RECT 132.2000 97.9000 132.6000 99.9000 ;
	    RECT 134.4000 98.2000 134.8000 99.9000 ;
	    RECT 134.4000 97.9000 135.4000 98.2000 ;
	    RECT 130.2000 97.5000 130.6000 97.9000 ;
	    RECT 132.3000 97.6000 132.6000 97.9000 ;
	    RECT 131.9000 97.3000 133.7000 97.6000 ;
	    RECT 135.0000 97.5000 135.4000 97.9000 ;
	    RECT 131.9000 97.2000 132.3000 97.3000 ;
	    RECT 133.3000 97.2000 133.7000 97.3000 ;
	    RECT 129.4000 97.0000 130.1000 97.2000 ;
	    RECT 129.4000 96.8000 130.5000 97.0000 ;
	    RECT 129.8000 96.6000 130.5000 96.8000 ;
	    RECT 130.2000 96.1000 130.5000 96.6000 ;
	    RECT 131.3000 96.5000 132.4000 96.8000 ;
	    RECT 131.3000 96.4000 131.7000 96.5000 ;
	    RECT 130.2000 95.8000 131.4000 96.1000 ;
	    RECT 127.8000 95.3000 129.9000 95.6000 ;
	    RECT 127.8000 93.6000 128.2000 95.3000 ;
	    RECT 129.5000 95.2000 129.9000 95.3000 ;
	    RECT 128.7000 94.9000 129.1000 95.0000 ;
	    RECT 128.7000 94.6000 130.6000 94.9000 ;
	    RECT 130.2000 94.5000 130.6000 94.6000 ;
	    RECT 131.1000 94.2000 131.4000 95.8000 ;
	    RECT 132.1000 95.9000 132.4000 96.5000 ;
	    RECT 132.7000 96.5000 133.1000 96.6000 ;
	    RECT 135.0000 96.5000 135.4000 96.6000 ;
	    RECT 132.7000 96.2000 135.4000 96.5000 ;
	    RECT 132.1000 95.7000 134.5000 95.9000 ;
	    RECT 136.6000 95.7000 137.0000 99.9000 ;
	    RECT 137.4000 96.2000 137.8000 99.9000 ;
	    RECT 139.0000 96.2000 139.4000 99.9000 ;
	    RECT 137.4000 95.9000 139.4000 96.2000 ;
	    RECT 139.8000 95.9000 140.2000 99.9000 ;
	    RECT 141.0000 96.8000 141.4000 97.2000 ;
	    RECT 141.0000 96.2000 141.3000 96.8000 ;
	    RECT 141.7000 96.2000 142.1000 99.9000 ;
	    RECT 145.1000 99.2000 145.5000 99.9000 ;
	    RECT 144.6000 98.8000 145.5000 99.2000 ;
	    RECT 140.6000 95.9000 141.3000 96.2000 ;
	    RECT 141.6000 95.9000 142.1000 96.2000 ;
	    RECT 145.1000 96.2000 145.5000 98.8000 ;
	    RECT 145.8000 96.8000 146.2000 97.2000 ;
	    RECT 145.9000 96.2000 146.2000 96.8000 ;
	    RECT 145.1000 95.9000 145.6000 96.2000 ;
	    RECT 145.9000 95.9000 146.6000 96.2000 ;
	    RECT 132.1000 95.6000 137.0000 95.7000 ;
	    RECT 134.1000 95.5000 137.0000 95.6000 ;
	    RECT 134.2000 95.4000 137.0000 95.5000 ;
	    RECT 137.8000 95.2000 138.2000 95.4000 ;
	    RECT 139.8000 95.2000 140.1000 95.9000 ;
	    RECT 140.6000 95.8000 141.0000 95.9000 ;
	    RECT 133.4000 95.1000 133.8000 95.2000 ;
	    RECT 133.4000 94.8000 135.9000 95.1000 ;
	    RECT 137.4000 94.9000 138.2000 95.2000 ;
	    RECT 139.0000 94.9000 140.2000 95.2000 ;
	    RECT 137.4000 94.8000 137.8000 94.9000 ;
	    RECT 134.2000 94.7000 134.6000 94.8000 ;
	    RECT 135.5000 94.7000 135.9000 94.8000 ;
	    RECT 134.7000 94.2000 135.1000 94.3000 ;
	    RECT 131.1000 93.9000 136.6000 94.2000 ;
	    RECT 131.3000 93.8000 131.7000 93.9000 ;
	    RECT 127.8000 93.3000 129.7000 93.6000 ;
	    RECT 127.8000 91.1000 128.2000 93.3000 ;
	    RECT 129.3000 93.2000 129.7000 93.3000 ;
	    RECT 134.2000 92.8000 134.5000 93.9000 ;
	    RECT 135.8000 93.8000 136.6000 93.9000 ;
	    RECT 138.2000 93.8000 138.6000 94.6000 ;
	    RECT 133.3000 92.7000 133.7000 92.8000 ;
	    RECT 130.2000 92.1000 130.6000 92.5000 ;
	    RECT 132.3000 92.4000 133.7000 92.7000 ;
	    RECT 134.2000 92.4000 134.6000 92.8000 ;
	    RECT 132.3000 92.1000 132.6000 92.4000 ;
	    RECT 135.0000 92.1000 135.4000 92.5000 ;
	    RECT 129.9000 91.8000 130.6000 92.1000 ;
	    RECT 129.9000 91.1000 130.5000 91.8000 ;
	    RECT 132.2000 91.1000 132.6000 92.1000 ;
	    RECT 134.4000 91.8000 135.4000 92.1000 ;
	    RECT 134.4000 91.1000 134.8000 91.8000 ;
	    RECT 136.6000 91.1000 137.0000 93.5000 ;
	    RECT 139.0000 93.1000 139.3000 94.9000 ;
	    RECT 139.8000 94.8000 140.2000 94.9000 ;
	    RECT 141.6000 94.2000 141.9000 95.9000 ;
	    RECT 142.2000 94.4000 142.6000 95.2000 ;
	    RECT 145.3000 94.2000 145.6000 95.9000 ;
	    RECT 146.2000 95.8000 146.6000 95.9000 ;
	    RECT 147.8000 95.6000 148.2000 99.9000 ;
	    RECT 149.4000 95.6000 149.8000 99.9000 ;
	    RECT 151.0000 95.6000 151.4000 99.9000 ;
	    RECT 152.6000 95.6000 153.0000 99.9000 ;
	    RECT 154.2000 95.7000 154.6000 99.9000 ;
	    RECT 156.4000 98.2000 156.8000 99.9000 ;
	    RECT 155.8000 97.9000 156.8000 98.2000 ;
	    RECT 158.6000 97.9000 159.0000 99.9000 ;
	    RECT 160.7000 97.9000 161.3000 99.9000 ;
	    RECT 155.8000 97.5000 156.2000 97.9000 ;
	    RECT 158.6000 97.6000 158.9000 97.9000 ;
	    RECT 157.5000 97.3000 159.3000 97.6000 ;
	    RECT 160.6000 97.5000 161.0000 97.9000 ;
	    RECT 157.5000 97.2000 157.9000 97.3000 ;
	    RECT 158.9000 97.2000 159.3000 97.3000 ;
	    RECT 161.1000 97.0000 161.8000 97.2000 ;
	    RECT 160.7000 96.8000 161.8000 97.0000 ;
	    RECT 155.8000 96.5000 156.2000 96.6000 ;
	    RECT 158.1000 96.5000 158.5000 96.6000 ;
	    RECT 155.8000 96.2000 158.5000 96.5000 ;
	    RECT 158.8000 96.5000 159.9000 96.8000 ;
	    RECT 158.8000 95.9000 159.1000 96.5000 ;
	    RECT 159.5000 96.4000 159.9000 96.5000 ;
	    RECT 160.7000 96.6000 161.4000 96.8000 ;
	    RECT 160.7000 96.1000 161.0000 96.6000 ;
	    RECT 156.7000 95.7000 159.1000 95.9000 ;
	    RECT 154.2000 95.6000 159.1000 95.7000 ;
	    RECT 159.8000 95.8000 161.0000 96.1000 ;
	    RECT 147.8000 95.2000 148.7000 95.6000 ;
	    RECT 149.4000 95.2000 150.5000 95.6000 ;
	    RECT 151.0000 95.2000 152.1000 95.6000 ;
	    RECT 152.6000 95.2000 153.8000 95.6000 ;
	    RECT 154.2000 95.5000 157.1000 95.6000 ;
	    RECT 154.2000 95.4000 157.0000 95.5000 ;
	    RECT 148.3000 94.5000 148.7000 95.2000 ;
	    RECT 150.1000 94.5000 150.5000 95.2000 ;
	    RECT 151.7000 94.5000 152.1000 95.2000 ;
	    RECT 140.6000 93.8000 141.9000 94.2000 ;
	    RECT 143.8000 94.1000 144.2000 94.2000 ;
	    RECT 143.8000 93.8000 144.6000 94.1000 ;
	    RECT 145.3000 93.8000 146.6000 94.2000 ;
	    RECT 148.3000 94.1000 149.6000 94.5000 ;
	    RECT 150.1000 94.1000 151.3000 94.5000 ;
	    RECT 151.7000 94.1000 153.0000 94.5000 ;
	    RECT 148.3000 93.8000 148.7000 94.1000 ;
	    RECT 150.1000 93.8000 150.5000 94.1000 ;
	    RECT 151.7000 93.8000 152.1000 94.1000 ;
	    RECT 153.4000 93.8000 153.8000 95.2000 ;
	    RECT 157.4000 95.1000 157.8000 95.2000 ;
	    RECT 155.3000 94.8000 157.8000 95.1000 ;
	    RECT 155.3000 94.7000 155.7000 94.8000 ;
	    RECT 156.1000 94.2000 156.5000 94.3000 ;
	    RECT 159.8000 94.2000 160.1000 95.8000 ;
	    RECT 163.0000 95.6000 163.4000 99.9000 ;
	    RECT 165.4000 95.9000 165.8000 99.9000 ;
	    RECT 166.2000 96.2000 166.6000 99.9000 ;
	    RECT 167.8000 96.2000 168.2000 99.9000 ;
	    RECT 166.2000 95.9000 168.2000 96.2000 ;
	    RECT 161.3000 95.3000 163.4000 95.6000 ;
	    RECT 161.3000 95.2000 161.7000 95.3000 ;
	    RECT 162.1000 94.9000 162.5000 95.0000 ;
	    RECT 160.6000 94.6000 162.5000 94.9000 ;
	    RECT 160.6000 94.5000 161.0000 94.6000 ;
	    RECT 154.6000 93.9000 160.1000 94.2000 ;
	    RECT 154.6000 93.8000 155.4000 93.9000 ;
	    RECT 139.8000 93.1000 140.2000 93.2000 ;
	    RECT 140.7000 93.1000 141.0000 93.8000 ;
	    RECT 144.2000 93.6000 144.6000 93.8000 ;
	    RECT 141.5000 93.1000 143.3000 93.3000 ;
	    RECT 143.9000 93.1000 145.7000 93.3000 ;
	    RECT 146.2000 93.1000 146.5000 93.8000 ;
	    RECT 147.8000 93.4000 148.7000 93.8000 ;
	    RECT 149.4000 93.4000 150.5000 93.8000 ;
	    RECT 151.0000 93.4000 152.1000 93.8000 ;
	    RECT 152.6000 93.4000 153.8000 93.8000 ;
	    RECT 139.0000 91.1000 139.4000 93.1000 ;
	    RECT 139.8000 92.8000 141.0000 93.1000 ;
	    RECT 139.7000 92.4000 140.1000 92.8000 ;
	    RECT 140.6000 91.1000 141.0000 92.8000 ;
	    RECT 141.4000 93.0000 143.4000 93.1000 ;
	    RECT 141.4000 91.1000 141.8000 93.0000 ;
	    RECT 143.0000 91.1000 143.4000 93.0000 ;
	    RECT 143.8000 93.0000 145.8000 93.1000 ;
	    RECT 143.8000 91.1000 144.2000 93.0000 ;
	    RECT 145.4000 91.1000 145.8000 93.0000 ;
	    RECT 146.2000 91.1000 146.6000 93.1000 ;
	    RECT 147.8000 91.1000 148.2000 93.4000 ;
	    RECT 149.4000 91.1000 149.8000 93.4000 ;
	    RECT 151.0000 91.1000 151.4000 93.4000 ;
	    RECT 152.6000 91.1000 153.0000 93.4000 ;
	    RECT 154.2000 91.1000 154.6000 93.5000 ;
	    RECT 156.7000 92.8000 157.0000 93.9000 ;
	    RECT 159.5000 93.8000 159.9000 93.9000 ;
	    RECT 163.0000 93.6000 163.4000 95.3000 ;
	    RECT 165.5000 95.2000 165.8000 95.9000 ;
	    RECT 168.6000 95.8000 169.0000 96.6000 ;
	    RECT 167.4000 95.2000 167.8000 95.4000 ;
	    RECT 164.6000 95.1000 165.0000 95.2000 ;
	    RECT 165.4000 95.1000 166.6000 95.2000 ;
	    RECT 164.6000 94.9000 166.6000 95.1000 ;
	    RECT 167.4000 94.9000 168.2000 95.2000 ;
	    RECT 164.6000 94.8000 165.8000 94.9000 ;
	    RECT 161.5000 93.3000 163.4000 93.6000 ;
	    RECT 161.5000 93.2000 161.9000 93.3000 ;
	    RECT 155.8000 92.1000 156.2000 92.5000 ;
	    RECT 156.6000 92.4000 157.0000 92.8000 ;
	    RECT 157.5000 92.7000 157.9000 92.8000 ;
	    RECT 157.5000 92.4000 158.9000 92.7000 ;
	    RECT 158.6000 92.1000 158.9000 92.4000 ;
	    RECT 160.6000 92.1000 161.0000 92.5000 ;
	    RECT 163.0000 92.1000 163.4000 93.3000 ;
	    RECT 165.4000 92.8000 165.8000 93.2000 ;
	    RECT 166.3000 93.1000 166.6000 94.9000 ;
	    RECT 167.8000 94.8000 168.2000 94.9000 ;
	    RECT 167.0000 94.1000 167.4000 94.6000 ;
	    RECT 169.4000 94.1000 169.8000 99.9000 ;
	    RECT 171.0000 96.2000 171.4000 99.9000 ;
	    RECT 172.6000 96.2000 173.0000 99.9000 ;
	    RECT 171.0000 95.9000 173.0000 96.2000 ;
	    RECT 173.4000 95.9000 173.8000 99.9000 ;
	    RECT 171.4000 95.2000 171.8000 95.4000 ;
	    RECT 173.4000 95.2000 173.7000 95.9000 ;
	    RECT 174.2000 95.7000 174.6000 99.9000 ;
	    RECT 176.4000 98.2000 176.8000 99.9000 ;
	    RECT 175.8000 97.9000 176.8000 98.2000 ;
	    RECT 178.6000 97.9000 179.0000 99.9000 ;
	    RECT 180.7000 97.9000 181.3000 99.9000 ;
	    RECT 175.8000 97.5000 176.2000 97.9000 ;
	    RECT 178.6000 97.6000 178.9000 97.9000 ;
	    RECT 177.5000 97.3000 179.3000 97.6000 ;
	    RECT 180.6000 97.5000 181.0000 97.9000 ;
	    RECT 177.5000 97.2000 177.9000 97.3000 ;
	    RECT 178.9000 97.2000 179.3000 97.3000 ;
	    RECT 175.8000 96.5000 176.2000 96.6000 ;
	    RECT 178.1000 96.5000 178.5000 96.6000 ;
	    RECT 175.8000 96.2000 178.5000 96.5000 ;
	    RECT 178.8000 96.5000 179.9000 96.8000 ;
	    RECT 178.8000 95.9000 179.1000 96.5000 ;
	    RECT 179.5000 96.4000 179.9000 96.5000 ;
	    RECT 180.7000 96.6000 181.4000 97.0000 ;
	    RECT 180.7000 96.1000 181.0000 96.6000 ;
	    RECT 176.7000 95.7000 179.1000 95.9000 ;
	    RECT 174.2000 95.6000 179.1000 95.7000 ;
	    RECT 179.8000 95.8000 181.0000 96.1000 ;
	    RECT 174.2000 95.5000 177.1000 95.6000 ;
	    RECT 174.2000 95.4000 177.0000 95.5000 ;
	    RECT 171.0000 94.9000 171.8000 95.2000 ;
	    RECT 172.6000 94.9000 173.8000 95.2000 ;
	    RECT 177.4000 95.1000 177.8000 95.2000 ;
	    RECT 171.0000 94.8000 171.4000 94.9000 ;
	    RECT 167.0000 93.8000 169.8000 94.1000 ;
	    RECT 169.4000 93.1000 169.8000 93.8000 ;
	    RECT 170.2000 93.4000 170.6000 94.2000 ;
	    RECT 171.8000 93.8000 172.2000 94.6000 ;
	    RECT 165.5000 92.4000 165.9000 92.8000 ;
	    RECT 164.6000 92.1000 165.0000 92.2000 ;
	    RECT 155.8000 91.8000 156.8000 92.1000 ;
	    RECT 156.4000 91.1000 156.8000 91.8000 ;
	    RECT 158.6000 91.1000 159.0000 92.1000 ;
	    RECT 160.6000 91.8000 161.3000 92.1000 ;
	    RECT 160.7000 91.1000 161.3000 91.8000 ;
	    RECT 163.0000 91.8000 165.0000 92.1000 ;
	    RECT 163.0000 91.1000 163.4000 91.8000 ;
	    RECT 166.2000 91.1000 166.6000 93.1000 ;
	    RECT 168.9000 92.8000 169.8000 93.1000 ;
	    RECT 172.6000 93.1000 172.9000 94.9000 ;
	    RECT 173.4000 94.8000 173.8000 94.9000 ;
	    RECT 175.3000 94.8000 177.8000 95.1000 ;
	    RECT 175.3000 94.7000 175.7000 94.8000 ;
	    RECT 176.1000 94.2000 176.5000 94.3000 ;
	    RECT 179.8000 94.2000 180.1000 95.8000 ;
	    RECT 183.0000 95.6000 183.4000 99.9000 ;
	    RECT 181.3000 95.3000 183.4000 95.6000 ;
	    RECT 181.3000 95.2000 181.7000 95.3000 ;
	    RECT 182.1000 94.9000 182.5000 95.0000 ;
	    RECT 180.6000 94.6000 182.5000 94.9000 ;
	    RECT 180.6000 94.5000 181.0000 94.6000 ;
	    RECT 174.6000 93.9000 180.1000 94.2000 ;
	    RECT 174.6000 93.8000 175.4000 93.9000 ;
	    RECT 168.9000 91.1000 169.3000 92.8000 ;
	    RECT 172.6000 91.1000 173.0000 93.1000 ;
	    RECT 173.4000 92.8000 173.8000 93.2000 ;
	    RECT 173.3000 92.4000 173.7000 92.8000 ;
	    RECT 174.2000 91.1000 174.6000 93.5000 ;
	    RECT 176.7000 92.8000 177.0000 93.9000 ;
	    RECT 179.5000 93.8000 179.9000 93.9000 ;
	    RECT 183.0000 93.6000 183.4000 95.3000 ;
	    RECT 181.5000 93.3000 183.4000 93.6000 ;
	    RECT 183.8000 93.4000 184.2000 94.2000 ;
	    RECT 181.5000 93.2000 181.9000 93.3000 ;
	    RECT 175.8000 92.1000 176.2000 92.5000 ;
	    RECT 176.6000 92.4000 177.0000 92.8000 ;
	    RECT 177.5000 92.7000 177.9000 92.8000 ;
	    RECT 177.5000 92.4000 178.9000 92.7000 ;
	    RECT 178.6000 92.1000 178.9000 92.4000 ;
	    RECT 180.6000 92.1000 181.0000 92.5000 ;
	    RECT 175.8000 91.8000 176.8000 92.1000 ;
	    RECT 176.4000 91.1000 176.8000 91.8000 ;
	    RECT 178.6000 91.1000 179.0000 92.1000 ;
	    RECT 180.6000 91.8000 181.3000 92.1000 ;
	    RECT 180.7000 91.1000 181.3000 91.8000 ;
	    RECT 183.0000 91.1000 183.4000 93.3000 ;
	    RECT 184.6000 93.1000 185.0000 99.9000 ;
	    RECT 185.4000 95.8000 185.8000 96.6000 ;
	    RECT 187.5000 96.2000 187.9000 99.9000 ;
	    RECT 188.2000 96.8000 188.6000 97.2000 ;
	    RECT 188.3000 96.2000 188.6000 96.8000 ;
	    RECT 187.0000 95.8000 188.0000 96.2000 ;
	    RECT 188.3000 96.1000 189.0000 96.2000 ;
	    RECT 189.4000 96.1000 189.8000 99.9000 ;
	    RECT 188.3000 95.9000 189.8000 96.1000 ;
	    RECT 188.6000 95.8000 189.8000 95.9000 ;
	    RECT 187.0000 94.4000 187.4000 95.2000 ;
	    RECT 187.7000 94.2000 188.0000 95.8000 ;
	    RECT 186.2000 94.1000 186.6000 94.2000 ;
	    RECT 186.2000 93.8000 187.0000 94.1000 ;
	    RECT 187.7000 93.8000 189.0000 94.2000 ;
	    RECT 186.6000 93.6000 187.0000 93.8000 ;
	    RECT 186.3000 93.1000 188.1000 93.3000 ;
	    RECT 188.6000 93.1000 188.9000 93.8000 ;
	    RECT 184.6000 92.8000 185.5000 93.1000 ;
	    RECT 185.1000 92.2000 185.5000 92.8000 ;
	    RECT 186.2000 93.0000 188.2000 93.1000 ;
	    RECT 185.1000 91.8000 185.8000 92.2000 ;
	    RECT 185.1000 91.1000 185.5000 91.8000 ;
	    RECT 186.2000 91.1000 186.6000 93.0000 ;
	    RECT 187.8000 91.1000 188.2000 93.0000 ;
	    RECT 188.6000 91.1000 189.0000 93.1000 ;
	    RECT 189.4000 91.1000 189.8000 95.8000 ;
	    RECT 191.0000 95.7000 191.4000 99.9000 ;
	    RECT 193.2000 98.2000 193.6000 99.9000 ;
	    RECT 192.6000 97.9000 193.6000 98.2000 ;
	    RECT 195.4000 97.9000 195.8000 99.9000 ;
	    RECT 197.5000 97.9000 198.1000 99.9000 ;
	    RECT 192.6000 97.5000 193.0000 97.9000 ;
	    RECT 195.4000 97.6000 195.7000 97.9000 ;
	    RECT 194.3000 97.3000 196.1000 97.6000 ;
	    RECT 197.4000 97.5000 197.8000 97.9000 ;
	    RECT 194.3000 97.2000 194.7000 97.3000 ;
	    RECT 195.7000 97.2000 196.1000 97.3000 ;
	    RECT 192.6000 96.5000 193.0000 96.6000 ;
	    RECT 194.9000 96.5000 195.3000 96.6000 ;
	    RECT 192.6000 96.2000 195.3000 96.5000 ;
	    RECT 195.6000 96.5000 196.7000 96.8000 ;
	    RECT 195.6000 95.9000 195.9000 96.5000 ;
	    RECT 196.3000 96.4000 196.7000 96.5000 ;
	    RECT 197.5000 96.6000 198.2000 97.0000 ;
	    RECT 197.5000 96.1000 197.8000 96.6000 ;
	    RECT 193.5000 95.7000 195.9000 95.9000 ;
	    RECT 191.0000 95.6000 195.9000 95.7000 ;
	    RECT 196.6000 95.8000 197.8000 96.1000 ;
	    RECT 191.0000 95.5000 193.9000 95.6000 ;
	    RECT 191.0000 95.4000 193.8000 95.5000 ;
	    RECT 196.6000 95.2000 196.9000 95.8000 ;
	    RECT 199.8000 95.6000 200.2000 99.9000 ;
	    RECT 200.6000 95.9000 201.0000 99.9000 ;
	    RECT 201.4000 96.2000 201.8000 99.9000 ;
	    RECT 203.0000 96.2000 203.4000 99.9000 ;
	    RECT 204.2000 96.8000 204.6000 97.2000 ;
	    RECT 204.2000 96.2000 204.5000 96.8000 ;
	    RECT 204.9000 96.2000 205.3000 99.9000 ;
	    RECT 201.4000 95.9000 203.4000 96.2000 ;
	    RECT 203.8000 95.9000 204.5000 96.2000 ;
	    RECT 204.8000 95.9000 205.3000 96.2000 ;
	    RECT 198.1000 95.3000 200.2000 95.6000 ;
	    RECT 198.1000 95.2000 198.5000 95.3000 ;
	    RECT 194.2000 95.1000 194.6000 95.2000 ;
	    RECT 195.0000 95.1000 195.4000 95.2000 ;
	    RECT 192.1000 94.8000 195.4000 95.1000 ;
	    RECT 196.6000 94.8000 197.0000 95.2000 ;
	    RECT 198.9000 94.9000 199.3000 95.0000 ;
	    RECT 192.1000 94.7000 192.5000 94.8000 ;
	    RECT 192.9000 94.2000 193.3000 94.3000 ;
	    RECT 196.6000 94.2000 196.9000 94.8000 ;
	    RECT 197.4000 94.6000 199.3000 94.9000 ;
	    RECT 197.4000 94.5000 197.8000 94.6000 ;
	    RECT 191.4000 93.9000 196.9000 94.2000 ;
	    RECT 191.4000 93.8000 192.2000 93.9000 ;
	    RECT 190.2000 92.4000 190.6000 93.2000 ;
	    RECT 191.0000 91.1000 191.4000 93.5000 ;
	    RECT 193.5000 92.8000 193.8000 93.9000 ;
	    RECT 196.3000 93.8000 196.7000 93.9000 ;
	    RECT 199.8000 93.6000 200.2000 95.3000 ;
	    RECT 200.7000 95.2000 201.0000 95.9000 ;
	    RECT 203.8000 95.8000 204.2000 95.9000 ;
	    RECT 202.6000 95.2000 203.0000 95.4000 ;
	    RECT 200.6000 94.9000 201.8000 95.2000 ;
	    RECT 202.6000 95.1000 203.4000 95.2000 ;
	    RECT 204.8000 95.1000 205.1000 95.9000 ;
	    RECT 202.6000 94.9000 205.1000 95.1000 ;
	    RECT 200.6000 94.8000 201.0000 94.9000 ;
	    RECT 198.3000 93.3000 200.2000 93.6000 ;
	    RECT 198.3000 93.2000 198.7000 93.3000 ;
	    RECT 192.6000 92.1000 193.0000 92.5000 ;
	    RECT 193.4000 92.4000 193.8000 92.8000 ;
	    RECT 194.3000 92.7000 194.7000 92.8000 ;
	    RECT 194.3000 92.4000 195.7000 92.7000 ;
	    RECT 195.4000 92.1000 195.7000 92.4000 ;
	    RECT 197.4000 92.1000 197.8000 92.5000 ;
	    RECT 192.6000 91.8000 193.6000 92.1000 ;
	    RECT 193.2000 91.1000 193.6000 91.8000 ;
	    RECT 195.4000 91.1000 195.8000 92.1000 ;
	    RECT 197.4000 91.8000 198.1000 92.1000 ;
	    RECT 197.5000 91.1000 198.1000 91.8000 ;
	    RECT 199.8000 91.1000 200.2000 93.3000 ;
	    RECT 200.6000 92.8000 201.0000 93.2000 ;
	    RECT 201.5000 93.1000 201.8000 94.9000 ;
	    RECT 203.0000 94.8000 205.1000 94.9000 ;
	    RECT 202.2000 93.8000 202.6000 94.6000 ;
	    RECT 204.8000 94.2000 205.1000 94.8000 ;
	    RECT 205.4000 94.4000 205.8000 95.2000 ;
	    RECT 203.8000 93.8000 205.1000 94.2000 ;
	    RECT 206.2000 94.1000 206.6000 94.2000 ;
	    RECT 205.8000 93.8000 206.6000 94.1000 ;
	    RECT 203.9000 93.1000 204.2000 93.8000 ;
	    RECT 205.8000 93.6000 206.2000 93.8000 ;
	    RECT 207.0000 93.4000 207.4000 94.2000 ;
	    RECT 204.7000 93.1000 206.5000 93.3000 ;
	    RECT 207.8000 93.1000 208.2000 99.9000 ;
	    RECT 208.6000 95.8000 209.0000 96.6000 ;
	    RECT 209.7000 96.3000 210.1000 99.9000 ;
	    RECT 209.7000 95.9000 210.6000 96.3000 ;
	    RECT 209.4000 94.8000 209.8000 95.6000 ;
	    RECT 210.2000 95.1000 210.5000 95.9000 ;
	    RECT 213.4000 95.8000 213.8000 96.6000 ;
	    RECT 213.4000 95.1000 213.7000 95.8000 ;
	    RECT 210.2000 94.8000 213.7000 95.1000 ;
	    RECT 210.2000 94.2000 210.5000 94.8000 ;
	    RECT 210.2000 93.8000 210.6000 94.2000 ;
	    RECT 200.7000 92.4000 201.1000 92.8000 ;
	    RECT 201.4000 91.1000 201.8000 93.1000 ;
	    RECT 203.8000 91.1000 204.2000 93.1000 ;
	    RECT 204.6000 93.0000 206.6000 93.1000 ;
	    RECT 204.6000 91.1000 205.0000 93.0000 ;
	    RECT 206.2000 91.1000 206.6000 93.0000 ;
	    RECT 207.8000 92.8000 208.7000 93.1000 ;
	    RECT 208.3000 92.2000 208.7000 92.8000 ;
	    RECT 208.3000 91.8000 209.0000 92.2000 ;
	    RECT 210.2000 92.1000 210.5000 93.8000 ;
	    RECT 211.0000 92.4000 211.4000 93.2000 ;
	    RECT 212.6000 93.1000 213.0000 93.2000 ;
	    RECT 214.2000 93.1000 214.6000 99.9000 ;
	    RECT 215.8000 96.2000 216.2000 99.9000 ;
	    RECT 216.7000 96.2000 217.1000 96.3000 ;
	    RECT 215.8000 95.9000 217.1000 96.2000 ;
	    RECT 218.0000 95.9000 218.8000 99.9000 ;
	    RECT 219.8000 96.2000 220.2000 96.3000 ;
	    RECT 220.6000 96.2000 221.0000 99.9000 ;
	    RECT 219.8000 95.9000 221.0000 96.2000 ;
	    RECT 221.7000 99.2000 222.1000 99.9000 ;
	    RECT 221.7000 98.8000 222.6000 99.2000 ;
	    RECT 221.7000 96.3000 222.1000 98.8000 ;
	    RECT 221.7000 95.9000 222.6000 96.3000 ;
	    RECT 223.8000 96.2000 224.2000 99.9000 ;
	    RECT 225.4000 96.4000 225.8000 99.9000 ;
	    RECT 223.8000 95.9000 225.1000 96.2000 ;
	    RECT 225.4000 95.9000 225.9000 96.4000 ;
	    RECT 217.3000 95.2000 217.7000 95.3000 ;
	    RECT 218.3000 95.2000 218.6000 95.9000 ;
	    RECT 216.9000 94.9000 217.7000 95.2000 ;
	    RECT 216.9000 94.8000 217.3000 94.9000 ;
	    RECT 218.2000 94.8000 218.6000 95.2000 ;
	    RECT 221.4000 94.8000 221.8000 95.6000 ;
	    RECT 217.6000 94.3000 218.0000 94.4000 ;
	    RECT 216.6000 94.2000 218.0000 94.3000 ;
	    RECT 215.0000 93.4000 215.4000 94.2000 ;
	    RECT 215.8000 94.0000 218.0000 94.2000 ;
	    RECT 218.3000 94.2000 218.6000 94.8000 ;
	    RECT 222.2000 94.2000 222.5000 95.9000 ;
	    RECT 223.8000 94.8000 224.3000 95.2000 ;
	    RECT 223.9000 94.4000 224.3000 94.8000 ;
	    RECT 224.8000 94.9000 225.1000 95.9000 ;
	    RECT 224.8000 94.5000 225.3000 94.9000 ;
	    RECT 215.8000 93.9000 216.9000 94.0000 ;
	    RECT 218.3000 93.9000 218.8000 94.2000 ;
	    RECT 215.8000 93.8000 216.6000 93.9000 ;
	    RECT 216.7000 93.4000 217.1000 93.5000 ;
	    RECT 212.6000 92.8000 214.6000 93.1000 ;
	    RECT 215.8000 93.1000 217.1000 93.4000 ;
	    RECT 217.4000 93.2000 218.2000 93.6000 ;
	    RECT 208.3000 91.1000 208.7000 91.8000 ;
	    RECT 210.2000 91.1000 210.6000 92.1000 ;
	    RECT 213.7000 91.1000 214.1000 92.8000 ;
	    RECT 215.8000 91.1000 216.2000 93.1000 ;
	    RECT 218.5000 92.9000 218.8000 93.9000 ;
	    RECT 219.2000 93.8000 219.6000 94.2000 ;
	    RECT 222.2000 93.8000 222.6000 94.2000 ;
	    RECT 219.2000 93.6000 219.5000 93.8000 ;
	    RECT 219.1000 93.2000 219.5000 93.6000 ;
	    RECT 219.8000 93.4000 220.2000 93.5000 ;
	    RECT 219.8000 93.1000 221.0000 93.4000 ;
	    RECT 218.0000 92.2000 218.8000 92.9000 ;
	    RECT 217.4000 91.8000 218.8000 92.2000 ;
	    RECT 218.0000 91.1000 218.8000 91.8000 ;
	    RECT 220.6000 91.1000 221.0000 93.1000 ;
	    RECT 222.2000 92.1000 222.5000 93.8000 ;
	    RECT 224.8000 93.7000 225.1000 94.5000 ;
	    RECT 225.6000 94.2000 225.9000 95.9000 ;
	    RECT 225.4000 93.8000 225.9000 94.2000 ;
	    RECT 223.8000 93.4000 225.1000 93.7000 ;
	    RECT 223.0000 92.4000 223.4000 93.2000 ;
	    RECT 222.2000 91.1000 222.6000 92.1000 ;
	    RECT 223.8000 91.1000 224.2000 93.4000 ;
	    RECT 225.6000 93.1000 225.9000 93.8000 ;
	    RECT 225.4000 92.8000 225.9000 93.1000 ;
	    RECT 225.4000 91.1000 225.8000 92.8000 ;
	    RECT 227.0000 91.1000 227.4000 99.9000 ;
	    RECT 227.8000 96.1000 228.2000 96.2000 ;
	    RECT 228.6000 96.1000 229.0000 96.6000 ;
	    RECT 227.8000 95.8000 229.0000 96.1000 ;
	    RECT 227.8000 93.1000 228.2000 93.2000 ;
	    RECT 229.4000 93.1000 229.8000 99.9000 ;
	    RECT 231.0000 95.8000 231.4000 96.6000 ;
	    RECT 230.2000 93.4000 230.6000 94.2000 ;
	    RECT 231.8000 93.1000 232.2000 99.9000 ;
	    RECT 233.4000 96.2000 233.8000 99.9000 ;
	    RECT 235.0000 96.4000 235.4000 99.9000 ;
	    RECT 233.4000 95.9000 234.7000 96.2000 ;
	    RECT 235.0000 95.9000 235.5000 96.4000 ;
	    RECT 236.9000 96.2000 237.3000 99.9000 ;
	    RECT 232.6000 95.1000 233.0000 95.2000 ;
	    RECT 233.4000 95.1000 233.9000 95.2000 ;
	    RECT 232.6000 94.8000 233.9000 95.1000 ;
	    RECT 233.5000 94.4000 233.9000 94.8000 ;
	    RECT 234.4000 94.9000 234.7000 95.9000 ;
	    RECT 234.4000 94.5000 234.9000 94.9000 ;
	    RECT 232.6000 93.4000 233.0000 94.2000 ;
	    RECT 234.4000 93.7000 234.7000 94.5000 ;
	    RECT 235.2000 94.2000 235.5000 95.9000 ;
	    RECT 236.6000 95.9000 237.3000 96.2000 ;
	    RECT 236.6000 95.2000 236.9000 95.9000 ;
	    RECT 239.0000 95.6000 239.4000 99.9000 ;
	    RECT 239.8000 95.8000 240.2000 96.6000 ;
	    RECT 237.4000 95.4000 239.4000 95.6000 ;
	    RECT 237.3000 95.3000 239.4000 95.4000 ;
	    RECT 236.6000 94.8000 237.0000 95.2000 ;
	    RECT 237.3000 95.0000 237.7000 95.3000 ;
	    RECT 235.0000 94.1000 235.5000 94.2000 ;
	    RECT 235.8000 94.1000 236.2000 94.2000 ;
	    RECT 235.0000 93.8000 236.2000 94.1000 ;
	    RECT 233.4000 93.4000 234.7000 93.7000 ;
	    RECT 227.8000 92.8000 229.8000 93.1000 ;
	    RECT 231.3000 92.8000 232.2000 93.1000 ;
	    RECT 227.8000 92.4000 228.2000 92.8000 ;
	    RECT 228.9000 91.1000 229.3000 92.8000 ;
	    RECT 231.3000 92.2000 231.7000 92.8000 ;
	    RECT 231.3000 91.8000 232.2000 92.2000 ;
	    RECT 231.3000 91.1000 231.7000 91.8000 ;
	    RECT 233.4000 91.1000 233.8000 93.4000 ;
	    RECT 235.2000 93.1000 235.5000 93.8000 ;
	    RECT 235.0000 92.8000 235.5000 93.1000 ;
	    RECT 236.6000 93.1000 236.9000 94.8000 ;
	    RECT 237.3000 93.5000 237.6000 95.0000 ;
	    RECT 238.0000 94.2000 238.4000 94.6000 ;
	    RECT 238.1000 93.8000 238.6000 94.2000 ;
	    RECT 237.3000 93.2000 238.5000 93.5000 ;
	    RECT 235.0000 91.1000 235.4000 92.8000 ;
	    RECT 236.6000 91.1000 237.0000 93.1000 ;
	    RECT 238.2000 92.1000 238.5000 93.2000 ;
	    RECT 239.0000 92.4000 239.4000 93.2000 ;
	    RECT 240.6000 93.1000 241.0000 99.9000 ;
	    RECT 243.5000 96.3000 243.9000 99.9000 ;
	    RECT 243.0000 95.9000 243.9000 96.3000 ;
	    RECT 244.9000 96.3000 245.3000 99.9000 ;
	    RECT 248.3000 96.3000 248.7000 99.9000 ;
	    RECT 244.9000 95.9000 245.8000 96.3000 ;
	    RECT 247.8000 95.9000 248.7000 96.3000 ;
	    RECT 249.4000 97.5000 249.8000 99.5000 ;
	    RECT 251.5000 99.2000 251.9000 99.9000 ;
	    RECT 251.5000 98.8000 252.2000 99.2000 ;
	    RECT 243.1000 94.2000 243.4000 95.9000 ;
	    RECT 243.8000 95.1000 244.2000 95.6000 ;
	    RECT 244.6000 95.1000 245.0000 95.6000 ;
	    RECT 243.8000 94.8000 245.0000 95.1000 ;
	    RECT 241.4000 93.4000 241.8000 94.2000 ;
	    RECT 243.0000 93.8000 243.4000 94.2000 ;
	    RECT 240.1000 92.8000 241.0000 93.1000 ;
	    RECT 240.1000 92.2000 240.5000 92.8000 ;
	    RECT 242.2000 92.4000 242.6000 93.2000 ;
	    RECT 243.1000 92.2000 243.4000 93.8000 ;
	    RECT 238.2000 91.1000 238.6000 92.1000 ;
	    RECT 240.1000 91.8000 241.0000 92.2000 ;
	    RECT 240.1000 91.1000 240.5000 91.8000 ;
	    RECT 243.0000 91.1000 243.4000 92.2000 ;
	    RECT 245.4000 94.2000 245.7000 95.9000 ;
	    RECT 247.9000 94.2000 248.2000 95.9000 ;
	    RECT 249.4000 95.8000 249.7000 97.5000 ;
	    RECT 251.5000 96.4000 251.9000 98.8000 ;
	    RECT 251.5000 96.1000 252.3000 96.4000 ;
	    RECT 255.5000 96.3000 255.9000 99.9000 ;
	    RECT 248.6000 94.8000 249.0000 95.6000 ;
	    RECT 249.4000 95.5000 251.3000 95.8000 ;
	    RECT 249.4000 94.4000 249.8000 95.2000 ;
	    RECT 250.2000 94.4000 250.6000 95.2000 ;
	    RECT 251.0000 94.5000 251.3000 95.5000 ;
	    RECT 245.4000 93.8000 245.8000 94.2000 ;
	    RECT 247.8000 93.8000 248.2000 94.2000 ;
	    RECT 251.0000 94.1000 251.7000 94.5000 ;
	    RECT 252.0000 94.2000 252.3000 96.1000 ;
	    RECT 255.0000 95.9000 255.9000 96.3000 ;
	    RECT 256.6000 96.2000 257.0000 99.9000 ;
	    RECT 257.5000 96.2000 257.9000 96.3000 ;
	    RECT 256.6000 95.9000 257.9000 96.2000 ;
	    RECT 258.8000 95.9000 259.6000 99.9000 ;
	    RECT 260.6000 96.2000 261.0000 96.3000 ;
	    RECT 261.4000 96.2000 261.8000 99.9000 ;
	    RECT 260.6000 95.9000 261.8000 96.2000 ;
	    RECT 262.2000 96.2000 262.6000 99.9000 ;
	    RECT 264.4000 97.2000 265.2000 99.9000 ;
	    RECT 263.8000 96.8000 265.2000 97.2000 ;
	    RECT 263.0000 96.2000 263.4000 96.3000 ;
	    RECT 264.4000 96.2000 265.2000 96.8000 ;
	    RECT 262.2000 95.9000 263.4000 96.2000 ;
	    RECT 264.2000 95.9000 265.2000 96.2000 ;
	    RECT 266.3000 96.2000 266.7000 96.3000 ;
	    RECT 267.0000 96.2000 267.4000 99.9000 ;
	    RECT 266.3000 95.9000 267.4000 96.2000 ;
	    RECT 268.1000 96.3000 268.5000 99.9000 ;
	    RECT 268.1000 95.9000 269.0000 96.3000 ;
	    RECT 252.6000 95.1000 253.0000 95.6000 ;
	    RECT 253.4000 95.1000 253.8000 95.2000 ;
	    RECT 252.6000 94.8000 253.8000 95.1000 ;
	    RECT 255.1000 94.2000 255.4000 95.9000 ;
	    RECT 258.1000 95.2000 258.5000 95.3000 ;
	    RECT 259.1000 95.2000 259.4000 95.9000 ;
	    RECT 264.2000 95.2000 264.5000 95.9000 ;
	    RECT 266.3000 95.6000 266.6000 95.9000 ;
	    RECT 264.9000 95.3000 266.6000 95.6000 ;
	    RECT 264.9000 95.2000 265.3000 95.3000 ;
	    RECT 257.7000 94.9000 258.5000 95.2000 ;
	    RECT 257.7000 94.8000 258.1000 94.9000 ;
	    RECT 259.0000 94.8000 259.4000 95.2000 ;
	    RECT 263.8000 94.9000 264.5000 95.2000 ;
	    RECT 267.8000 95.1000 268.2000 95.6000 ;
	    RECT 266.0000 94.9000 266.4000 95.0000 ;
	    RECT 263.8000 94.8000 264.7000 94.9000 ;
	    RECT 258.4000 94.3000 258.8000 94.4000 ;
	    RECT 257.4000 94.2000 258.8000 94.3000 ;
	    RECT 251.0000 93.9000 251.5000 94.1000 ;
	    RECT 245.4000 92.2000 245.7000 93.8000 ;
	    RECT 246.2000 92.4000 246.6000 93.2000 ;
	    RECT 247.0000 92.4000 247.4000 93.2000 ;
	    RECT 247.9000 92.2000 248.2000 93.8000 ;
	    RECT 245.4000 91.1000 245.8000 92.2000 ;
	    RECT 247.8000 91.1000 248.2000 92.2000 ;
	    RECT 249.4000 93.6000 251.5000 93.9000 ;
	    RECT 252.0000 93.8000 253.0000 94.2000 ;
	    RECT 255.0000 94.1000 255.4000 94.2000 ;
	    RECT 256.6000 94.1000 258.8000 94.2000 ;
	    RECT 255.0000 94.0000 258.8000 94.1000 ;
	    RECT 259.1000 94.2000 259.4000 94.8000 ;
	    RECT 264.2000 94.6000 264.7000 94.8000 ;
	    RECT 255.0000 93.9000 257.7000 94.0000 ;
	    RECT 259.1000 93.9000 259.6000 94.2000 ;
	    RECT 255.0000 93.8000 257.4000 93.9000 ;
	    RECT 249.4000 92.5000 249.7000 93.6000 ;
	    RECT 252.0000 93.5000 252.3000 93.8000 ;
	    RECT 251.9000 93.3000 252.3000 93.5000 ;
	    RECT 251.5000 93.0000 252.3000 93.3000 ;
	    RECT 249.4000 91.5000 249.8000 92.5000 ;
	    RECT 251.5000 91.5000 251.9000 93.0000 ;
	    RECT 254.2000 92.4000 254.6000 93.2000 ;
	    RECT 255.1000 92.1000 255.4000 93.8000 ;
	    RECT 257.5000 93.4000 257.9000 93.5000 ;
	    RECT 255.0000 91.1000 255.4000 92.1000 ;
	    RECT 256.6000 93.1000 257.9000 93.4000 ;
	    RECT 258.2000 93.2000 259.0000 93.6000 ;
	    RECT 256.6000 91.1000 257.0000 93.1000 ;
	    RECT 259.3000 92.9000 259.6000 93.9000 ;
	    RECT 260.0000 93.8000 260.4000 94.2000 ;
	    RECT 263.6000 93.8000 264.0000 94.2000 ;
	    RECT 260.0000 93.6000 260.3000 93.8000 ;
	    RECT 259.9000 93.2000 260.3000 93.6000 ;
	    RECT 263.7000 93.6000 264.0000 93.8000 ;
	    RECT 260.6000 93.4000 261.0000 93.5000 ;
	    RECT 263.0000 93.4000 263.4000 93.5000 ;
	    RECT 260.6000 93.1000 261.8000 93.4000 ;
	    RECT 258.8000 92.2000 259.6000 92.9000 ;
	    RECT 258.2000 91.8000 259.6000 92.2000 ;
	    RECT 258.8000 91.1000 259.6000 91.8000 ;
	    RECT 261.4000 91.1000 261.8000 93.1000 ;
	    RECT 262.2000 93.1000 263.4000 93.4000 ;
	    RECT 263.7000 93.2000 264.1000 93.6000 ;
	    RECT 262.2000 91.1000 262.6000 93.1000 ;
	    RECT 264.4000 92.9000 264.7000 94.6000 ;
	    RECT 265.1000 94.6000 266.4000 94.9000 ;
	    RECT 267.0000 94.8000 268.2000 95.1000 ;
	    RECT 265.1000 94.3000 265.4000 94.6000 ;
	    RECT 265.0000 93.9000 265.4000 94.3000 ;
	    RECT 267.0000 94.2000 267.3000 94.8000 ;
	    RECT 268.6000 94.2000 268.9000 95.9000 ;
	    RECT 266.6000 94.1000 267.4000 94.2000 ;
	    RECT 265.7000 93.8000 267.4000 94.1000 ;
	    RECT 268.6000 93.8000 269.0000 94.2000 ;
	    RECT 265.7000 93.6000 266.0000 93.8000 ;
	    RECT 265.0000 93.3000 266.0000 93.6000 ;
	    RECT 266.3000 93.4000 266.7000 93.5000 ;
	    RECT 265.0000 93.2000 265.8000 93.3000 ;
	    RECT 266.3000 93.1000 267.4000 93.4000 ;
	    RECT 264.4000 91.1000 265.2000 92.9000 ;
	    RECT 267.0000 91.1000 267.4000 93.1000 ;
	    RECT 268.6000 92.2000 268.9000 93.8000 ;
	    RECT 268.6000 91.1000 269.0000 92.2000 ;
	    RECT 0.6000 87.9000 1.0000 89.9000 ;
	    RECT 1.4000 88.0000 1.8000 89.9000 ;
	    RECT 3.0000 88.0000 3.4000 89.9000 ;
	    RECT 1.4000 87.9000 3.4000 88.0000 ;
	    RECT 0.7000 87.2000 1.0000 87.9000 ;
	    RECT 1.5000 87.7000 3.3000 87.9000 ;
	    RECT 2.6000 87.2000 3.0000 87.4000 ;
	    RECT 0.6000 86.8000 1.9000 87.2000 ;
	    RECT 2.6000 87.1000 3.4000 87.2000 ;
	    RECT 3.8000 87.1000 4.2000 89.9000 ;
	    RECT 6.9000 89.2000 7.7000 89.9000 ;
	    RECT 6.9000 88.8000 8.2000 89.2000 ;
	    RECT 6.9000 87.9000 7.7000 88.8000 ;
	    RECT 2.6000 86.9000 4.2000 87.1000 ;
	    RECT 3.0000 86.8000 4.2000 86.9000 ;
	    RECT 1.6000 85.2000 1.9000 86.8000 ;
	    RECT 3.8000 86.1000 4.2000 86.8000 ;
	    RECT 7.1000 86.2000 7.4000 87.9000 ;
	    RECT 7.8000 87.1000 8.2000 87.2000 ;
	    RECT 9.4000 87.1000 9.8000 89.9000 ;
	    RECT 11.0000 87.9000 11.4000 89.9000 ;
	    RECT 13.2000 89.2000 14.0000 89.9000 ;
	    RECT 13.2000 88.8000 14.6000 89.2000 ;
	    RECT 13.2000 88.1000 14.0000 88.8000 ;
	    RECT 11.0000 87.6000 12.3000 87.9000 ;
	    RECT 11.9000 87.5000 12.3000 87.6000 ;
	    RECT 12.6000 87.4000 13.4000 87.8000 ;
	    RECT 13.7000 87.1000 14.0000 88.1000 ;
	    RECT 15.8000 87.9000 16.2000 89.9000 ;
	    RECT 16.9000 88.2000 17.3000 89.9000 ;
	    RECT 19.8000 88.9000 20.2000 89.9000 ;
	    RECT 16.9000 87.9000 17.8000 88.2000 ;
	    RECT 14.3000 87.4000 14.7000 87.8000 ;
	    RECT 15.0000 87.6000 16.2000 87.9000 ;
	    RECT 15.0000 87.5000 15.4000 87.6000 ;
	    RECT 7.8000 86.8000 9.8000 87.1000 ;
	    RECT 7.8000 86.6000 8.1000 86.8000 ;
	    RECT 7.7000 86.2000 8.1000 86.6000 ;
	    RECT 5.4000 86.1000 5.8000 86.2000 ;
	    RECT 3.8000 85.8000 6.2000 86.1000 ;
	    RECT 7.0000 85.8000 7.4000 86.2000 ;
	    RECT 0.6000 85.1000 1.0000 85.2000 ;
	    RECT 0.6000 84.8000 1.3000 85.1000 ;
	    RECT 1.6000 84.8000 2.6000 85.2000 ;
	    RECT 1.0000 84.2000 1.3000 84.8000 ;
	    RECT 1.0000 83.8000 1.4000 84.2000 ;
	    RECT 1.7000 81.1000 2.1000 84.8000 ;
	    RECT 3.8000 81.1000 4.2000 85.8000 ;
	    RECT 5.8000 85.6000 6.2000 85.8000 ;
	    RECT 7.1000 85.7000 7.4000 85.8000 ;
	    RECT 7.1000 85.4000 8.1000 85.7000 ;
	    RECT 7.8000 85.1000 8.1000 85.4000 ;
	    RECT 5.4000 84.8000 7.4000 85.1000 ;
	    RECT 5.4000 81.1000 5.8000 84.8000 ;
	    RECT 7.0000 81.4000 7.4000 84.8000 ;
	    RECT 7.8000 81.7000 8.2000 85.1000 ;
	    RECT 8.6000 81.4000 9.0000 85.1000 ;
	    RECT 7.0000 81.1000 9.0000 81.4000 ;
	    RECT 9.4000 81.1000 9.8000 86.8000 ;
	    RECT 13.5000 86.8000 14.0000 87.1000 ;
	    RECT 14.4000 87.2000 14.7000 87.4000 ;
	    RECT 14.4000 86.8000 14.8000 87.2000 ;
	    RECT 13.5000 86.2000 13.8000 86.8000 ;
	    RECT 12.1000 86.1000 12.5000 86.2000 ;
	    RECT 12.1000 85.8000 12.9000 86.1000 ;
	    RECT 13.4000 85.8000 13.8000 86.2000 ;
	    RECT 12.5000 85.7000 12.9000 85.8000 ;
	    RECT 13.5000 85.1000 13.8000 85.8000 ;
	    RECT 11.0000 84.8000 12.3000 85.1000 ;
	    RECT 11.0000 81.1000 11.4000 84.8000 ;
	    RECT 11.9000 84.7000 12.3000 84.8000 ;
	    RECT 13.2000 81.1000 14.0000 85.1000 ;
	    RECT 15.0000 84.8000 16.2000 85.1000 ;
	    RECT 15.0000 84.7000 15.4000 84.8000 ;
	    RECT 15.8000 81.1000 16.2000 84.8000 ;
	    RECT 16.6000 84.4000 17.0000 85.2000 ;
	    RECT 17.4000 81.1000 17.8000 87.9000 ;
	    RECT 19.0000 87.8000 19.4000 88.6000 ;
	    RECT 18.2000 87.1000 18.6000 87.6000 ;
	    RECT 19.9000 87.2000 20.2000 88.9000 ;
	    RECT 21.4000 87.9000 21.8000 89.9000 ;
	    RECT 23.6000 89.2000 24.4000 89.9000 ;
	    RECT 23.6000 88.8000 25.0000 89.2000 ;
	    RECT 23.6000 88.1000 24.4000 88.8000 ;
	    RECT 21.4000 87.6000 22.5000 87.9000 ;
	    RECT 22.1000 87.5000 22.5000 87.6000 ;
	    RECT 19.8000 87.1000 20.2000 87.2000 ;
	    RECT 18.2000 86.8000 20.2000 87.1000 ;
	    RECT 19.9000 85.1000 20.2000 86.8000 ;
	    RECT 23.4000 86.7000 23.8000 87.1000 ;
	    RECT 23.4000 86.4000 23.7000 86.7000 ;
	    RECT 20.6000 85.4000 21.0000 86.2000 ;
	    RECT 22.4000 86.1000 23.7000 86.4000 ;
	    RECT 24.1000 86.4000 24.4000 88.1000 ;
	    RECT 26.2000 87.9000 26.6000 89.9000 ;
	    RECT 25.4000 87.6000 26.6000 87.9000 ;
	    RECT 27.0000 87.9000 27.4000 89.9000 ;
	    RECT 29.2000 88.1000 30.0000 89.9000 ;
	    RECT 27.0000 87.6000 28.2000 87.9000 ;
	    RECT 25.4000 87.5000 25.8000 87.6000 ;
	    RECT 27.8000 87.5000 28.2000 87.6000 ;
	    RECT 29.2000 86.4000 29.5000 88.1000 ;
	    RECT 31.8000 87.9000 32.2000 89.9000 ;
	    RECT 31.1000 87.6000 32.2000 87.9000 ;
	    RECT 32.6000 87.9000 33.0000 89.9000 ;
	    RECT 34.8000 88.1000 35.6000 89.9000 ;
	    RECT 32.6000 87.6000 33.9000 87.9000 ;
	    RECT 31.1000 87.5000 31.5000 87.6000 ;
	    RECT 33.5000 87.5000 33.9000 87.6000 ;
	    RECT 34.2000 87.4000 35.0000 87.8000 ;
	    RECT 35.3000 87.1000 35.6000 88.1000 ;
	    RECT 37.4000 87.9000 37.8000 89.9000 ;
	    RECT 35.9000 87.4000 36.3000 87.8000 ;
	    RECT 36.6000 87.6000 37.8000 87.9000 ;
	    RECT 38.2000 87.7000 38.6000 89.9000 ;
	    RECT 40.3000 89.2000 40.9000 89.9000 ;
	    RECT 40.3000 88.9000 41.0000 89.2000 ;
	    RECT 42.6000 88.9000 43.0000 89.9000 ;
	    RECT 44.8000 89.2000 45.2000 89.9000 ;
	    RECT 44.8000 88.9000 45.8000 89.2000 ;
	    RECT 40.6000 88.5000 41.0000 88.9000 ;
	    RECT 42.7000 88.6000 43.0000 88.9000 ;
	    RECT 42.7000 88.3000 44.1000 88.6000 ;
	    RECT 43.7000 88.2000 44.1000 88.3000 ;
	    RECT 44.6000 88.2000 45.0000 88.6000 ;
	    RECT 45.4000 88.5000 45.8000 88.9000 ;
	    RECT 39.7000 87.7000 40.1000 87.8000 ;
	    RECT 36.6000 87.5000 37.0000 87.6000 ;
	    RECT 29.8000 86.7000 30.2000 87.1000 ;
	    RECT 24.1000 86.2000 24.6000 86.4000 ;
	    RECT 29.0000 86.2000 29.5000 86.4000 ;
	    RECT 24.1000 86.1000 25.0000 86.2000 ;
	    RECT 22.4000 86.0000 22.8000 86.1000 ;
	    RECT 24.3000 85.8000 25.0000 86.1000 ;
	    RECT 28.6000 86.1000 29.5000 86.2000 ;
	    RECT 29.9000 86.4000 30.2000 86.7000 ;
	    RECT 35.1000 86.8000 35.6000 87.1000 ;
	    RECT 36.0000 87.2000 36.3000 87.4000 ;
	    RECT 38.2000 87.4000 40.1000 87.7000 ;
	    RECT 36.0000 86.8000 36.4000 87.2000 ;
	    RECT 29.9000 86.1000 31.2000 86.4000 ;
	    RECT 35.1000 86.2000 35.4000 86.8000 ;
	    RECT 28.6000 85.8000 29.3000 86.1000 ;
	    RECT 30.8000 86.0000 31.2000 86.1000 ;
	    RECT 33.7000 86.1000 34.1000 86.2000 ;
	    RECT 33.7000 85.8000 34.5000 86.1000 ;
	    RECT 35.0000 85.8000 35.4000 86.2000 ;
	    RECT 23.5000 85.7000 23.9000 85.8000 ;
	    RECT 22.2000 85.4000 23.9000 85.7000 ;
	    RECT 22.2000 85.1000 22.5000 85.4000 ;
	    RECT 24.3000 85.1000 24.6000 85.8000 ;
	    RECT 29.0000 85.1000 29.3000 85.8000 ;
	    RECT 29.7000 85.7000 30.1000 85.8000 ;
	    RECT 34.1000 85.7000 34.5000 85.8000 ;
	    RECT 29.7000 85.4000 31.4000 85.7000 ;
	    RECT 31.1000 85.1000 31.4000 85.4000 ;
	    RECT 35.1000 85.1000 35.4000 85.8000 ;
	    RECT 38.2000 85.7000 38.6000 87.4000 ;
	    RECT 41.7000 87.1000 42.1000 87.2000 ;
	    RECT 44.6000 87.1000 44.9000 88.2000 ;
	    RECT 47.0000 87.5000 47.4000 89.9000 ;
	    RECT 48.6000 88.8000 49.0000 89.9000 ;
	    RECT 48.6000 87.2000 48.9000 88.8000 ;
	    RECT 49.4000 87.8000 49.8000 88.6000 ;
	    RECT 46.2000 87.1000 47.0000 87.2000 ;
	    RECT 41.5000 86.8000 47.0000 87.1000 ;
	    RECT 48.6000 86.8000 49.0000 87.2000 ;
	    RECT 50.8000 87.1000 51.2000 89.9000 ;
	    RECT 50.3000 86.9000 51.2000 87.1000 ;
	    RECT 53.4000 87.9000 53.8000 89.9000 ;
	    RECT 55.0000 88.9000 55.4000 89.9000 ;
	    RECT 50.3000 86.8000 51.1000 86.9000 ;
	    RECT 40.6000 86.4000 41.0000 86.5000 ;
	    RECT 39.1000 86.1000 41.0000 86.4000 ;
	    RECT 39.1000 86.0000 39.5000 86.1000 ;
	    RECT 39.9000 85.7000 40.3000 85.8000 ;
	    RECT 38.2000 85.4000 40.3000 85.7000 ;
	    RECT 19.8000 84.7000 20.7000 85.1000 ;
	    RECT 20.3000 81.1000 20.7000 84.7000 ;
	    RECT 21.4000 84.8000 22.5000 85.1000 ;
	    RECT 21.4000 81.1000 21.8000 84.8000 ;
	    RECT 22.1000 84.7000 22.5000 84.8000 ;
	    RECT 23.6000 84.8000 24.6000 85.1000 ;
	    RECT 25.4000 84.8000 26.6000 85.1000 ;
	    RECT 23.6000 81.1000 24.4000 84.8000 ;
	    RECT 25.4000 84.7000 25.8000 84.8000 ;
	    RECT 26.2000 81.1000 26.6000 84.8000 ;
	    RECT 27.0000 84.8000 28.2000 85.1000 ;
	    RECT 29.0000 84.8000 30.0000 85.1000 ;
	    RECT 27.0000 81.1000 27.4000 84.8000 ;
	    RECT 27.8000 84.7000 28.2000 84.8000 ;
	    RECT 29.2000 81.1000 30.0000 84.8000 ;
	    RECT 31.1000 84.8000 32.2000 85.1000 ;
	    RECT 31.1000 84.7000 31.5000 84.8000 ;
	    RECT 31.8000 81.1000 32.2000 84.8000 ;
	    RECT 32.6000 84.8000 33.9000 85.1000 ;
	    RECT 32.6000 81.1000 33.0000 84.8000 ;
	    RECT 33.5000 84.7000 33.9000 84.8000 ;
	    RECT 34.8000 81.1000 35.6000 85.1000 ;
	    RECT 36.6000 84.8000 37.8000 85.1000 ;
	    RECT 36.6000 84.7000 37.0000 84.8000 ;
	    RECT 37.4000 81.1000 37.8000 84.8000 ;
	    RECT 38.2000 81.1000 38.6000 85.4000 ;
	    RECT 41.5000 85.2000 41.8000 86.8000 ;
	    RECT 45.1000 86.7000 45.5000 86.8000 ;
	    RECT 44.6000 86.2000 45.0000 86.3000 ;
	    RECT 45.9000 86.2000 46.3000 86.3000 ;
	    RECT 43.8000 85.9000 46.3000 86.2000 ;
	    RECT 43.8000 85.8000 44.2000 85.9000 ;
	    RECT 44.6000 85.5000 47.4000 85.6000 ;
	    RECT 44.5000 85.4000 47.4000 85.5000 ;
	    RECT 47.8000 85.4000 48.2000 86.2000 ;
	    RECT 40.6000 84.9000 41.8000 85.2000 ;
	    RECT 42.5000 85.3000 47.4000 85.4000 ;
	    RECT 42.5000 85.1000 44.9000 85.3000 ;
	    RECT 40.6000 84.4000 40.9000 84.9000 ;
	    RECT 40.2000 84.0000 40.9000 84.4000 ;
	    RECT 41.7000 84.5000 42.1000 84.6000 ;
	    RECT 42.5000 84.5000 42.8000 85.1000 ;
	    RECT 41.7000 84.2000 42.8000 84.5000 ;
	    RECT 43.1000 84.5000 45.8000 84.8000 ;
	    RECT 43.1000 84.4000 43.5000 84.5000 ;
	    RECT 45.4000 84.4000 45.8000 84.5000 ;
	    RECT 42.3000 83.7000 42.7000 83.8000 ;
	    RECT 43.7000 83.7000 44.1000 83.8000 ;
	    RECT 40.6000 83.1000 41.0000 83.5000 ;
	    RECT 42.3000 83.4000 44.1000 83.7000 ;
	    RECT 42.7000 83.1000 43.0000 83.4000 ;
	    RECT 45.4000 83.1000 45.8000 83.5000 ;
	    RECT 40.3000 81.1000 40.9000 83.1000 ;
	    RECT 42.6000 81.1000 43.0000 83.1000 ;
	    RECT 44.8000 82.8000 45.8000 83.1000 ;
	    RECT 44.8000 81.1000 45.2000 82.8000 ;
	    RECT 47.0000 81.1000 47.4000 85.3000 ;
	    RECT 48.6000 85.1000 48.9000 86.8000 ;
	    RECT 50.3000 85.2000 50.6000 86.8000 ;
	    RECT 53.4000 86.2000 53.7000 87.9000 ;
	    RECT 55.0000 87.8000 55.3000 88.9000 ;
	    RECT 55.8000 87.8000 56.2000 88.6000 ;
	    RECT 56.9000 88.2000 57.3000 89.9000 ;
	    RECT 56.9000 87.9000 57.8000 88.2000 ;
	    RECT 60.6000 87.9000 61.0000 89.9000 ;
	    RECT 61.4000 88.0000 61.8000 89.9000 ;
	    RECT 63.0000 88.0000 63.4000 89.9000 ;
	    RECT 61.4000 87.9000 63.4000 88.0000 ;
	    RECT 54.1000 87.5000 55.3000 87.8000 ;
	    RECT 51.4000 85.8000 52.2000 86.2000 ;
	    RECT 53.4000 85.8000 53.8000 86.2000 ;
	    RECT 54.1000 86.0000 54.4000 87.5000 ;
	    RECT 54.9000 87.1000 55.4000 87.2000 ;
	    RECT 55.8000 87.1000 56.2000 87.2000 ;
	    RECT 54.9000 86.8000 56.2000 87.1000 ;
	    RECT 54.8000 86.4000 55.2000 86.8000 ;
	    RECT 48.1000 84.7000 49.0000 85.1000 ;
	    RECT 50.2000 84.8000 50.6000 85.2000 ;
	    RECT 52.6000 85.1000 53.0000 85.6000 ;
	    RECT 53.4000 85.1000 53.7000 85.8000 ;
	    RECT 54.1000 85.7000 54.5000 86.0000 ;
	    RECT 54.1000 85.6000 56.2000 85.7000 ;
	    RECT 54.2000 85.4000 56.2000 85.6000 ;
	    RECT 52.6000 84.8000 54.1000 85.1000 ;
	    RECT 48.1000 81.1000 48.5000 84.7000 ;
	    RECT 50.3000 83.5000 50.6000 84.8000 ;
	    RECT 51.0000 83.8000 51.4000 84.6000 ;
	    RECT 50.3000 83.2000 52.1000 83.5000 ;
	    RECT 50.3000 83.1000 50.6000 83.2000 ;
	    RECT 50.2000 81.1000 50.6000 83.1000 ;
	    RECT 51.8000 83.1000 52.1000 83.2000 ;
	    RECT 51.8000 81.1000 52.2000 83.1000 ;
	    RECT 53.7000 81.1000 54.1000 84.8000 ;
	    RECT 55.8000 81.1000 56.2000 85.4000 ;
	    RECT 56.6000 84.4000 57.0000 85.2000 ;
	    RECT 57.4000 81.1000 57.8000 87.9000 ;
	    RECT 58.2000 86.8000 58.6000 87.6000 ;
	    RECT 60.7000 87.2000 61.0000 87.9000 ;
	    RECT 61.5000 87.7000 63.3000 87.9000 ;
	    RECT 62.6000 87.2000 63.0000 87.4000 ;
	    RECT 60.6000 86.8000 61.9000 87.2000 ;
	    RECT 62.6000 86.9000 63.4000 87.2000 ;
	    RECT 64.4000 87.1000 64.8000 89.9000 ;
	    RECT 63.0000 86.8000 63.4000 86.9000 ;
	    RECT 63.9000 86.9000 64.8000 87.1000 ;
	    RECT 67.0000 87.7000 67.4000 89.9000 ;
	    RECT 69.1000 89.2000 69.7000 89.9000 ;
	    RECT 69.1000 88.9000 69.8000 89.2000 ;
	    RECT 71.4000 88.9000 71.8000 89.9000 ;
	    RECT 73.6000 89.2000 74.0000 89.9000 ;
	    RECT 73.6000 88.9000 74.6000 89.2000 ;
	    RECT 69.4000 88.5000 69.8000 88.9000 ;
	    RECT 71.5000 88.6000 71.8000 88.9000 ;
	    RECT 71.5000 88.3000 72.9000 88.6000 ;
	    RECT 72.5000 88.2000 72.9000 88.3000 ;
	    RECT 73.4000 88.2000 73.8000 88.6000 ;
	    RECT 74.2000 88.5000 74.6000 88.9000 ;
	    RECT 68.5000 87.7000 68.9000 87.8000 ;
	    RECT 67.0000 87.4000 68.9000 87.7000 ;
	    RECT 63.9000 86.8000 64.7000 86.9000 ;
	    RECT 59.0000 85.1000 59.4000 85.2000 ;
	    RECT 60.6000 85.1000 61.0000 85.2000 ;
	    RECT 61.6000 85.1000 61.9000 86.8000 ;
	    RECT 62.2000 85.8000 62.6000 86.6000 ;
	    RECT 63.9000 85.2000 64.2000 86.8000 ;
	    RECT 65.0000 85.8000 65.8000 86.2000 ;
	    RECT 67.0000 85.7000 67.4000 87.4000 ;
	    RECT 70.5000 87.1000 70.9000 87.2000 ;
	    RECT 73.4000 87.1000 73.7000 88.2000 ;
	    RECT 75.8000 87.5000 76.2000 89.9000 ;
	    RECT 77.4000 88.9000 77.8000 89.9000 ;
	    RECT 76.6000 87.8000 77.0000 88.6000 ;
	    RECT 77.5000 87.2000 77.8000 88.9000 ;
	    RECT 79.0000 87.5000 79.4000 89.9000 ;
	    RECT 81.2000 89.2000 81.6000 89.9000 ;
	    RECT 80.6000 88.9000 81.6000 89.2000 ;
	    RECT 83.4000 88.9000 83.8000 89.9000 ;
	    RECT 85.5000 89.2000 86.1000 89.9000 ;
	    RECT 85.4000 88.9000 86.1000 89.2000 ;
	    RECT 80.6000 88.5000 81.0000 88.9000 ;
	    RECT 83.4000 88.6000 83.7000 88.9000 ;
	    RECT 81.4000 88.2000 81.8000 88.6000 ;
	    RECT 82.3000 88.3000 83.7000 88.6000 ;
	    RECT 85.4000 88.5000 85.8000 88.9000 ;
	    RECT 82.3000 88.2000 82.7000 88.3000 ;
	    RECT 75.0000 87.1000 75.8000 87.2000 ;
	    RECT 70.3000 86.8000 75.8000 87.1000 ;
	    RECT 76.6000 86.8000 77.0000 87.2000 ;
	    RECT 77.4000 86.8000 77.8000 87.2000 ;
	    RECT 79.4000 87.1000 80.2000 87.2000 ;
	    RECT 81.5000 87.1000 81.8000 88.2000 ;
	    RECT 86.3000 87.7000 86.7000 87.8000 ;
	    RECT 87.8000 87.7000 88.2000 89.9000 ;
	    RECT 86.3000 87.4000 88.2000 87.7000 ;
	    RECT 84.3000 87.1000 84.7000 87.2000 ;
	    RECT 79.4000 86.8000 84.9000 87.1000 ;
	    RECT 69.4000 86.4000 69.8000 86.5000 ;
	    RECT 67.9000 86.1000 69.8000 86.4000 ;
	    RECT 67.9000 86.0000 68.3000 86.1000 ;
	    RECT 68.7000 85.7000 69.1000 85.8000 ;
	    RECT 59.0000 84.8000 61.3000 85.1000 ;
	    RECT 61.6000 84.8000 62.1000 85.1000 ;
	    RECT 63.8000 84.8000 64.2000 85.2000 ;
	    RECT 61.0000 84.2000 61.3000 84.8000 ;
	    RECT 61.0000 83.8000 61.4000 84.2000 ;
	    RECT 61.7000 81.1000 62.1000 84.8000 ;
	    RECT 63.9000 83.5000 64.2000 84.8000 ;
	    RECT 66.2000 84.8000 66.6000 85.6000 ;
	    RECT 67.0000 85.4000 69.1000 85.7000 ;
	    RECT 64.6000 83.8000 65.0000 84.6000 ;
	    RECT 66.2000 84.1000 66.5000 84.8000 ;
	    RECT 67.0000 84.1000 67.4000 85.4000 ;
	    RECT 70.3000 85.2000 70.6000 86.8000 ;
	    RECT 73.9000 86.7000 74.3000 86.8000 ;
	    RECT 73.4000 86.2000 73.8000 86.3000 ;
	    RECT 74.7000 86.2000 75.1000 86.3000 ;
	    RECT 72.6000 85.9000 75.1000 86.2000 ;
	    RECT 76.6000 86.1000 76.9000 86.8000 ;
	    RECT 77.5000 86.1000 77.8000 86.8000 ;
	    RECT 80.9000 86.7000 81.3000 86.8000 ;
	    RECT 80.1000 86.2000 80.5000 86.3000 ;
	    RECT 81.4000 86.2000 81.8000 86.3000 ;
	    RECT 84.6000 86.2000 84.9000 86.8000 ;
	    RECT 85.4000 86.4000 85.8000 86.5000 ;
	    RECT 72.6000 85.8000 73.0000 85.9000 ;
	    RECT 76.6000 85.8000 77.8000 86.1000 ;
	    RECT 73.4000 85.5000 76.2000 85.6000 ;
	    RECT 73.3000 85.4000 76.2000 85.5000 ;
	    RECT 69.4000 84.9000 70.6000 85.2000 ;
	    RECT 71.3000 85.3000 76.2000 85.4000 ;
	    RECT 71.3000 85.1000 73.7000 85.3000 ;
	    RECT 69.4000 84.4000 69.7000 84.9000 ;
	    RECT 66.2000 83.8000 67.4000 84.1000 ;
	    RECT 69.0000 84.0000 69.7000 84.4000 ;
	    RECT 70.5000 84.5000 70.9000 84.6000 ;
	    RECT 71.3000 84.5000 71.6000 85.1000 ;
	    RECT 70.5000 84.2000 71.6000 84.5000 ;
	    RECT 71.9000 84.5000 74.6000 84.8000 ;
	    RECT 71.9000 84.4000 72.3000 84.5000 ;
	    RECT 74.2000 84.4000 74.6000 84.5000 ;
	    RECT 63.9000 83.2000 65.7000 83.5000 ;
	    RECT 63.9000 83.1000 64.2000 83.2000 ;
	    RECT 63.8000 81.1000 64.2000 83.1000 ;
	    RECT 65.4000 83.1000 65.7000 83.2000 ;
	    RECT 65.4000 81.1000 65.8000 83.1000 ;
	    RECT 67.0000 81.1000 67.4000 83.8000 ;
	    RECT 71.1000 83.7000 71.5000 83.8000 ;
	    RECT 72.5000 83.7000 72.9000 83.8000 ;
	    RECT 69.4000 83.1000 69.8000 83.5000 ;
	    RECT 71.1000 83.4000 72.9000 83.7000 ;
	    RECT 71.5000 83.1000 71.8000 83.4000 ;
	    RECT 74.2000 83.1000 74.6000 83.5000 ;
	    RECT 69.1000 81.1000 69.7000 83.1000 ;
	    RECT 71.4000 81.1000 71.8000 83.1000 ;
	    RECT 73.6000 82.8000 74.6000 83.1000 ;
	    RECT 73.6000 81.1000 74.0000 82.8000 ;
	    RECT 75.8000 81.1000 76.2000 85.3000 ;
	    RECT 77.5000 85.1000 77.8000 85.8000 ;
	    RECT 78.2000 85.4000 78.6000 86.2000 ;
	    RECT 80.1000 85.9000 82.6000 86.2000 ;
	    RECT 82.2000 85.8000 82.6000 85.9000 ;
	    RECT 84.6000 85.8000 85.0000 86.2000 ;
	    RECT 85.4000 86.1000 87.3000 86.4000 ;
	    RECT 86.9000 86.0000 87.3000 86.1000 ;
	    RECT 79.0000 85.5000 81.8000 85.6000 ;
	    RECT 79.0000 85.4000 81.9000 85.5000 ;
	    RECT 79.0000 85.3000 83.9000 85.4000 ;
	    RECT 77.4000 84.7000 78.3000 85.1000 ;
	    RECT 77.9000 81.1000 78.3000 84.7000 ;
	    RECT 79.0000 81.1000 79.4000 85.3000 ;
	    RECT 81.5000 85.1000 83.9000 85.3000 ;
	    RECT 80.6000 84.5000 83.3000 84.8000 ;
	    RECT 80.6000 84.4000 81.0000 84.5000 ;
	    RECT 82.9000 84.4000 83.3000 84.5000 ;
	    RECT 83.6000 84.5000 83.9000 85.1000 ;
	    RECT 84.6000 85.2000 84.9000 85.8000 ;
	    RECT 86.1000 85.7000 86.5000 85.8000 ;
	    RECT 87.8000 85.7000 88.2000 87.4000 ;
	    RECT 86.1000 85.4000 88.2000 85.7000 ;
	    RECT 84.6000 84.9000 85.8000 85.2000 ;
	    RECT 84.3000 84.5000 84.7000 84.6000 ;
	    RECT 83.6000 84.2000 84.7000 84.5000 ;
	    RECT 85.5000 84.4000 85.8000 84.9000 ;
	    RECT 85.5000 84.0000 86.2000 84.4000 ;
	    RECT 82.3000 83.7000 82.7000 83.8000 ;
	    RECT 83.7000 83.7000 84.1000 83.8000 ;
	    RECT 80.6000 83.1000 81.0000 83.5000 ;
	    RECT 82.3000 83.4000 84.1000 83.7000 ;
	    RECT 83.4000 83.1000 83.7000 83.4000 ;
	    RECT 85.4000 83.1000 85.8000 83.5000 ;
	    RECT 80.6000 82.8000 81.6000 83.1000 ;
	    RECT 81.2000 81.1000 81.6000 82.8000 ;
	    RECT 83.4000 81.1000 83.8000 83.1000 ;
	    RECT 85.5000 81.1000 86.1000 83.1000 ;
	    RECT 87.8000 81.1000 88.2000 85.4000 ;
	    RECT 88.6000 87.7000 89.0000 89.9000 ;
	    RECT 90.7000 89.2000 91.3000 89.9000 ;
	    RECT 90.7000 88.9000 91.4000 89.2000 ;
	    RECT 93.0000 88.9000 93.4000 89.9000 ;
	    RECT 95.2000 89.2000 95.6000 89.9000 ;
	    RECT 95.2000 88.9000 96.2000 89.2000 ;
	    RECT 91.0000 88.5000 91.4000 88.9000 ;
	    RECT 93.1000 88.6000 93.4000 88.9000 ;
	    RECT 93.1000 88.3000 94.5000 88.6000 ;
	    RECT 94.1000 88.2000 94.5000 88.3000 ;
	    RECT 95.0000 88.2000 95.4000 88.6000 ;
	    RECT 95.8000 88.5000 96.2000 88.9000 ;
	    RECT 90.1000 87.7000 90.5000 87.8000 ;
	    RECT 88.6000 87.4000 90.5000 87.7000 ;
	    RECT 88.6000 85.7000 89.0000 87.4000 ;
	    RECT 92.1000 87.1000 92.5000 87.2000 ;
	    RECT 95.0000 87.1000 95.3000 88.2000 ;
	    RECT 97.4000 87.5000 97.8000 89.9000 ;
	    RECT 98.2000 88.0000 98.6000 89.9000 ;
	    RECT 99.8000 88.0000 100.2000 89.9000 ;
	    RECT 98.2000 87.9000 100.2000 88.0000 ;
	    RECT 100.6000 87.9000 101.0000 89.9000 ;
	    RECT 102.2000 88.2000 102.6000 89.9000 ;
	    RECT 102.1000 87.9000 102.6000 88.2000 ;
	    RECT 98.3000 87.7000 100.1000 87.9000 ;
	    RECT 98.6000 87.2000 99.0000 87.4000 ;
	    RECT 100.6000 87.2000 100.9000 87.9000 ;
	    RECT 102.1000 87.2000 102.4000 87.9000 ;
	    RECT 103.8000 87.6000 104.2000 89.9000 ;
	    RECT 102.9000 87.3000 104.2000 87.6000 ;
	    RECT 105.4000 87.6000 105.8000 89.9000 ;
	    RECT 107.0000 87.6000 107.4000 89.9000 ;
	    RECT 110.3000 88.2000 110.7000 88.6000 ;
	    RECT 108.6000 88.1000 109.0000 88.2000 ;
	    RECT 110.2000 88.1000 110.6000 88.2000 ;
	    RECT 108.6000 87.8000 110.6000 88.1000 ;
	    RECT 111.0000 87.9000 111.4000 89.9000 ;
	    RECT 96.6000 87.1000 97.4000 87.2000 ;
	    RECT 91.9000 86.8000 97.4000 87.1000 ;
	    RECT 98.2000 86.9000 99.0000 87.2000 ;
	    RECT 98.2000 86.8000 98.6000 86.9000 ;
	    RECT 99.7000 86.8000 101.0000 87.2000 ;
	    RECT 101.4000 87.1000 101.8000 87.2000 ;
	    RECT 102.1000 87.1000 102.6000 87.2000 ;
	    RECT 101.4000 86.8000 102.6000 87.1000 ;
	    RECT 91.0000 86.4000 91.4000 86.5000 ;
	    RECT 89.5000 86.1000 91.4000 86.4000 ;
	    RECT 89.5000 86.0000 89.9000 86.1000 ;
	    RECT 90.3000 85.7000 90.7000 85.8000 ;
	    RECT 88.6000 85.4000 90.7000 85.7000 ;
	    RECT 88.6000 81.1000 89.0000 85.4000 ;
	    RECT 91.9000 85.2000 92.2000 86.8000 ;
	    RECT 95.5000 86.7000 95.9000 86.8000 ;
	    RECT 96.3000 86.2000 96.7000 86.3000 ;
	    RECT 94.2000 85.9000 96.7000 86.2000 ;
	    RECT 98.2000 86.1000 98.6000 86.2000 ;
	    RECT 99.0000 86.1000 99.4000 86.6000 ;
	    RECT 94.2000 85.8000 94.6000 85.9000 ;
	    RECT 98.2000 85.8000 99.4000 86.1000 ;
	    RECT 99.7000 86.1000 100.0000 86.8000 ;
	    RECT 101.4000 86.1000 101.8000 86.2000 ;
	    RECT 99.7000 85.8000 101.8000 86.1000 ;
	    RECT 95.0000 85.5000 97.8000 85.6000 ;
	    RECT 94.9000 85.4000 97.8000 85.5000 ;
	    RECT 91.0000 84.9000 92.2000 85.2000 ;
	    RECT 92.9000 85.3000 97.8000 85.4000 ;
	    RECT 92.9000 85.1000 95.3000 85.3000 ;
	    RECT 91.0000 84.4000 91.3000 84.9000 ;
	    RECT 90.6000 84.0000 91.3000 84.4000 ;
	    RECT 92.1000 84.5000 92.5000 84.6000 ;
	    RECT 92.9000 84.5000 93.2000 85.1000 ;
	    RECT 92.1000 84.2000 93.2000 84.5000 ;
	    RECT 93.5000 84.5000 96.2000 84.8000 ;
	    RECT 93.5000 84.4000 93.9000 84.5000 ;
	    RECT 95.8000 84.4000 96.2000 84.5000 ;
	    RECT 92.7000 83.7000 93.1000 83.8000 ;
	    RECT 94.1000 83.7000 94.5000 83.8000 ;
	    RECT 91.0000 83.1000 91.4000 83.5000 ;
	    RECT 92.7000 83.4000 94.5000 83.7000 ;
	    RECT 93.1000 83.1000 93.4000 83.4000 ;
	    RECT 95.8000 83.1000 96.2000 83.5000 ;
	    RECT 90.7000 81.1000 91.3000 83.1000 ;
	    RECT 93.0000 81.1000 93.4000 83.1000 ;
	    RECT 95.2000 82.8000 96.2000 83.1000 ;
	    RECT 95.2000 81.1000 95.6000 82.8000 ;
	    RECT 97.4000 81.1000 97.8000 85.3000 ;
	    RECT 99.7000 85.1000 100.0000 85.8000 ;
	    RECT 100.6000 85.1000 101.0000 85.2000 ;
	    RECT 99.5000 84.8000 100.0000 85.1000 ;
	    RECT 100.3000 84.8000 101.0000 85.1000 ;
	    RECT 102.1000 85.1000 102.4000 86.8000 ;
	    RECT 102.9000 86.5000 103.2000 87.3000 ;
	    RECT 105.4000 87.2000 107.4000 87.6000 ;
	    RECT 102.7000 86.1000 103.2000 86.5000 ;
	    RECT 102.9000 85.1000 103.2000 86.1000 ;
	    RECT 103.7000 86.2000 104.1000 86.6000 ;
	    RECT 103.7000 86.1000 104.2000 86.2000 ;
	    RECT 104.6000 86.1000 105.0000 86.2000 ;
	    RECT 103.7000 85.8000 105.0000 86.1000 ;
	    RECT 105.4000 85.8000 105.8000 87.2000 ;
	    RECT 107.8000 86.8000 108.2000 87.6000 ;
	    RECT 110.2000 86.1000 110.6000 86.2000 ;
	    RECT 111.1000 86.1000 111.4000 87.9000 ;
	    RECT 115.2000 87.2000 115.6000 89.9000 ;
	    RECT 116.6000 87.8000 117.0000 88.6000 ;
	    RECT 111.8000 86.4000 112.2000 87.2000 ;
	    RECT 115.0000 87.1000 115.6000 87.2000 ;
	    RECT 115.0000 86.8000 116.1000 87.1000 ;
	    RECT 112.6000 86.1000 113.0000 86.2000 ;
	    RECT 110.2000 85.8000 111.4000 86.1000 ;
	    RECT 112.2000 85.8000 113.0000 86.1000 ;
	    RECT 105.4000 85.4000 107.4000 85.8000 ;
	    RECT 99.5000 81.1000 99.9000 84.8000 ;
	    RECT 100.3000 84.2000 100.6000 84.8000 ;
	    RECT 102.1000 84.6000 102.6000 85.1000 ;
	    RECT 102.9000 84.8000 104.2000 85.1000 ;
	    RECT 100.2000 83.8000 100.6000 84.2000 ;
	    RECT 102.2000 81.1000 102.6000 84.6000 ;
	    RECT 103.8000 81.1000 104.2000 84.8000 ;
	    RECT 105.4000 81.1000 105.8000 85.4000 ;
	    RECT 107.0000 81.1000 107.4000 85.4000 ;
	    RECT 110.3000 85.1000 110.6000 85.8000 ;
	    RECT 112.2000 85.6000 112.6000 85.8000 ;
	    RECT 110.2000 81.1000 110.6000 85.1000 ;
	    RECT 111.0000 84.8000 113.0000 85.1000 ;
	    RECT 113.4000 84.8000 113.8000 86.2000 ;
	    RECT 114.2000 85.8000 115.0000 86.2000 ;
	    RECT 115.8000 85.2000 116.1000 86.8000 ;
	    RECT 115.8000 84.8000 116.2000 85.2000 ;
	    RECT 117.4000 85.1000 117.8000 89.9000 ;
	    RECT 118.5000 89.2000 118.9000 89.9000 ;
	    RECT 118.2000 88.8000 118.9000 89.2000 ;
	    RECT 118.5000 88.2000 118.9000 88.8000 ;
	    RECT 118.5000 87.9000 119.4000 88.2000 ;
	    RECT 118.2000 85.1000 118.6000 85.2000 ;
	    RECT 117.4000 84.8000 118.6000 85.1000 ;
	    RECT 111.0000 81.1000 111.4000 84.8000 ;
	    RECT 112.6000 81.1000 113.0000 84.8000 ;
	    RECT 115.0000 83.8000 115.4000 84.6000 ;
	    RECT 115.8000 83.5000 116.1000 84.8000 ;
	    RECT 114.3000 83.2000 116.1000 83.5000 ;
	    RECT 114.3000 83.1000 114.6000 83.2000 ;
	    RECT 114.2000 81.1000 114.6000 83.1000 ;
	    RECT 115.8000 83.1000 116.1000 83.2000 ;
	    RECT 115.8000 81.1000 116.2000 83.1000 ;
	    RECT 117.4000 81.1000 117.8000 84.8000 ;
	    RECT 118.2000 84.4000 118.6000 84.8000 ;
	    RECT 119.0000 81.1000 119.4000 87.9000 ;
	    RECT 120.6000 87.7000 121.0000 89.9000 ;
	    RECT 122.7000 89.2000 123.3000 89.9000 ;
	    RECT 122.7000 88.9000 123.4000 89.2000 ;
	    RECT 125.0000 88.9000 125.4000 89.9000 ;
	    RECT 127.2000 89.2000 127.6000 89.9000 ;
	    RECT 127.2000 88.9000 128.2000 89.2000 ;
	    RECT 123.0000 88.5000 123.4000 88.9000 ;
	    RECT 125.1000 88.6000 125.4000 88.9000 ;
	    RECT 125.1000 88.3000 126.5000 88.6000 ;
	    RECT 126.1000 88.2000 126.5000 88.3000 ;
	    RECT 127.0000 88.2000 127.4000 88.6000 ;
	    RECT 127.8000 88.5000 128.2000 88.9000 ;
	    RECT 122.1000 87.7000 122.5000 87.8000 ;
	    RECT 119.8000 87.1000 120.2000 87.6000 ;
	    RECT 120.6000 87.4000 122.5000 87.7000 ;
	    RECT 120.6000 87.1000 121.0000 87.4000 ;
	    RECT 124.1000 87.1000 124.5000 87.2000 ;
	    RECT 127.0000 87.1000 127.3000 88.2000 ;
	    RECT 129.4000 87.5000 129.8000 89.9000 ;
	    RECT 131.0000 88.9000 131.4000 89.9000 ;
	    RECT 130.2000 87.8000 130.6000 88.6000 ;
	    RECT 131.1000 87.2000 131.4000 88.9000 ;
	    RECT 131.8000 88.1000 132.2000 88.2000 ;
	    RECT 132.6000 88.1000 133.0000 88.6000 ;
	    RECT 131.8000 87.8000 133.0000 88.1000 ;
	    RECT 133.4000 88.1000 133.8000 89.9000 ;
	    RECT 135.0000 88.9000 135.4000 89.9000 ;
	    RECT 134.2000 88.1000 134.6000 88.6000 ;
	    RECT 133.4000 87.8000 134.6000 88.1000 ;
	    RECT 128.6000 87.1000 129.4000 87.2000 ;
	    RECT 119.8000 86.8000 121.0000 87.1000 ;
	    RECT 120.6000 85.7000 121.0000 86.8000 ;
	    RECT 123.9000 86.8000 129.4000 87.1000 ;
	    RECT 130.2000 86.8000 130.6000 87.2000 ;
	    RECT 131.0000 86.8000 131.4000 87.2000 ;
	    RECT 123.0000 86.4000 123.4000 86.5000 ;
	    RECT 121.5000 86.1000 123.4000 86.4000 ;
	    RECT 123.9000 86.1000 124.2000 86.8000 ;
	    RECT 127.5000 86.7000 127.9000 86.8000 ;
	    RECT 127.0000 86.2000 127.4000 86.3000 ;
	    RECT 128.3000 86.2000 128.7000 86.3000 ;
	    RECT 124.6000 86.1000 125.0000 86.2000 ;
	    RECT 121.5000 86.0000 121.9000 86.1000 ;
	    RECT 123.8000 85.8000 125.0000 86.1000 ;
	    RECT 126.2000 85.9000 128.7000 86.2000 ;
	    RECT 130.2000 86.1000 130.5000 86.8000 ;
	    RECT 131.1000 86.1000 131.4000 86.8000 ;
	    RECT 126.2000 85.8000 126.6000 85.9000 ;
	    RECT 130.2000 85.8000 131.4000 86.1000 ;
	    RECT 122.3000 85.7000 122.7000 85.8000 ;
	    RECT 120.6000 85.4000 122.7000 85.7000 ;
	    RECT 120.6000 81.1000 121.0000 85.4000 ;
	    RECT 123.9000 85.2000 124.2000 85.8000 ;
	    RECT 127.0000 85.5000 129.8000 85.6000 ;
	    RECT 126.9000 85.4000 129.8000 85.5000 ;
	    RECT 123.0000 84.9000 124.2000 85.2000 ;
	    RECT 124.9000 85.3000 129.8000 85.4000 ;
	    RECT 124.9000 85.1000 127.3000 85.3000 ;
	    RECT 123.0000 84.4000 123.3000 84.9000 ;
	    RECT 122.6000 84.0000 123.3000 84.4000 ;
	    RECT 124.1000 84.5000 124.5000 84.6000 ;
	    RECT 124.9000 84.5000 125.2000 85.1000 ;
	    RECT 124.1000 84.2000 125.2000 84.5000 ;
	    RECT 125.5000 84.5000 128.2000 84.8000 ;
	    RECT 125.5000 84.4000 125.9000 84.5000 ;
	    RECT 127.8000 84.4000 128.2000 84.5000 ;
	    RECT 124.7000 83.7000 125.1000 83.8000 ;
	    RECT 126.1000 83.7000 126.5000 83.8000 ;
	    RECT 123.0000 83.1000 123.4000 83.5000 ;
	    RECT 124.7000 83.4000 126.5000 83.7000 ;
	    RECT 125.1000 83.1000 125.4000 83.4000 ;
	    RECT 127.8000 83.1000 128.2000 83.5000 ;
	    RECT 122.7000 81.1000 123.3000 83.1000 ;
	    RECT 125.0000 81.1000 125.4000 83.1000 ;
	    RECT 127.2000 82.8000 128.2000 83.1000 ;
	    RECT 127.2000 81.1000 127.6000 82.8000 ;
	    RECT 129.4000 81.1000 129.8000 85.3000 ;
	    RECT 131.1000 85.1000 131.4000 85.8000 ;
	    RECT 131.8000 85.4000 132.2000 86.2000 ;
	    RECT 131.0000 84.7000 131.9000 85.1000 ;
	    RECT 131.5000 81.1000 131.9000 84.7000 ;
	    RECT 133.4000 81.1000 133.8000 87.8000 ;
	    RECT 135.1000 87.2000 135.4000 88.9000 ;
	    RECT 136.6000 87.5000 137.0000 89.9000 ;
	    RECT 138.8000 89.2000 139.2000 89.9000 ;
	    RECT 138.2000 88.9000 139.2000 89.2000 ;
	    RECT 141.0000 88.9000 141.4000 89.9000 ;
	    RECT 143.1000 89.2000 143.7000 89.9000 ;
	    RECT 143.0000 88.9000 143.7000 89.2000 ;
	    RECT 138.2000 88.5000 138.6000 88.9000 ;
	    RECT 141.0000 88.6000 141.3000 88.9000 ;
	    RECT 139.0000 88.2000 139.4000 88.6000 ;
	    RECT 139.9000 88.3000 141.3000 88.6000 ;
	    RECT 143.0000 88.5000 143.4000 88.9000 ;
	    RECT 139.9000 88.2000 140.3000 88.3000 ;
	    RECT 134.2000 87.1000 134.6000 87.2000 ;
	    RECT 135.0000 87.1000 135.4000 87.2000 ;
	    RECT 134.2000 86.8000 135.4000 87.1000 ;
	    RECT 135.8000 87.1000 136.2000 87.2000 ;
	    RECT 137.0000 87.1000 137.8000 87.2000 ;
	    RECT 139.1000 87.1000 139.4000 88.2000 ;
	    RECT 143.9000 87.7000 144.3000 87.8000 ;
	    RECT 145.4000 87.7000 145.8000 89.9000 ;
	    RECT 143.9000 87.4000 145.8000 87.7000 ;
	    RECT 141.9000 87.1000 142.3000 87.2000 ;
	    RECT 135.8000 86.8000 142.5000 87.1000 ;
	    RECT 135.1000 85.1000 135.4000 86.8000 ;
	    RECT 138.5000 86.7000 138.9000 86.8000 ;
	    RECT 137.7000 86.2000 138.1000 86.3000 ;
	    RECT 139.0000 86.2000 139.4000 86.3000 ;
	    RECT 135.8000 85.4000 136.2000 86.2000 ;
	    RECT 137.7000 85.9000 140.2000 86.2000 ;
	    RECT 139.8000 85.8000 140.2000 85.9000 ;
	    RECT 141.4000 86.1000 141.8000 86.2000 ;
	    RECT 142.2000 86.1000 142.5000 86.8000 ;
	    RECT 143.0000 86.4000 143.4000 86.5000 ;
	    RECT 143.0000 86.1000 144.9000 86.4000 ;
	    RECT 141.4000 85.8000 142.5000 86.1000 ;
	    RECT 144.5000 86.0000 144.9000 86.1000 ;
	    RECT 136.6000 85.5000 139.4000 85.6000 ;
	    RECT 136.6000 85.4000 139.5000 85.5000 ;
	    RECT 136.6000 85.3000 141.5000 85.4000 ;
	    RECT 135.0000 84.7000 135.9000 85.1000 ;
	    RECT 135.5000 81.1000 135.9000 84.7000 ;
	    RECT 136.6000 81.1000 137.0000 85.3000 ;
	    RECT 139.1000 85.1000 141.5000 85.3000 ;
	    RECT 138.2000 84.5000 140.9000 84.8000 ;
	    RECT 138.2000 84.4000 138.6000 84.5000 ;
	    RECT 140.5000 84.4000 140.9000 84.5000 ;
	    RECT 141.2000 84.5000 141.5000 85.1000 ;
	    RECT 142.2000 85.2000 142.5000 85.8000 ;
	    RECT 143.7000 85.7000 144.1000 85.8000 ;
	    RECT 145.4000 85.7000 145.8000 87.4000 ;
	    RECT 143.7000 85.4000 145.8000 85.7000 ;
	    RECT 142.2000 84.9000 143.4000 85.2000 ;
	    RECT 141.9000 84.5000 142.3000 84.6000 ;
	    RECT 141.2000 84.2000 142.3000 84.5000 ;
	    RECT 143.1000 84.4000 143.4000 84.9000 ;
	    RECT 143.1000 84.0000 143.8000 84.4000 ;
	    RECT 139.9000 83.7000 140.3000 83.8000 ;
	    RECT 141.3000 83.7000 141.7000 83.8000 ;
	    RECT 138.2000 83.1000 138.6000 83.5000 ;
	    RECT 139.9000 83.4000 141.7000 83.7000 ;
	    RECT 141.0000 83.1000 141.3000 83.4000 ;
	    RECT 143.0000 83.1000 143.4000 83.5000 ;
	    RECT 138.2000 82.8000 139.2000 83.1000 ;
	    RECT 138.8000 81.1000 139.2000 82.8000 ;
	    RECT 141.0000 81.1000 141.4000 83.1000 ;
	    RECT 143.1000 81.1000 143.7000 83.1000 ;
	    RECT 145.4000 81.1000 145.8000 85.4000 ;
	    RECT 146.2000 87.7000 146.6000 89.9000 ;
	    RECT 148.3000 89.2000 148.9000 89.9000 ;
	    RECT 148.3000 88.9000 149.0000 89.2000 ;
	    RECT 150.6000 88.9000 151.0000 89.9000 ;
	    RECT 152.8000 89.2000 153.2000 89.9000 ;
	    RECT 152.8000 88.9000 153.8000 89.2000 ;
	    RECT 148.6000 88.5000 149.0000 88.9000 ;
	    RECT 150.7000 88.6000 151.0000 88.9000 ;
	    RECT 150.7000 88.3000 152.1000 88.6000 ;
	    RECT 151.7000 88.2000 152.1000 88.3000 ;
	    RECT 152.6000 87.8000 153.0000 88.6000 ;
	    RECT 153.4000 88.5000 153.8000 88.9000 ;
	    RECT 147.7000 87.7000 148.1000 87.8000 ;
	    RECT 146.2000 87.4000 148.1000 87.7000 ;
	    RECT 146.2000 85.7000 146.6000 87.4000 ;
	    RECT 149.7000 87.1000 150.1000 87.2000 ;
	    RECT 152.6000 87.1000 152.9000 87.8000 ;
	    RECT 155.0000 87.5000 155.4000 89.9000 ;
	    RECT 157.1000 89.2000 157.5000 89.9000 ;
	    RECT 157.1000 88.8000 157.8000 89.2000 ;
	    RECT 157.1000 88.2000 157.5000 88.8000 ;
	    RECT 156.6000 87.9000 157.5000 88.2000 ;
	    RECT 158.2000 87.9000 158.6000 89.9000 ;
	    RECT 159.0000 88.0000 159.4000 89.9000 ;
	    RECT 160.6000 88.0000 161.0000 89.9000 ;
	    RECT 163.1000 88.2000 163.5000 88.6000 ;
	    RECT 159.0000 87.9000 161.0000 88.0000 ;
	    RECT 154.2000 87.1000 155.0000 87.2000 ;
	    RECT 149.5000 86.8000 155.0000 87.1000 ;
	    RECT 155.8000 86.8000 156.2000 87.6000 ;
	    RECT 148.6000 86.4000 149.0000 86.5000 ;
	    RECT 147.1000 86.1000 149.0000 86.4000 ;
	    RECT 147.1000 86.0000 147.5000 86.1000 ;
	    RECT 147.9000 85.7000 148.3000 85.8000 ;
	    RECT 146.2000 85.4000 148.3000 85.7000 ;
	    RECT 146.2000 81.1000 146.6000 85.4000 ;
	    RECT 149.5000 85.2000 149.8000 86.8000 ;
	    RECT 153.1000 86.7000 153.5000 86.8000 ;
	    RECT 152.6000 86.2000 153.0000 86.3000 ;
	    RECT 153.9000 86.2000 154.3000 86.3000 ;
	    RECT 151.8000 85.9000 154.3000 86.2000 ;
	    RECT 151.8000 85.8000 152.2000 85.9000 ;
	    RECT 152.6000 85.5000 155.4000 85.6000 ;
	    RECT 152.5000 85.4000 155.4000 85.5000 ;
	    RECT 148.6000 84.9000 149.8000 85.2000 ;
	    RECT 150.5000 85.3000 155.4000 85.4000 ;
	    RECT 150.5000 85.1000 152.9000 85.3000 ;
	    RECT 148.6000 84.4000 148.9000 84.9000 ;
	    RECT 148.2000 84.0000 148.9000 84.4000 ;
	    RECT 149.7000 84.5000 150.1000 84.6000 ;
	    RECT 150.5000 84.5000 150.8000 85.1000 ;
	    RECT 149.7000 84.2000 150.8000 84.5000 ;
	    RECT 151.1000 84.5000 153.8000 84.8000 ;
	    RECT 151.1000 84.4000 151.5000 84.5000 ;
	    RECT 153.4000 84.4000 153.8000 84.5000 ;
	    RECT 150.3000 83.7000 150.7000 83.8000 ;
	    RECT 151.7000 83.7000 152.1000 83.8000 ;
	    RECT 148.6000 83.1000 149.0000 83.5000 ;
	    RECT 150.3000 83.4000 152.1000 83.7000 ;
	    RECT 150.7000 83.1000 151.0000 83.4000 ;
	    RECT 153.4000 83.1000 153.8000 83.5000 ;
	    RECT 148.3000 81.1000 148.9000 83.1000 ;
	    RECT 150.6000 81.1000 151.0000 83.1000 ;
	    RECT 152.8000 82.8000 153.8000 83.1000 ;
	    RECT 152.8000 81.1000 153.2000 82.8000 ;
	    RECT 155.0000 81.1000 155.4000 85.3000 ;
	    RECT 156.6000 81.1000 157.0000 87.9000 ;
	    RECT 158.3000 87.2000 158.6000 87.9000 ;
	    RECT 159.1000 87.7000 160.9000 87.9000 ;
	    RECT 163.0000 87.8000 163.4000 88.2000 ;
	    RECT 163.8000 87.9000 164.2000 89.9000 ;
	    RECT 160.2000 87.2000 160.6000 87.4000 ;
	    RECT 158.2000 86.8000 159.5000 87.2000 ;
	    RECT 160.2000 86.9000 161.0000 87.2000 ;
	    RECT 160.6000 86.8000 161.0000 86.9000 ;
	    RECT 157.4000 85.1000 157.8000 85.2000 ;
	    RECT 158.2000 85.1000 158.6000 85.2000 ;
	    RECT 159.2000 85.1000 159.5000 86.8000 ;
	    RECT 159.8000 85.8000 160.2000 86.6000 ;
	    RECT 161.4000 86.1000 161.8000 86.2000 ;
	    RECT 163.0000 86.1000 163.4000 86.2000 ;
	    RECT 163.9000 86.1000 164.2000 87.9000 ;
	    RECT 166.2000 87.8000 166.6000 88.6000 ;
	    RECT 164.6000 86.4000 165.0000 87.2000 ;
	    RECT 167.0000 87.1000 167.4000 89.9000 ;
	    RECT 169.1000 89.2000 169.5000 89.9000 ;
	    RECT 169.1000 88.8000 169.8000 89.2000 ;
	    RECT 169.1000 88.2000 169.5000 88.8000 ;
	    RECT 168.6000 87.9000 169.5000 88.2000 ;
	    RECT 170.5000 88.2000 170.9000 89.9000 ;
	    RECT 170.5000 87.9000 171.4000 88.2000 ;
	    RECT 167.8000 87.1000 168.2000 87.6000 ;
	    RECT 167.0000 86.8000 168.2000 87.1000 ;
	    RECT 165.4000 86.1000 165.8000 86.2000 ;
	    RECT 161.4000 85.8000 164.2000 86.1000 ;
	    RECT 165.0000 85.8000 165.8000 86.1000 ;
	    RECT 163.1000 85.1000 163.4000 85.8000 ;
	    RECT 165.0000 85.6000 165.4000 85.8000 ;
	    RECT 157.4000 84.8000 158.9000 85.1000 ;
	    RECT 159.2000 84.8000 159.7000 85.1000 ;
	    RECT 157.4000 84.4000 157.8000 84.8000 ;
	    RECT 158.6000 84.2000 158.9000 84.8000 ;
	    RECT 158.6000 83.8000 159.0000 84.2000 ;
	    RECT 159.3000 81.1000 159.7000 84.8000 ;
	    RECT 163.0000 81.1000 163.4000 85.1000 ;
	    RECT 163.8000 84.8000 165.8000 85.1000 ;
	    RECT 163.8000 81.1000 164.2000 84.8000 ;
	    RECT 165.4000 81.1000 165.8000 84.8000 ;
	    RECT 167.0000 81.1000 167.4000 86.8000 ;
	    RECT 168.6000 81.1000 169.0000 87.9000 ;
	    RECT 171.0000 86.1000 171.4000 87.9000 ;
	    RECT 171.8000 86.8000 172.2000 87.6000 ;
	    RECT 172.6000 87.5000 173.0000 89.9000 ;
	    RECT 174.8000 89.2000 175.2000 89.9000 ;
	    RECT 174.2000 88.9000 175.2000 89.2000 ;
	    RECT 177.0000 88.9000 177.4000 89.9000 ;
	    RECT 179.1000 89.2000 179.7000 89.9000 ;
	    RECT 179.0000 88.9000 179.7000 89.2000 ;
	    RECT 174.2000 88.5000 174.6000 88.9000 ;
	    RECT 177.0000 88.6000 177.3000 88.9000 ;
	    RECT 175.0000 87.8000 175.4000 88.6000 ;
	    RECT 175.9000 88.3000 177.3000 88.6000 ;
	    RECT 179.0000 88.5000 179.4000 88.9000 ;
	    RECT 175.9000 88.2000 176.3000 88.3000 ;
	    RECT 173.0000 87.1000 173.8000 87.2000 ;
	    RECT 175.1000 87.1000 175.4000 87.8000 ;
	    RECT 179.9000 87.7000 180.3000 87.8000 ;
	    RECT 181.4000 87.7000 181.8000 89.9000 ;
	    RECT 179.9000 87.4000 181.8000 87.7000 ;
	    RECT 177.9000 87.1000 178.3000 87.2000 ;
	    RECT 173.0000 86.8000 178.5000 87.1000 ;
	    RECT 174.5000 86.7000 174.9000 86.8000 ;
	    RECT 169.4000 85.8000 171.4000 86.1000 ;
	    RECT 173.7000 86.2000 174.1000 86.3000 ;
	    RECT 173.7000 85.9000 176.2000 86.2000 ;
	    RECT 175.8000 85.8000 176.2000 85.9000 ;
	    RECT 169.4000 85.2000 169.7000 85.8000 ;
	    RECT 169.4000 84.4000 169.8000 85.2000 ;
	    RECT 170.2000 84.4000 170.6000 85.2000 ;
	    RECT 171.0000 81.1000 171.4000 85.8000 ;
	    RECT 172.6000 85.5000 175.4000 85.6000 ;
	    RECT 172.6000 85.4000 175.5000 85.5000 ;
	    RECT 172.6000 85.3000 177.5000 85.4000 ;
	    RECT 172.6000 81.1000 173.0000 85.3000 ;
	    RECT 175.1000 85.1000 177.5000 85.3000 ;
	    RECT 174.2000 84.5000 176.9000 84.8000 ;
	    RECT 174.2000 84.4000 174.6000 84.5000 ;
	    RECT 176.5000 84.4000 176.9000 84.5000 ;
	    RECT 177.2000 84.5000 177.5000 85.1000 ;
	    RECT 178.2000 85.2000 178.5000 86.8000 ;
	    RECT 179.0000 86.4000 179.4000 86.5000 ;
	    RECT 179.0000 86.1000 180.9000 86.4000 ;
	    RECT 180.5000 86.0000 180.9000 86.1000 ;
	    RECT 179.7000 85.7000 180.1000 85.8000 ;
	    RECT 181.4000 85.7000 181.8000 87.4000 ;
	    RECT 179.7000 85.4000 181.8000 85.7000 ;
	    RECT 178.2000 84.9000 179.4000 85.2000 ;
	    RECT 177.9000 84.5000 178.3000 84.6000 ;
	    RECT 177.2000 84.2000 178.3000 84.5000 ;
	    RECT 179.1000 84.4000 179.4000 84.9000 ;
	    RECT 179.1000 84.0000 179.8000 84.4000 ;
	    RECT 175.9000 83.7000 176.3000 83.8000 ;
	    RECT 177.3000 83.7000 177.7000 83.8000 ;
	    RECT 174.2000 83.1000 174.6000 83.5000 ;
	    RECT 175.9000 83.4000 177.7000 83.7000 ;
	    RECT 177.0000 83.1000 177.3000 83.4000 ;
	    RECT 179.0000 83.1000 179.4000 83.5000 ;
	    RECT 174.2000 82.8000 175.2000 83.1000 ;
	    RECT 174.8000 81.1000 175.2000 82.8000 ;
	    RECT 177.0000 81.1000 177.4000 83.1000 ;
	    RECT 179.1000 81.1000 179.7000 83.1000 ;
	    RECT 181.4000 81.1000 181.8000 85.4000 ;
	    RECT 182.2000 81.1000 182.6000 89.9000 ;
	    RECT 184.6000 88.9000 185.0000 89.9000 ;
	    RECT 186.5000 89.2000 186.9000 89.9000 ;
	    RECT 183.0000 87.8000 183.4000 88.6000 ;
	    RECT 183.8000 87.8000 184.2000 88.6000 ;
	    RECT 184.7000 87.2000 185.0000 88.9000 ;
	    RECT 186.2000 88.8000 186.9000 89.2000 ;
	    RECT 186.5000 88.2000 186.9000 88.8000 ;
	    RECT 188.7000 88.2000 189.1000 88.6000 ;
	    RECT 186.5000 87.9000 187.4000 88.2000 ;
	    RECT 184.6000 86.8000 185.0000 87.2000 ;
	    RECT 184.7000 85.1000 185.0000 86.8000 ;
	    RECT 185.4000 85.4000 185.8000 86.2000 ;
	    RECT 184.6000 84.7000 185.5000 85.1000 ;
	    RECT 185.1000 84.1000 185.5000 84.7000 ;
	    RECT 186.2000 84.1000 186.6000 85.2000 ;
	    RECT 185.1000 83.8000 186.6000 84.1000 ;
	    RECT 185.1000 81.1000 185.5000 83.8000 ;
	    RECT 187.0000 81.1000 187.4000 87.9000 ;
	    RECT 188.6000 87.8000 189.0000 88.2000 ;
	    RECT 189.4000 87.9000 189.8000 89.9000 ;
	    RECT 187.8000 86.8000 188.2000 87.6000 ;
	    RECT 188.6000 86.1000 189.0000 86.2000 ;
	    RECT 189.5000 86.1000 189.8000 87.9000 ;
	    RECT 192.6000 88.9000 193.0000 89.9000 ;
	    RECT 192.6000 87.2000 192.9000 88.9000 ;
	    RECT 193.4000 87.8000 193.8000 88.6000 ;
	    RECT 190.2000 86.4000 190.6000 87.2000 ;
	    RECT 192.6000 87.1000 193.0000 87.2000 ;
	    RECT 194.8000 87.1000 195.2000 89.9000 ;
	    RECT 191.0000 86.8000 193.0000 87.1000 ;
	    RECT 194.3000 86.9000 195.2000 87.1000 ;
	    RECT 197.4000 87.8000 197.8000 88.6000 ;
	    RECT 197.4000 87.2000 197.7000 87.8000 ;
	    RECT 194.3000 86.8000 195.1000 86.9000 ;
	    RECT 197.4000 86.8000 197.8000 87.2000 ;
	    RECT 191.0000 86.2000 191.3000 86.8000 ;
	    RECT 191.0000 86.1000 191.4000 86.2000 ;
	    RECT 188.6000 85.8000 189.8000 86.1000 ;
	    RECT 190.6000 85.8000 191.4000 86.1000 ;
	    RECT 188.7000 85.1000 189.0000 85.8000 ;
	    RECT 190.6000 85.6000 191.0000 85.8000 ;
	    RECT 191.8000 85.4000 192.2000 86.2000 ;
	    RECT 192.6000 85.1000 192.9000 86.8000 ;
	    RECT 194.3000 85.2000 194.6000 86.8000 ;
	    RECT 195.4000 85.8000 196.2000 86.2000 ;
	    RECT 188.6000 81.1000 189.0000 85.1000 ;
	    RECT 189.4000 84.8000 191.4000 85.1000 ;
	    RECT 189.4000 81.1000 189.8000 84.8000 ;
	    RECT 191.0000 81.1000 191.4000 84.8000 ;
	    RECT 192.1000 84.7000 193.0000 85.1000 ;
	    RECT 194.2000 84.8000 194.6000 85.2000 ;
	    RECT 196.6000 84.8000 197.0000 85.6000 ;
	    RECT 192.1000 81.1000 192.5000 84.7000 ;
	    RECT 194.3000 83.5000 194.6000 84.8000 ;
	    RECT 195.0000 83.8000 195.4000 84.6000 ;
	    RECT 194.3000 83.2000 196.1000 83.5000 ;
	    RECT 194.3000 83.1000 194.6000 83.2000 ;
	    RECT 194.2000 81.1000 194.6000 83.1000 ;
	    RECT 195.8000 81.1000 196.2000 83.2000 ;
	    RECT 198.2000 81.1000 198.6000 89.9000 ;
	    RECT 199.8000 88.9000 200.2000 89.9000 ;
	    RECT 199.8000 87.2000 200.1000 88.9000 ;
	    RECT 200.6000 87.8000 201.0000 88.6000 ;
	    RECT 201.4000 88.0000 201.8000 89.9000 ;
	    RECT 203.0000 88.0000 203.4000 89.9000 ;
	    RECT 201.4000 87.9000 203.4000 88.0000 ;
	    RECT 203.8000 87.9000 204.2000 89.9000 ;
	    RECT 204.9000 88.2000 205.3000 89.9000 ;
	    RECT 207.8000 88.9000 208.2000 89.9000 ;
	    RECT 204.9000 87.9000 205.8000 88.2000 ;
	    RECT 201.5000 87.7000 203.3000 87.9000 ;
	    RECT 201.8000 87.2000 202.2000 87.4000 ;
	    RECT 203.8000 87.2000 204.1000 87.9000 ;
	    RECT 199.8000 86.8000 200.2000 87.2000 ;
	    RECT 201.4000 86.9000 202.2000 87.2000 ;
	    RECT 201.4000 86.8000 201.8000 86.9000 ;
	    RECT 202.9000 86.8000 204.2000 87.2000 ;
	    RECT 199.0000 85.4000 199.4000 86.2000 ;
	    RECT 199.8000 85.2000 200.1000 86.8000 ;
	    RECT 200.6000 86.1000 201.0000 86.2000 ;
	    RECT 202.2000 86.1000 202.6000 86.6000 ;
	    RECT 200.6000 85.8000 202.6000 86.1000 ;
	    RECT 202.9000 86.2000 203.2000 86.8000 ;
	    RECT 202.9000 85.8000 203.4000 86.2000 ;
	    RECT 199.8000 85.1000 200.2000 85.2000 ;
	    RECT 202.9000 85.1000 203.2000 85.8000 ;
	    RECT 203.8000 85.1000 204.2000 85.2000 ;
	    RECT 199.3000 84.7000 200.2000 85.1000 ;
	    RECT 202.7000 84.8000 203.2000 85.1000 ;
	    RECT 203.5000 84.8000 204.2000 85.1000 ;
	    RECT 199.3000 81.1000 199.7000 84.7000 ;
	    RECT 202.7000 81.1000 203.1000 84.8000 ;
	    RECT 203.5000 84.2000 203.8000 84.8000 ;
	    RECT 204.6000 84.4000 205.0000 85.2000 ;
	    RECT 203.4000 83.8000 203.8000 84.2000 ;
	    RECT 205.4000 81.1000 205.8000 87.9000 ;
	    RECT 207.0000 87.8000 207.4000 88.6000 ;
	    RECT 206.2000 86.8000 206.6000 87.6000 ;
	    RECT 207.9000 87.2000 208.2000 88.9000 ;
	    RECT 208.6000 88.1000 209.0000 88.2000 ;
	    RECT 209.4000 88.1000 209.8000 88.6000 ;
	    RECT 208.6000 87.8000 209.8000 88.1000 ;
	    RECT 207.8000 86.8000 208.2000 87.2000 ;
	    RECT 207.0000 86.1000 207.4000 86.2000 ;
	    RECT 207.9000 86.1000 208.2000 86.8000 ;
	    RECT 210.2000 87.1000 210.6000 89.9000 ;
	    RECT 212.6000 88.0000 213.0000 89.9000 ;
	    RECT 214.2000 88.0000 214.6000 89.9000 ;
	    RECT 212.6000 87.9000 214.6000 88.0000 ;
	    RECT 215.0000 87.9000 215.4000 89.9000 ;
	    RECT 215.8000 87.9000 216.2000 89.9000 ;
	    RECT 216.6000 88.0000 217.0000 89.9000 ;
	    RECT 218.2000 88.0000 218.6000 89.9000 ;
	    RECT 219.1000 88.2000 219.5000 88.6000 ;
	    RECT 216.6000 87.9000 218.6000 88.0000 ;
	    RECT 212.7000 87.7000 214.5000 87.9000 ;
	    RECT 213.0000 87.2000 213.4000 87.4000 ;
	    RECT 215.0000 87.2000 215.3000 87.9000 ;
	    RECT 215.9000 87.2000 216.2000 87.9000 ;
	    RECT 216.7000 87.7000 218.5000 87.9000 ;
	    RECT 219.0000 87.8000 219.4000 88.2000 ;
	    RECT 219.8000 87.9000 220.2000 89.9000 ;
	    RECT 222.2000 88.0000 222.6000 89.9000 ;
	    RECT 223.8000 88.0000 224.2000 89.9000 ;
	    RECT 222.2000 87.9000 224.2000 88.0000 ;
	    RECT 217.8000 87.2000 218.2000 87.4000 ;
	    RECT 212.6000 87.1000 213.4000 87.2000 ;
	    RECT 210.2000 86.9000 213.4000 87.1000 ;
	    RECT 210.2000 86.8000 213.0000 86.9000 ;
	    RECT 214.1000 86.8000 215.4000 87.2000 ;
	    RECT 215.8000 86.8000 217.1000 87.2000 ;
	    RECT 217.8000 87.1000 218.6000 87.2000 ;
	    RECT 219.9000 87.1000 220.2000 87.9000 ;
	    RECT 222.3000 87.7000 224.1000 87.9000 ;
	    RECT 224.6000 87.8000 225.0000 89.9000 ;
	    RECT 225.4000 88.0000 225.8000 89.9000 ;
	    RECT 227.0000 88.0000 227.4000 89.9000 ;
	    RECT 225.4000 87.9000 227.4000 88.0000 ;
	    RECT 227.8000 87.9000 228.2000 89.9000 ;
	    RECT 222.6000 87.2000 223.0000 87.4000 ;
	    RECT 224.6000 87.2000 224.9000 87.8000 ;
	    RECT 225.5000 87.7000 227.3000 87.9000 ;
	    RECT 225.8000 87.2000 226.2000 87.4000 ;
	    RECT 227.8000 87.2000 228.1000 87.9000 ;
	    RECT 217.8000 86.9000 220.2000 87.1000 ;
	    RECT 218.2000 86.8000 220.2000 86.9000 ;
	    RECT 207.0000 85.8000 208.2000 86.1000 ;
	    RECT 207.9000 85.1000 208.2000 85.8000 ;
	    RECT 208.6000 86.1000 209.0000 86.2000 ;
	    RECT 209.4000 86.1000 209.8000 86.2000 ;
	    RECT 208.6000 85.8000 209.8000 86.1000 ;
	    RECT 208.6000 85.4000 209.0000 85.8000 ;
	    RECT 207.8000 84.7000 208.7000 85.1000 ;
	    RECT 208.3000 81.1000 208.7000 84.7000 ;
	    RECT 210.2000 81.1000 210.6000 86.8000 ;
	    RECT 213.4000 85.8000 213.8000 86.6000 ;
	    RECT 214.1000 86.1000 214.4000 86.8000 ;
	    RECT 214.1000 85.8000 216.1000 86.1000 ;
	    RECT 214.1000 85.1000 214.4000 85.8000 ;
	    RECT 215.8000 85.2000 216.1000 85.8000 ;
	    RECT 215.0000 85.1000 215.4000 85.2000 ;
	    RECT 213.9000 84.8000 214.4000 85.1000 ;
	    RECT 214.7000 84.8000 215.4000 85.1000 ;
	    RECT 215.8000 85.1000 216.2000 85.2000 ;
	    RECT 216.8000 85.1000 217.1000 86.8000 ;
	    RECT 217.4000 85.8000 217.8000 86.6000 ;
	    RECT 219.0000 86.1000 219.4000 86.2000 ;
	    RECT 219.9000 86.1000 220.2000 86.8000 ;
	    RECT 220.6000 87.1000 221.0000 87.2000 ;
	    RECT 221.4000 87.1000 221.8000 87.2000 ;
	    RECT 220.6000 86.8000 221.8000 87.1000 ;
	    RECT 222.2000 86.9000 223.0000 87.2000 ;
	    RECT 222.2000 86.8000 222.6000 86.9000 ;
	    RECT 223.7000 86.8000 225.0000 87.2000 ;
	    RECT 225.4000 86.9000 226.2000 87.2000 ;
	    RECT 225.4000 86.8000 225.8000 86.9000 ;
	    RECT 226.9000 86.8000 228.2000 87.2000 ;
	    RECT 220.6000 86.4000 221.0000 86.8000 ;
	    RECT 221.4000 86.1000 221.8000 86.2000 ;
	    RECT 222.2000 86.1000 222.6000 86.2000 ;
	    RECT 219.0000 85.8000 220.2000 86.1000 ;
	    RECT 221.0000 85.8000 222.6000 86.1000 ;
	    RECT 223.0000 85.8000 223.4000 86.6000 ;
	    RECT 219.1000 85.1000 219.4000 85.8000 ;
	    RECT 221.0000 85.6000 221.4000 85.8000 ;
	    RECT 223.7000 85.1000 224.0000 86.8000 ;
	    RECT 225.4000 86.1000 225.7000 86.8000 ;
	    RECT 224.6000 85.8000 225.7000 86.1000 ;
	    RECT 226.2000 85.8000 226.6000 86.6000 ;
	    RECT 224.6000 85.2000 224.9000 85.8000 ;
	    RECT 224.6000 85.1000 225.0000 85.2000 ;
	    RECT 226.9000 85.1000 227.2000 86.8000 ;
	    RECT 227.8000 85.1000 228.2000 85.2000 ;
	    RECT 228.6000 85.1000 229.0000 89.9000 ;
	    RECT 229.4000 87.8000 229.8000 88.6000 ;
	    RECT 215.8000 84.8000 216.5000 85.1000 ;
	    RECT 216.8000 84.8000 217.3000 85.1000 ;
	    RECT 213.9000 81.1000 214.3000 84.8000 ;
	    RECT 214.7000 84.2000 215.0000 84.8000 ;
	    RECT 214.6000 83.8000 215.0000 84.2000 ;
	    RECT 216.2000 84.2000 216.5000 84.8000 ;
	    RECT 216.2000 83.8000 216.6000 84.2000 ;
	    RECT 216.9000 82.2000 217.3000 84.8000 ;
	    RECT 216.9000 81.8000 217.8000 82.2000 ;
	    RECT 216.9000 81.1000 217.3000 81.8000 ;
	    RECT 219.0000 81.1000 219.4000 85.1000 ;
	    RECT 219.8000 84.8000 221.8000 85.1000 ;
	    RECT 219.8000 81.1000 220.2000 84.8000 ;
	    RECT 221.4000 81.1000 221.8000 84.8000 ;
	    RECT 223.5000 84.8000 224.0000 85.1000 ;
	    RECT 224.3000 84.8000 225.0000 85.1000 ;
	    RECT 226.7000 84.8000 227.2000 85.1000 ;
	    RECT 227.5000 84.8000 229.0000 85.1000 ;
	    RECT 223.5000 81.1000 223.9000 84.8000 ;
	    RECT 224.3000 84.2000 224.6000 84.8000 ;
	    RECT 224.2000 83.8000 224.6000 84.2000 ;
	    RECT 226.7000 81.1000 227.1000 84.8000 ;
	    RECT 227.5000 84.2000 227.8000 84.8000 ;
	    RECT 227.4000 83.8000 227.8000 84.2000 ;
	    RECT 228.6000 81.1000 229.0000 84.8000 ;
	    RECT 229.4000 84.1000 229.8000 84.2000 ;
	    RECT 230.2000 84.1000 230.6000 89.9000 ;
	    RECT 231.0000 87.8000 231.4000 88.6000 ;
	    RECT 231.8000 87.9000 232.2000 89.9000 ;
	    RECT 234.0000 88.1000 234.8000 89.9000 ;
	    RECT 231.8000 87.6000 233.1000 87.9000 ;
	    RECT 232.7000 87.5000 233.1000 87.6000 ;
	    RECT 233.4000 87.4000 234.2000 87.8000 ;
	    RECT 231.8000 87.1000 232.6000 87.2000 ;
	    RECT 234.5000 87.1000 234.8000 88.1000 ;
	    RECT 236.6000 87.9000 237.0000 89.9000 ;
	    RECT 235.1000 87.4000 235.5000 87.8000 ;
	    RECT 235.8000 87.6000 237.0000 87.9000 ;
	    RECT 237.4000 87.8000 237.8000 88.6000 ;
	    RECT 235.8000 87.5000 236.2000 87.6000 ;
	    RECT 231.8000 87.0000 232.9000 87.1000 ;
	    RECT 231.8000 86.8000 234.0000 87.0000 ;
	    RECT 232.6000 86.7000 234.0000 86.8000 ;
	    RECT 233.6000 86.6000 234.0000 86.7000 ;
	    RECT 234.3000 86.8000 234.8000 87.1000 ;
	    RECT 235.2000 87.2000 235.5000 87.4000 ;
	    RECT 235.2000 86.8000 235.6000 87.2000 ;
	    RECT 234.3000 86.2000 234.6000 86.8000 ;
	    RECT 232.9000 86.1000 233.3000 86.2000 ;
	    RECT 234.2000 86.1000 234.6000 86.2000 ;
	    RECT 235.0000 86.1000 235.4000 86.2000 ;
	    RECT 232.9000 85.8000 233.7000 86.1000 ;
	    RECT 234.2000 85.8000 235.4000 86.1000 ;
	    RECT 238.2000 86.1000 238.6000 89.9000 ;
	    RECT 239.0000 86.8000 239.4000 87.2000 ;
	    RECT 239.0000 86.1000 239.3000 86.8000 ;
	    RECT 238.2000 85.8000 239.3000 86.1000 ;
	    RECT 233.3000 85.7000 233.7000 85.8000 ;
	    RECT 234.3000 85.1000 234.6000 85.8000 ;
	    RECT 229.4000 83.8000 230.6000 84.1000 ;
	    RECT 230.2000 81.1000 230.6000 83.8000 ;
	    RECT 231.8000 84.8000 233.1000 85.1000 ;
	    RECT 231.8000 81.1000 232.2000 84.8000 ;
	    RECT 232.7000 84.7000 233.1000 84.8000 ;
	    RECT 234.0000 81.1000 234.8000 85.1000 ;
	    RECT 235.8000 84.8000 237.0000 85.1000 ;
	    RECT 235.8000 84.7000 236.2000 84.8000 ;
	    RECT 236.6000 81.1000 237.0000 84.8000 ;
	    RECT 238.2000 81.1000 238.6000 85.8000 ;
	    RECT 239.8000 81.1000 240.2000 89.9000 ;
	    RECT 241.4000 87.8000 241.8000 88.6000 ;
	    RECT 240.6000 86.8000 241.0000 87.6000 ;
	    RECT 242.2000 86.1000 242.6000 89.9000 ;
	    RECT 243.0000 88.0000 243.4000 89.9000 ;
	    RECT 244.6000 88.0000 245.0000 89.9000 ;
	    RECT 243.0000 87.9000 245.0000 88.0000 ;
	    RECT 245.4000 87.9000 245.8000 89.9000 ;
	    RECT 246.2000 88.0000 246.6000 89.9000 ;
	    RECT 247.8000 88.0000 248.2000 89.9000 ;
	    RECT 246.2000 87.9000 248.2000 88.0000 ;
	    RECT 248.6000 87.9000 249.0000 89.9000 ;
	    RECT 250.2000 88.9000 250.6000 89.9000 ;
	    RECT 243.1000 87.7000 244.9000 87.9000 ;
	    RECT 243.4000 87.2000 243.8000 87.4000 ;
	    RECT 245.4000 87.2000 245.7000 87.9000 ;
	    RECT 246.3000 87.7000 248.1000 87.9000 ;
	    RECT 246.6000 87.2000 247.0000 87.4000 ;
	    RECT 248.6000 87.2000 248.9000 87.9000 ;
	    RECT 250.2000 87.2000 250.5000 88.9000 ;
	    RECT 251.0000 87.8000 251.4000 88.6000 ;
	    RECT 251.8000 88.0000 252.2000 89.9000 ;
	    RECT 253.4000 88.0000 253.8000 89.9000 ;
	    RECT 251.8000 87.9000 253.8000 88.0000 ;
	    RECT 254.2000 87.9000 254.6000 89.9000 ;
	    RECT 255.0000 88.0000 255.4000 89.9000 ;
	    RECT 256.6000 88.0000 257.0000 89.9000 ;
	    RECT 255.0000 87.9000 257.0000 88.0000 ;
	    RECT 257.4000 87.9000 257.8000 89.9000 ;
	    RECT 258.2000 87.9000 258.6000 89.9000 ;
	    RECT 260.4000 89.2000 261.2000 89.9000 ;
	    RECT 259.8000 88.8000 261.2000 89.2000 ;
	    RECT 260.4000 88.1000 261.2000 88.8000 ;
	    RECT 251.9000 87.7000 253.7000 87.9000 ;
	    RECT 252.2000 87.2000 252.6000 87.4000 ;
	    RECT 254.2000 87.2000 254.5000 87.9000 ;
	    RECT 255.1000 87.7000 256.9000 87.9000 ;
	    RECT 255.4000 87.2000 255.8000 87.4000 ;
	    RECT 257.4000 87.2000 257.7000 87.9000 ;
	    RECT 258.2000 87.6000 259.5000 87.9000 ;
	    RECT 259.1000 87.5000 259.5000 87.6000 ;
	    RECT 259.8000 87.4000 260.6000 87.8000 ;
	    RECT 243.0000 86.9000 243.8000 87.2000 ;
	    RECT 244.5000 87.1000 245.8000 87.2000 ;
	    RECT 246.2000 87.1000 247.0000 87.2000 ;
	    RECT 244.5000 86.9000 247.0000 87.1000 ;
	    RECT 243.0000 86.8000 243.4000 86.9000 ;
	    RECT 244.5000 86.8000 246.6000 86.9000 ;
	    RECT 247.7000 86.8000 249.0000 87.2000 ;
	    RECT 250.2000 87.1000 250.6000 87.2000 ;
	    RECT 251.8000 87.1000 252.6000 87.2000 ;
	    RECT 250.2000 86.9000 252.6000 87.1000 ;
	    RECT 250.2000 86.8000 252.2000 86.9000 ;
	    RECT 253.3000 86.8000 254.6000 87.2000 ;
	    RECT 255.0000 86.9000 255.8000 87.2000 ;
	    RECT 255.0000 86.8000 255.4000 86.9000 ;
	    RECT 256.5000 86.8000 257.8000 87.2000 ;
	    RECT 260.9000 87.1000 261.2000 88.1000 ;
	    RECT 263.0000 87.9000 263.4000 89.9000 ;
	    RECT 261.5000 87.4000 261.9000 87.8000 ;
	    RECT 262.2000 87.6000 263.4000 87.9000 ;
	    RECT 263.8000 87.9000 264.2000 89.9000 ;
	    RECT 266.0000 89.2000 266.8000 89.9000 ;
	    RECT 265.4000 88.8000 266.8000 89.2000 ;
	    RECT 266.0000 88.1000 266.8000 88.8000 ;
	    RECT 263.8000 87.6000 265.0000 87.9000 ;
	    RECT 262.2000 87.5000 262.6000 87.6000 ;
	    RECT 264.6000 87.5000 265.0000 87.6000 ;
	    RECT 260.7000 86.8000 261.2000 87.1000 ;
	    RECT 261.6000 87.2000 261.9000 87.4000 ;
	    RECT 265.3000 87.4000 265.7000 87.8000 ;
	    RECT 265.3000 87.2000 265.6000 87.4000 ;
	    RECT 261.6000 86.8000 262.0000 87.2000 ;
	    RECT 265.2000 86.8000 265.6000 87.2000 ;
	    RECT 243.8000 86.1000 244.2000 86.6000 ;
	    RECT 242.2000 85.8000 244.2000 86.1000 ;
	    RECT 242.2000 81.1000 242.6000 85.8000 ;
	    RECT 244.5000 85.1000 244.8000 86.8000 ;
	    RECT 245.4000 86.1000 245.8000 86.2000 ;
	    RECT 247.0000 86.1000 247.4000 86.6000 ;
	    RECT 245.4000 85.8000 247.4000 86.1000 ;
	    RECT 247.7000 86.1000 248.0000 86.8000 ;
	    RECT 249.4000 86.1000 249.8000 86.2000 ;
	    RECT 247.7000 85.8000 249.8000 86.1000 ;
	    RECT 245.4000 85.1000 245.8000 85.2000 ;
	    RECT 247.7000 85.1000 248.0000 85.8000 ;
	    RECT 249.4000 85.4000 249.8000 85.8000 ;
	    RECT 248.6000 85.1000 249.0000 85.2000 ;
	    RECT 250.2000 85.1000 250.5000 86.8000 ;
	    RECT 252.6000 85.8000 253.0000 86.6000 ;
	    RECT 253.3000 85.1000 253.6000 86.8000 ;
	    RECT 255.8000 85.8000 256.2000 86.6000 ;
	    RECT 256.5000 86.1000 256.8000 86.8000 ;
	    RECT 260.7000 86.2000 261.0000 86.8000 ;
	    RECT 266.0000 86.4000 266.3000 88.1000 ;
	    RECT 268.6000 87.9000 269.0000 89.9000 ;
	    RECT 266.6000 87.7000 267.4000 87.8000 ;
	    RECT 266.6000 87.4000 267.6000 87.7000 ;
	    RECT 267.9000 87.6000 269.0000 87.9000 ;
	    RECT 267.9000 87.5000 268.3000 87.6000 ;
	    RECT 267.3000 87.2000 267.6000 87.4000 ;
	    RECT 266.6000 86.7000 267.0000 87.1000 ;
	    RECT 267.3000 86.9000 269.0000 87.2000 ;
	    RECT 268.2000 86.8000 269.0000 86.9000 ;
	    RECT 265.8000 86.2000 266.3000 86.4000 ;
	    RECT 257.4000 86.1000 257.8000 86.2000 ;
	    RECT 256.5000 85.8000 257.8000 86.1000 ;
	    RECT 259.3000 86.1000 259.7000 86.2000 ;
	    RECT 259.3000 85.8000 260.1000 86.1000 ;
	    RECT 260.6000 85.8000 261.0000 86.2000 ;
	    RECT 265.4000 86.1000 266.3000 86.2000 ;
	    RECT 266.7000 86.4000 267.0000 86.7000 ;
	    RECT 266.7000 86.1000 268.0000 86.4000 ;
	    RECT 265.4000 85.8000 266.1000 86.1000 ;
	    RECT 267.6000 86.0000 268.0000 86.1000 ;
	    RECT 254.2000 85.1000 254.6000 85.2000 ;
	    RECT 256.5000 85.1000 256.8000 85.8000 ;
	    RECT 259.7000 85.7000 260.1000 85.8000 ;
	    RECT 257.4000 85.1000 257.8000 85.2000 ;
	    RECT 260.7000 85.1000 261.0000 85.8000 ;
	    RECT 265.8000 85.1000 266.1000 85.8000 ;
	    RECT 266.5000 85.7000 266.9000 85.8000 ;
	    RECT 266.5000 85.4000 268.2000 85.7000 ;
	    RECT 267.9000 85.1000 268.2000 85.4000 ;
	    RECT 244.3000 84.8000 244.8000 85.1000 ;
	    RECT 245.1000 84.8000 245.8000 85.1000 ;
	    RECT 247.5000 84.8000 248.0000 85.1000 ;
	    RECT 248.3000 84.8000 249.0000 85.1000 ;
	    RECT 244.3000 81.1000 244.7000 84.8000 ;
	    RECT 245.1000 84.2000 245.4000 84.8000 ;
	    RECT 245.0000 83.8000 245.4000 84.2000 ;
	    RECT 247.5000 81.1000 247.9000 84.8000 ;
	    RECT 248.3000 84.2000 248.6000 84.8000 ;
	    RECT 248.2000 83.8000 248.6000 84.2000 ;
	    RECT 249.7000 84.7000 250.6000 85.1000 ;
	    RECT 253.1000 84.8000 253.6000 85.1000 ;
	    RECT 253.9000 84.8000 254.6000 85.1000 ;
	    RECT 256.3000 84.8000 256.8000 85.1000 ;
	    RECT 257.1000 84.8000 257.8000 85.1000 ;
	    RECT 258.2000 84.8000 259.5000 85.1000 ;
	    RECT 249.7000 81.1000 250.1000 84.7000 ;
	    RECT 253.1000 81.1000 253.5000 84.8000 ;
	    RECT 253.9000 84.2000 254.2000 84.8000 ;
	    RECT 253.8000 83.8000 254.2000 84.2000 ;
	    RECT 256.3000 81.1000 256.7000 84.8000 ;
	    RECT 257.1000 84.2000 257.4000 84.8000 ;
	    RECT 257.0000 83.8000 257.4000 84.2000 ;
	    RECT 258.2000 81.1000 258.6000 84.8000 ;
	    RECT 259.1000 84.7000 259.5000 84.8000 ;
	    RECT 260.4000 81.1000 261.2000 85.1000 ;
	    RECT 262.2000 84.8000 263.4000 85.1000 ;
	    RECT 262.2000 84.7000 262.6000 84.8000 ;
	    RECT 263.0000 81.1000 263.4000 84.8000 ;
	    RECT 263.8000 84.8000 265.0000 85.1000 ;
	    RECT 265.8000 84.8000 266.8000 85.1000 ;
	    RECT 263.8000 81.1000 264.2000 84.8000 ;
	    RECT 264.6000 84.7000 265.0000 84.8000 ;
	    RECT 266.0000 81.1000 266.8000 84.8000 ;
	    RECT 267.9000 84.8000 269.0000 85.1000 ;
	    RECT 267.9000 84.7000 268.3000 84.8000 ;
	    RECT 268.6000 81.1000 269.0000 84.8000 ;
	    RECT 1.4000 75.1000 1.8000 79.9000 ;
	    RECT 2.2000 79.6000 4.2000 79.9000 ;
	    RECT 2.2000 75.9000 2.6000 79.6000 ;
	    RECT 3.0000 75.9000 3.4000 79.3000 ;
	    RECT 3.8000 76.2000 4.2000 79.6000 ;
	    RECT 5.4000 76.2000 5.8000 79.9000 ;
	    RECT 3.8000 75.9000 5.8000 76.2000 ;
	    RECT 7.5000 78.2000 8.5000 79.9000 ;
	    RECT 7.5000 77.8000 9.0000 78.2000 ;
	    RECT 7.5000 75.9000 8.5000 77.8000 ;
	    RECT 3.1000 75.6000 3.4000 75.9000 ;
	    RECT 2.2000 75.1000 2.6000 75.6000 ;
	    RECT 3.1000 75.3000 4.1000 75.6000 ;
	    RECT 1.4000 74.8000 2.6000 75.1000 ;
	    RECT 3.8000 75.2000 4.1000 75.3000 ;
	    RECT 5.0000 75.2000 5.4000 75.4000 ;
	    RECT 3.8000 74.8000 4.2000 75.2000 ;
	    RECT 5.0000 74.9000 5.8000 75.2000 ;
	    RECT 5.4000 74.8000 5.8000 74.9000 ;
	    RECT 1.4000 71.1000 1.8000 74.8000 ;
	    RECT 3.8000 73.1000 4.1000 74.8000 ;
	    RECT 6.2000 73.8000 6.6000 74.6000 ;
	    RECT 7.9000 74.2000 8.2000 75.9000 ;
	    RECT 7.8000 74.1000 8.2000 74.2000 ;
	    RECT 9.4000 74.1000 9.8000 74.2000 ;
	    RECT 10.2000 74.1000 10.6000 79.9000 ;
	    RECT 7.0000 73.8000 8.2000 74.1000 ;
	    RECT 9.0000 73.8000 10.6000 74.1000 ;
	    RECT 7.0000 73.1000 7.3000 73.8000 ;
	    RECT 9.0000 73.6000 9.4000 73.8000 ;
	    RECT 7.9000 73.1000 9.7000 73.3000 ;
	    RECT 3.5000 71.1000 4.3000 73.1000 ;
	    RECT 6.2000 71.4000 6.6000 73.1000 ;
	    RECT 7.0000 71.7000 7.4000 73.1000 ;
	    RECT 7.8000 73.0000 9.8000 73.1000 ;
	    RECT 7.8000 71.4000 8.2000 73.0000 ;
	    RECT 6.2000 71.1000 8.2000 71.4000 ;
	    RECT 9.4000 71.1000 9.8000 73.0000 ;
	    RECT 10.2000 71.1000 10.6000 73.8000 ;
	    RECT 12.6000 74.1000 13.0000 79.9000 ;
	    RECT 13.4000 79.6000 15.4000 79.9000 ;
	    RECT 13.4000 75.9000 13.8000 79.6000 ;
	    RECT 14.2000 75.9000 14.6000 79.3000 ;
	    RECT 15.0000 76.2000 15.4000 79.6000 ;
	    RECT 16.6000 76.2000 17.0000 79.9000 ;
	    RECT 17.8000 76.8000 18.2000 77.2000 ;
	    RECT 17.8000 76.2000 18.1000 76.8000 ;
	    RECT 18.5000 76.2000 18.9000 79.9000 ;
	    RECT 15.0000 75.9000 17.0000 76.2000 ;
	    RECT 17.4000 75.9000 18.1000 76.2000 ;
	    RECT 18.4000 75.9000 18.9000 76.2000 ;
	    RECT 20.6000 76.1000 21.0000 79.9000 ;
	    RECT 21.4000 76.1000 21.8000 76.2000 ;
	    RECT 14.3000 75.6000 14.6000 75.9000 ;
	    RECT 17.4000 75.8000 17.8000 75.9000 ;
	    RECT 14.3000 75.3000 15.3000 75.6000 ;
	    RECT 15.0000 75.2000 15.3000 75.3000 ;
	    RECT 16.2000 75.2000 16.6000 75.4000 ;
	    RECT 15.0000 74.8000 15.4000 75.2000 ;
	    RECT 16.2000 74.9000 17.0000 75.2000 ;
	    RECT 16.6000 74.8000 17.0000 74.9000 ;
	    RECT 14.3000 74.4000 14.7000 74.8000 ;
	    RECT 14.3000 74.2000 14.6000 74.4000 ;
	    RECT 14.2000 74.1000 14.6000 74.2000 ;
	    RECT 12.6000 73.8000 14.6000 74.1000 ;
	    RECT 12.6000 71.1000 13.0000 73.8000 ;
	    RECT 15.0000 73.2000 15.3000 74.8000 ;
	    RECT 18.4000 74.2000 18.7000 75.9000 ;
	    RECT 20.6000 75.8000 21.8000 76.1000 ;
	    RECT 17.4000 73.8000 18.7000 74.2000 ;
	    RECT 19.8000 74.1000 20.2000 74.2000 ;
	    RECT 20.6000 74.1000 21.0000 75.8000 ;
	    RECT 19.4000 73.8000 21.0000 74.1000 ;
	    RECT 15.0000 73.1000 15.4000 73.2000 ;
	    RECT 17.5000 73.1000 17.8000 73.8000 ;
	    RECT 19.4000 73.6000 19.8000 73.8000 ;
	    RECT 18.3000 73.1000 20.1000 73.3000 ;
	    RECT 14.7000 71.1000 15.5000 73.1000 ;
	    RECT 17.4000 71.1000 17.8000 73.1000 ;
	    RECT 18.2000 73.0000 20.2000 73.1000 ;
	    RECT 18.2000 71.1000 18.6000 73.0000 ;
	    RECT 19.8000 71.1000 20.2000 73.0000 ;
	    RECT 20.6000 71.1000 21.0000 73.8000 ;
	    RECT 22.2000 73.4000 22.6000 74.2000 ;
	    RECT 23.0000 73.1000 23.4000 79.9000 ;
	    RECT 25.4000 77.9000 25.8000 79.9000 ;
	    RECT 23.8000 75.8000 24.2000 76.6000 ;
	    RECT 25.5000 75.8000 25.8000 77.9000 ;
	    RECT 27.0000 75.8000 27.4000 79.9000 ;
	    RECT 29.1000 76.2000 29.5000 79.9000 ;
	    RECT 29.8000 76.8000 30.2000 77.2000 ;
	    RECT 29.9000 76.2000 30.2000 76.8000 ;
	    RECT 29.1000 75.9000 29.6000 76.2000 ;
	    RECT 29.9000 75.9000 30.6000 76.2000 ;
	    RECT 25.5000 75.5000 26.7000 75.8000 ;
	    RECT 25.4000 74.8000 25.8000 75.2000 ;
	    RECT 24.6000 73.8000 25.0000 74.6000 ;
	    RECT 25.5000 74.4000 25.8000 74.8000 ;
	    RECT 25.5000 74.1000 26.0000 74.4000 ;
	    RECT 25.6000 74.0000 26.0000 74.1000 ;
	    RECT 26.4000 73.8000 26.7000 75.5000 ;
	    RECT 27.1000 75.2000 27.4000 75.8000 ;
	    RECT 27.0000 74.8000 27.4000 75.2000 ;
	    RECT 26.4000 73.7000 26.8000 73.8000 ;
	    RECT 25.3000 73.5000 26.8000 73.7000 ;
	    RECT 24.7000 73.4000 26.8000 73.5000 ;
	    RECT 24.7000 73.2000 25.6000 73.4000 ;
	    RECT 24.7000 73.1000 25.0000 73.2000 ;
	    RECT 27.1000 73.1000 27.4000 74.8000 ;
	    RECT 28.6000 74.4000 29.0000 75.2000 ;
	    RECT 29.3000 74.2000 29.6000 75.9000 ;
	    RECT 30.2000 75.8000 30.6000 75.9000 ;
	    RECT 31.0000 75.8000 31.4000 76.6000 ;
	    RECT 27.8000 74.1000 28.2000 74.2000 ;
	    RECT 27.8000 73.8000 28.6000 74.1000 ;
	    RECT 29.3000 73.8000 30.6000 74.2000 ;
	    RECT 28.2000 73.6000 28.6000 73.8000 ;
	    RECT 27.9000 73.1000 29.7000 73.3000 ;
	    RECT 30.2000 73.1000 30.5000 73.8000 ;
	    RECT 31.8000 73.1000 32.2000 79.9000 ;
	    RECT 34.7000 76.3000 35.1000 79.9000 ;
	    RECT 34.2000 75.9000 35.1000 76.3000 ;
	    RECT 35.8000 76.2000 36.2000 79.9000 ;
	    RECT 36.6000 76.2000 37.0000 76.3000 ;
	    RECT 35.8000 75.9000 37.0000 76.2000 ;
	    RECT 38.0000 75.9000 38.8000 79.9000 ;
	    RECT 39.7000 76.2000 40.1000 76.3000 ;
	    RECT 40.6000 76.2000 41.0000 79.9000 ;
	    RECT 39.7000 75.9000 41.0000 76.2000 ;
	    RECT 34.3000 74.2000 34.6000 75.9000 ;
	    RECT 35.0000 74.8000 35.4000 75.6000 ;
	    RECT 38.2000 75.2000 38.5000 75.9000 ;
	    RECT 39.1000 75.2000 39.5000 75.3000 ;
	    RECT 38.2000 74.8000 38.6000 75.2000 ;
	    RECT 39.1000 74.9000 39.9000 75.2000 ;
	    RECT 39.5000 74.8000 39.9000 74.9000 ;
	    RECT 38.2000 74.2000 38.5000 74.8000 ;
	    RECT 32.6000 74.1000 33.0000 74.2000 ;
	    RECT 34.2000 74.1000 34.6000 74.2000 ;
	    RECT 32.6000 73.8000 34.6000 74.1000 ;
	    RECT 37.2000 73.8000 37.6000 74.2000 ;
	    RECT 32.6000 73.4000 33.0000 73.8000 ;
	    RECT 23.0000 72.8000 23.9000 73.1000 ;
	    RECT 23.5000 72.2000 23.9000 72.8000 ;
	    RECT 23.0000 71.8000 23.9000 72.2000 ;
	    RECT 23.5000 71.1000 23.9000 71.8000 ;
	    RECT 24.6000 71.1000 25.0000 73.1000 ;
	    RECT 26.7000 72.6000 27.4000 73.1000 ;
	    RECT 27.8000 73.0000 29.8000 73.1000 ;
	    RECT 26.7000 71.1000 27.1000 72.6000 ;
	    RECT 27.8000 71.1000 28.2000 73.0000 ;
	    RECT 29.4000 71.1000 29.8000 73.0000 ;
	    RECT 30.2000 71.1000 30.6000 73.1000 ;
	    RECT 31.3000 72.8000 32.2000 73.1000 ;
	    RECT 31.3000 72.2000 31.7000 72.8000 ;
	    RECT 33.4000 72.4000 33.8000 73.2000 ;
	    RECT 31.0000 71.8000 31.7000 72.2000 ;
	    RECT 34.3000 72.1000 34.6000 73.8000 ;
	    RECT 37.3000 73.6000 37.6000 73.8000 ;
	    RECT 38.0000 73.9000 38.5000 74.2000 ;
	    RECT 41.4000 74.1000 41.8000 74.2000 ;
	    RECT 42.2000 74.1000 42.6000 79.9000 ;
	    RECT 43.4000 76.8000 43.8000 77.2000 ;
	    RECT 43.4000 76.2000 43.7000 76.8000 ;
	    RECT 44.1000 76.2000 44.5000 79.9000 ;
	    RECT 46.2000 76.2000 46.6000 79.9000 ;
	    RECT 47.8000 79.6000 49.8000 79.9000 ;
	    RECT 47.8000 76.2000 48.2000 79.6000 ;
	    RECT 43.0000 75.9000 43.7000 76.2000 ;
	    RECT 43.0000 75.8000 43.4000 75.9000 ;
	    RECT 44.0000 75.8000 45.0000 76.2000 ;
	    RECT 46.2000 75.9000 48.2000 76.2000 ;
	    RECT 48.6000 75.9000 49.0000 79.3000 ;
	    RECT 49.4000 75.9000 49.8000 79.6000 ;
	    RECT 44.0000 74.2000 44.3000 75.8000 ;
	    RECT 48.6000 75.6000 48.9000 75.9000 ;
	    RECT 46.6000 75.2000 47.0000 75.4000 ;
	    RECT 47.9000 75.3000 48.9000 75.6000 ;
	    RECT 47.9000 75.2000 48.2000 75.3000 ;
	    RECT 44.6000 74.4000 45.0000 75.2000 ;
	    RECT 46.2000 74.9000 47.0000 75.2000 ;
	    RECT 46.2000 74.8000 46.6000 74.9000 ;
	    RECT 47.8000 74.8000 48.2000 75.2000 ;
	    RECT 49.4000 74.8000 49.8000 75.6000 ;
	    RECT 36.6000 73.4000 37.0000 73.5000 ;
	    RECT 31.3000 71.1000 31.7000 71.8000 ;
	    RECT 34.2000 71.1000 34.6000 72.1000 ;
	    RECT 35.8000 73.1000 37.0000 73.4000 ;
	    RECT 37.3000 73.2000 37.7000 73.6000 ;
	    RECT 35.8000 71.1000 36.2000 73.1000 ;
	    RECT 38.0000 72.9000 38.3000 73.9000 ;
	    RECT 41.4000 73.8000 42.6000 74.1000 ;
	    RECT 43.0000 73.8000 44.3000 74.2000 ;
	    RECT 45.4000 74.1000 45.8000 74.2000 ;
	    RECT 46.2000 74.1000 46.5000 74.8000 ;
	    RECT 45.0000 73.8000 46.5000 74.1000 ;
	    RECT 47.0000 73.8000 47.4000 74.6000 ;
	    RECT 38.6000 73.2000 39.4000 73.6000 ;
	    RECT 39.7000 73.4000 40.1000 73.5000 ;
	    RECT 39.7000 73.1000 41.0000 73.4000 ;
	    RECT 38.0000 72.2000 38.8000 72.9000 ;
	    RECT 37.4000 71.8000 38.8000 72.2000 ;
	    RECT 38.0000 71.1000 38.8000 71.8000 ;
	    RECT 40.6000 71.1000 41.0000 73.1000 ;
	    RECT 41.4000 72.4000 41.8000 73.2000 ;
	    RECT 42.2000 71.1000 42.6000 73.8000 ;
	    RECT 43.1000 73.1000 43.4000 73.8000 ;
	    RECT 45.0000 73.6000 45.4000 73.8000 ;
	    RECT 43.9000 73.1000 45.7000 73.3000 ;
	    RECT 47.9000 73.1000 48.2000 74.8000 ;
	    RECT 48.5000 74.4000 48.9000 74.8000 ;
	    RECT 48.6000 74.2000 48.9000 74.4000 ;
	    RECT 48.6000 74.1000 49.0000 74.2000 ;
	    RECT 50.2000 74.1000 50.6000 79.9000 ;
	    RECT 53.1000 76.2000 53.5000 79.9000 ;
	    RECT 55.8000 77.9000 56.2000 79.9000 ;
	    RECT 55.9000 77.8000 56.2000 77.9000 ;
	    RECT 57.4000 79.1000 57.8000 79.9000 ;
	    RECT 58.2000 79.1000 58.6000 79.2000 ;
	    RECT 57.4000 78.8000 58.6000 79.1000 ;
	    RECT 57.4000 77.9000 57.8000 78.8000 ;
	    RECT 57.4000 77.8000 57.7000 77.9000 ;
	    RECT 55.9000 77.5000 57.7000 77.8000 ;
	    RECT 53.8000 76.8000 54.2000 77.2000 ;
	    RECT 53.9000 76.2000 54.2000 76.8000 ;
	    RECT 56.6000 76.4000 57.0000 77.2000 ;
	    RECT 57.4000 76.2000 57.7000 77.5000 ;
	    RECT 53.1000 75.9000 53.6000 76.2000 ;
	    RECT 53.9000 75.9000 54.6000 76.2000 ;
	    RECT 51.0000 75.1000 51.4000 75.2000 ;
	    RECT 52.6000 75.1000 53.0000 75.2000 ;
	    RECT 51.0000 74.8000 53.0000 75.1000 ;
	    RECT 52.6000 74.4000 53.0000 74.8000 ;
	    RECT 53.3000 74.2000 53.6000 75.9000 ;
	    RECT 54.2000 75.8000 54.6000 75.9000 ;
	    RECT 55.0000 75.4000 55.4000 76.2000 ;
	    RECT 57.4000 75.8000 57.8000 76.2000 ;
	    RECT 54.2000 74.8000 54.6000 75.2000 ;
	    RECT 55.8000 74.8000 56.6000 75.2000 ;
	    RECT 54.2000 74.2000 54.5000 74.8000 ;
	    RECT 57.4000 74.2000 57.7000 75.8000 ;
	    RECT 48.6000 73.8000 50.6000 74.1000 ;
	    RECT 51.8000 74.1000 52.2000 74.2000 ;
	    RECT 51.8000 73.8000 52.6000 74.1000 ;
	    RECT 53.3000 73.8000 54.6000 74.2000 ;
	    RECT 56.9000 74.1000 57.7000 74.2000 ;
	    RECT 56.8000 73.9000 57.7000 74.1000 ;
	    RECT 59.8000 75.6000 60.2000 79.9000 ;
	    RECT 61.9000 77.9000 62.5000 79.9000 ;
	    RECT 64.2000 77.9000 64.6000 79.9000 ;
	    RECT 66.4000 78.2000 66.8000 79.9000 ;
	    RECT 66.4000 77.9000 67.4000 78.2000 ;
	    RECT 62.2000 77.5000 62.6000 77.9000 ;
	    RECT 64.3000 77.6000 64.6000 77.9000 ;
	    RECT 63.9000 77.3000 65.7000 77.6000 ;
	    RECT 67.0000 77.5000 67.4000 77.9000 ;
	    RECT 63.9000 77.2000 64.3000 77.3000 ;
	    RECT 65.3000 77.2000 65.7000 77.3000 ;
	    RECT 61.8000 76.6000 62.5000 77.0000 ;
	    RECT 62.2000 76.1000 62.5000 76.6000 ;
	    RECT 63.3000 76.5000 64.4000 76.8000 ;
	    RECT 63.3000 76.4000 63.7000 76.5000 ;
	    RECT 62.2000 75.8000 63.4000 76.1000 ;
	    RECT 59.8000 75.3000 61.9000 75.6000 ;
	    RECT 43.0000 71.1000 43.4000 73.1000 ;
	    RECT 43.8000 73.0000 45.8000 73.1000 ;
	    RECT 43.8000 71.1000 44.2000 73.0000 ;
	    RECT 45.4000 71.1000 45.8000 73.0000 ;
	    RECT 47.7000 71.1000 48.5000 73.1000 ;
	    RECT 50.2000 71.1000 50.6000 73.8000 ;
	    RECT 52.2000 73.6000 52.6000 73.8000 ;
	    RECT 51.0000 72.4000 51.4000 73.2000 ;
	    RECT 51.9000 73.1000 53.7000 73.3000 ;
	    RECT 54.2000 73.1000 54.5000 73.8000 ;
	    RECT 51.8000 73.0000 53.8000 73.1000 ;
	    RECT 51.8000 71.1000 52.2000 73.0000 ;
	    RECT 53.4000 71.1000 53.8000 73.0000 ;
	    RECT 54.2000 71.1000 54.6000 73.1000 ;
	    RECT 56.8000 71.1000 57.2000 73.9000 ;
	    RECT 59.8000 73.6000 60.2000 75.3000 ;
	    RECT 61.5000 75.2000 61.9000 75.3000 ;
	    RECT 60.7000 74.9000 61.1000 75.0000 ;
	    RECT 60.7000 74.6000 62.6000 74.9000 ;
	    RECT 62.2000 74.5000 62.6000 74.6000 ;
	    RECT 63.1000 74.2000 63.4000 75.8000 ;
	    RECT 64.1000 75.9000 64.4000 76.5000 ;
	    RECT 64.7000 76.5000 65.1000 76.6000 ;
	    RECT 67.0000 76.5000 67.4000 76.6000 ;
	    RECT 64.7000 76.2000 67.4000 76.5000 ;
	    RECT 64.1000 75.7000 66.5000 75.9000 ;
	    RECT 68.6000 75.7000 69.0000 79.9000 ;
	    RECT 69.4000 75.9000 69.8000 79.9000 ;
	    RECT 70.2000 76.2000 70.6000 79.9000 ;
	    RECT 71.8000 76.2000 72.2000 79.9000 ;
	    RECT 73.0000 76.8000 73.4000 77.2000 ;
	    RECT 73.0000 76.2000 73.3000 76.8000 ;
	    RECT 73.7000 76.2000 74.1000 79.9000 ;
	    RECT 76.9000 79.2000 77.3000 79.9000 ;
	    RECT 76.9000 78.8000 77.8000 79.2000 ;
	    RECT 76.2000 76.8000 76.6000 77.2000 ;
	    RECT 76.2000 76.2000 76.5000 76.8000 ;
	    RECT 76.9000 76.2000 77.3000 78.8000 ;
	    RECT 70.2000 75.9000 72.2000 76.2000 ;
	    RECT 72.6000 75.9000 73.3000 76.2000 ;
	    RECT 73.6000 75.9000 74.1000 76.2000 ;
	    RECT 75.8000 75.9000 76.5000 76.2000 ;
	    RECT 76.8000 75.9000 77.3000 76.2000 ;
	    RECT 64.1000 75.6000 69.0000 75.7000 ;
	    RECT 66.1000 75.5000 69.0000 75.6000 ;
	    RECT 66.2000 75.4000 69.0000 75.5000 ;
	    RECT 69.5000 75.2000 69.8000 75.9000 ;
	    RECT 72.6000 75.8000 73.0000 75.9000 ;
	    RECT 71.4000 75.2000 71.8000 75.4000 ;
	    RECT 65.4000 75.1000 65.8000 75.2000 ;
	    RECT 65.4000 74.8000 67.9000 75.1000 ;
	    RECT 66.2000 74.7000 66.6000 74.8000 ;
	    RECT 67.5000 74.7000 67.9000 74.8000 ;
	    RECT 69.4000 74.9000 70.6000 75.2000 ;
	    RECT 71.4000 74.9000 72.2000 75.2000 ;
	    RECT 69.4000 74.8000 69.8000 74.9000 ;
	    RECT 66.7000 74.2000 67.1000 74.3000 ;
	    RECT 69.4000 74.2000 69.7000 74.8000 ;
	    RECT 63.1000 73.9000 68.6000 74.2000 ;
	    RECT 63.3000 73.8000 63.7000 73.9000 ;
	    RECT 59.8000 73.3000 61.7000 73.6000 ;
	    RECT 59.8000 71.1000 60.2000 73.3000 ;
	    RECT 61.3000 73.2000 61.7000 73.3000 ;
	    RECT 66.2000 72.8000 66.5000 73.9000 ;
	    RECT 67.8000 73.8000 68.6000 73.9000 ;
	    RECT 69.4000 73.8000 69.8000 74.2000 ;
	    RECT 65.3000 72.7000 65.7000 72.8000 ;
	    RECT 62.2000 72.1000 62.6000 72.5000 ;
	    RECT 64.3000 72.4000 65.7000 72.7000 ;
	    RECT 66.2000 72.4000 66.6000 72.8000 ;
	    RECT 64.3000 72.1000 64.6000 72.4000 ;
	    RECT 67.0000 72.1000 67.4000 72.5000 ;
	    RECT 61.9000 71.8000 62.6000 72.1000 ;
	    RECT 61.9000 71.1000 62.5000 71.8000 ;
	    RECT 64.2000 71.1000 64.6000 72.1000 ;
	    RECT 66.4000 71.8000 67.4000 72.1000 ;
	    RECT 66.4000 71.1000 66.8000 71.8000 ;
	    RECT 68.6000 71.1000 69.0000 73.5000 ;
	    RECT 69.4000 72.8000 69.8000 73.2000 ;
	    RECT 70.3000 73.1000 70.6000 74.9000 ;
	    RECT 71.8000 74.8000 72.2000 74.9000 ;
	    RECT 71.0000 74.1000 71.4000 74.6000 ;
	    RECT 73.6000 74.2000 73.9000 75.9000 ;
	    RECT 75.8000 75.8000 76.2000 75.9000 ;
	    RECT 74.2000 74.4000 74.6000 75.2000 ;
	    RECT 76.8000 74.2000 77.1000 75.9000 ;
	    RECT 79.0000 75.6000 79.4000 79.9000 ;
	    RECT 81.1000 77.9000 81.7000 79.9000 ;
	    RECT 83.4000 77.9000 83.8000 79.9000 ;
	    RECT 85.6000 78.2000 86.0000 79.9000 ;
	    RECT 85.6000 77.9000 86.6000 78.2000 ;
	    RECT 81.4000 77.5000 81.8000 77.9000 ;
	    RECT 83.5000 77.6000 83.8000 77.9000 ;
	    RECT 83.1000 77.3000 84.9000 77.6000 ;
	    RECT 86.2000 77.5000 86.6000 77.9000 ;
	    RECT 83.1000 77.2000 83.5000 77.3000 ;
	    RECT 84.5000 77.2000 84.9000 77.3000 ;
	    RECT 81.0000 76.6000 81.7000 77.0000 ;
	    RECT 81.4000 76.1000 81.7000 76.6000 ;
	    RECT 82.5000 76.5000 83.6000 76.8000 ;
	    RECT 82.5000 76.4000 82.9000 76.5000 ;
	    RECT 81.4000 75.8000 82.6000 76.1000 ;
	    RECT 79.0000 75.3000 81.1000 75.6000 ;
	    RECT 77.4000 74.4000 77.8000 75.2000 ;
	    RECT 72.6000 74.1000 73.9000 74.2000 ;
	    RECT 75.0000 74.1000 75.4000 74.2000 ;
	    RECT 71.0000 73.8000 73.9000 74.1000 ;
	    RECT 74.6000 73.8000 75.4000 74.1000 ;
	    RECT 75.8000 73.8000 77.1000 74.2000 ;
	    RECT 78.2000 74.1000 78.6000 74.2000 ;
	    RECT 77.8000 73.8000 78.6000 74.1000 ;
	    RECT 72.7000 73.1000 73.0000 73.8000 ;
	    RECT 74.6000 73.6000 75.0000 73.8000 ;
	    RECT 73.5000 73.1000 75.3000 73.3000 ;
	    RECT 75.9000 73.1000 76.2000 73.8000 ;
	    RECT 77.8000 73.6000 78.2000 73.8000 ;
	    RECT 79.0000 73.6000 79.4000 75.3000 ;
	    RECT 80.7000 75.2000 81.1000 75.3000 ;
	    RECT 79.9000 74.9000 80.3000 75.0000 ;
	    RECT 79.9000 74.6000 81.8000 74.9000 ;
	    RECT 81.4000 74.5000 81.8000 74.6000 ;
	    RECT 82.3000 74.2000 82.6000 75.8000 ;
	    RECT 83.3000 75.9000 83.6000 76.5000 ;
	    RECT 83.9000 76.5000 84.3000 76.6000 ;
	    RECT 86.2000 76.5000 86.6000 76.6000 ;
	    RECT 83.9000 76.2000 86.6000 76.5000 ;
	    RECT 83.3000 75.7000 85.7000 75.9000 ;
	    RECT 87.8000 75.7000 88.2000 79.9000 ;
	    RECT 83.3000 75.6000 88.2000 75.7000 ;
	    RECT 85.3000 75.5000 88.2000 75.6000 ;
	    RECT 85.4000 75.4000 88.2000 75.5000 ;
	    RECT 84.6000 75.1000 85.0000 75.2000 ;
	    RECT 88.6000 75.1000 89.0000 79.9000 ;
	    RECT 89.4000 75.8000 89.8000 76.2000 ;
	    RECT 90.2000 75.8000 90.6000 76.6000 ;
	    RECT 89.4000 75.1000 89.7000 75.8000 ;
	    RECT 84.6000 74.8000 87.1000 75.1000 ;
	    RECT 85.4000 74.7000 85.8000 74.8000 ;
	    RECT 86.7000 74.7000 87.1000 74.8000 ;
	    RECT 88.6000 74.8000 89.7000 75.1000 ;
	    RECT 85.9000 74.2000 86.3000 74.3000 ;
	    RECT 82.3000 73.9000 87.8000 74.2000 ;
	    RECT 82.5000 73.8000 82.9000 73.9000 ;
	    RECT 84.6000 73.8000 85.0000 73.9000 ;
	    RECT 79.0000 73.3000 80.9000 73.6000 ;
	    RECT 76.7000 73.1000 78.5000 73.3000 ;
	    RECT 69.5000 72.4000 69.9000 72.8000 ;
	    RECT 70.2000 71.1000 70.6000 73.1000 ;
	    RECT 72.6000 71.1000 73.0000 73.1000 ;
	    RECT 73.4000 73.0000 75.4000 73.1000 ;
	    RECT 73.4000 71.1000 73.8000 73.0000 ;
	    RECT 75.0000 71.1000 75.4000 73.0000 ;
	    RECT 75.8000 71.1000 76.2000 73.1000 ;
	    RECT 76.6000 73.0000 78.6000 73.1000 ;
	    RECT 76.6000 71.1000 77.0000 73.0000 ;
	    RECT 78.2000 71.1000 78.6000 73.0000 ;
	    RECT 79.0000 71.1000 79.4000 73.3000 ;
	    RECT 80.5000 73.2000 80.9000 73.3000 ;
	    RECT 85.4000 72.8000 85.7000 73.9000 ;
	    RECT 87.0000 73.8000 87.8000 73.9000 ;
	    RECT 84.5000 72.7000 84.9000 72.8000 ;
	    RECT 81.4000 72.1000 81.8000 72.5000 ;
	    RECT 83.5000 72.4000 84.9000 72.7000 ;
	    RECT 85.4000 72.4000 85.8000 72.8000 ;
	    RECT 83.5000 72.1000 83.8000 72.4000 ;
	    RECT 86.2000 72.1000 86.6000 72.5000 ;
	    RECT 81.1000 71.8000 81.8000 72.1000 ;
	    RECT 81.1000 71.1000 81.7000 71.8000 ;
	    RECT 83.4000 71.1000 83.8000 72.1000 ;
	    RECT 85.6000 71.8000 86.6000 72.1000 ;
	    RECT 85.6000 71.1000 86.0000 71.8000 ;
	    RECT 87.8000 71.1000 88.2000 73.5000 ;
	    RECT 88.6000 71.1000 89.0000 74.8000 ;
	    RECT 89.4000 73.1000 89.8000 73.2000 ;
	    RECT 91.0000 73.1000 91.4000 79.9000 ;
	    RECT 93.9000 76.2000 94.3000 79.9000 ;
	    RECT 94.6000 76.8000 95.0000 77.2000 ;
	    RECT 94.7000 76.2000 95.0000 76.8000 ;
	    RECT 96.1000 76.3000 96.5000 79.9000 ;
	    RECT 99.0000 76.4000 99.4000 79.9000 ;
	    RECT 93.9000 75.9000 94.4000 76.2000 ;
	    RECT 94.7000 75.9000 95.4000 76.2000 ;
	    RECT 96.1000 75.9000 97.0000 76.3000 ;
	    RECT 98.9000 75.9000 99.4000 76.4000 ;
	    RECT 100.6000 76.2000 101.0000 79.9000 ;
	    RECT 99.7000 75.9000 101.0000 76.2000 ;
	    RECT 101.4000 76.2000 101.8000 79.9000 ;
	    RECT 103.0000 76.2000 103.4000 79.9000 ;
	    RECT 101.4000 75.9000 103.4000 76.2000 ;
	    RECT 103.8000 75.9000 104.2000 79.9000 ;
	    RECT 93.4000 75.1000 93.8000 75.2000 ;
	    RECT 91.8000 74.8000 93.8000 75.1000 ;
	    RECT 91.8000 74.2000 92.1000 74.8000 ;
	    RECT 93.4000 74.4000 93.8000 74.8000 ;
	    RECT 94.1000 74.2000 94.4000 75.9000 ;
	    RECT 95.0000 75.8000 95.4000 75.9000 ;
	    RECT 95.8000 74.8000 96.2000 75.6000 ;
	    RECT 96.6000 75.1000 96.9000 75.9000 ;
	    RECT 96.6000 74.8000 97.7000 75.1000 ;
	    RECT 96.6000 74.2000 96.9000 74.8000 ;
	    RECT 97.4000 74.2000 97.7000 74.8000 ;
	    RECT 98.9000 74.2000 99.2000 75.9000 ;
	    RECT 99.7000 74.9000 100.0000 75.9000 ;
	    RECT 101.8000 75.2000 102.2000 75.4000 ;
	    RECT 103.8000 75.2000 104.1000 75.9000 ;
	    RECT 106.2000 75.7000 106.6000 79.9000 ;
	    RECT 108.4000 78.2000 108.8000 79.9000 ;
	    RECT 107.8000 77.9000 108.8000 78.2000 ;
	    RECT 110.6000 77.9000 111.0000 79.9000 ;
	    RECT 112.7000 77.9000 113.3000 79.9000 ;
	    RECT 107.8000 77.5000 108.2000 77.9000 ;
	    RECT 110.6000 77.6000 110.9000 77.9000 ;
	    RECT 109.5000 77.3000 111.3000 77.6000 ;
	    RECT 112.6000 77.5000 113.0000 77.9000 ;
	    RECT 109.5000 77.2000 109.9000 77.3000 ;
	    RECT 110.9000 77.2000 111.3000 77.3000 ;
	    RECT 107.8000 76.5000 108.2000 76.6000 ;
	    RECT 110.1000 76.5000 110.5000 76.6000 ;
	    RECT 107.8000 76.2000 110.5000 76.5000 ;
	    RECT 110.8000 76.5000 111.9000 76.8000 ;
	    RECT 110.8000 75.9000 111.1000 76.5000 ;
	    RECT 111.5000 76.4000 111.9000 76.5000 ;
	    RECT 112.7000 76.6000 113.4000 77.0000 ;
	    RECT 112.7000 76.1000 113.0000 76.6000 ;
	    RECT 108.7000 75.7000 111.1000 75.9000 ;
	    RECT 106.2000 75.6000 111.1000 75.7000 ;
	    RECT 111.8000 75.8000 113.0000 76.1000 ;
	    RECT 106.2000 75.5000 109.1000 75.6000 ;
	    RECT 106.2000 75.4000 109.0000 75.5000 ;
	    RECT 111.8000 75.2000 112.1000 75.8000 ;
	    RECT 115.0000 75.6000 115.4000 79.9000 ;
	    RECT 115.8000 76.2000 116.2000 79.9000 ;
	    RECT 117.4000 76.4000 117.8000 79.9000 ;
	    RECT 115.8000 75.9000 117.1000 76.2000 ;
	    RECT 117.4000 75.9000 117.9000 76.4000 ;
	    RECT 113.3000 75.3000 115.4000 75.6000 ;
	    RECT 113.3000 75.2000 113.7000 75.3000 ;
	    RECT 99.5000 74.5000 100.0000 74.9000 ;
	    RECT 91.8000 73.4000 92.2000 74.2000 ;
	    RECT 92.6000 74.1000 93.0000 74.2000 ;
	    RECT 92.6000 73.8000 93.4000 74.1000 ;
	    RECT 94.1000 73.8000 95.4000 74.2000 ;
	    RECT 95.8000 73.8000 96.2000 74.2000 ;
	    RECT 96.6000 73.8000 97.0000 74.2000 ;
	    RECT 97.4000 73.8000 97.8000 74.2000 ;
	    RECT 98.9000 73.8000 99.4000 74.2000 ;
	    RECT 93.0000 73.6000 93.4000 73.8000 ;
	    RECT 92.7000 73.1000 94.5000 73.3000 ;
	    RECT 95.0000 73.1000 95.3000 73.8000 ;
	    RECT 95.8000 73.1000 96.1000 73.8000 ;
	    RECT 89.4000 72.8000 91.4000 73.1000 ;
	    RECT 92.6000 73.0000 94.6000 73.1000 ;
	    RECT 89.4000 72.4000 89.8000 72.8000 ;
	    RECT 90.5000 71.1000 90.9000 72.8000 ;
	    RECT 92.6000 71.1000 93.0000 73.0000 ;
	    RECT 94.2000 71.1000 94.6000 73.0000 ;
	    RECT 95.0000 72.8000 96.1000 73.1000 ;
	    RECT 95.0000 71.1000 95.4000 72.8000 ;
	    RECT 96.6000 72.1000 96.9000 73.8000 ;
	    RECT 97.4000 72.4000 97.8000 73.2000 ;
	    RECT 98.9000 73.1000 99.2000 73.8000 ;
	    RECT 99.7000 73.7000 100.0000 74.5000 ;
	    RECT 100.5000 74.8000 101.0000 75.2000 ;
	    RECT 101.4000 74.9000 102.2000 75.2000 ;
	    RECT 103.0000 74.9000 104.2000 75.2000 ;
	    RECT 109.4000 75.1000 109.8000 75.2000 ;
	    RECT 101.4000 74.8000 101.8000 74.9000 ;
	    RECT 100.5000 74.4000 100.9000 74.8000 ;
	    RECT 102.2000 73.8000 102.6000 74.6000 ;
	    RECT 99.7000 73.4000 101.0000 73.7000 ;
	    RECT 98.9000 72.8000 99.4000 73.1000 ;
	    RECT 96.6000 71.1000 97.0000 72.1000 ;
	    RECT 99.0000 71.1000 99.4000 72.8000 ;
	    RECT 100.6000 71.1000 101.0000 73.4000 ;
	    RECT 103.0000 73.1000 103.3000 74.9000 ;
	    RECT 103.8000 74.8000 104.2000 74.9000 ;
	    RECT 107.3000 74.8000 109.8000 75.1000 ;
	    RECT 111.8000 74.8000 112.2000 75.2000 ;
	    RECT 114.1000 74.9000 114.5000 75.0000 ;
	    RECT 107.3000 74.7000 107.7000 74.8000 ;
	    RECT 108.6000 74.7000 109.0000 74.8000 ;
	    RECT 108.1000 74.2000 108.5000 74.3000 ;
	    RECT 111.8000 74.2000 112.1000 74.8000 ;
	    RECT 112.6000 74.6000 114.5000 74.9000 ;
	    RECT 112.6000 74.5000 113.0000 74.6000 ;
	    RECT 106.6000 73.9000 112.1000 74.2000 ;
	    RECT 106.6000 73.8000 107.4000 73.9000 ;
	    RECT 103.0000 71.1000 103.4000 73.1000 ;
	    RECT 103.8000 72.8000 104.2000 73.2000 ;
	    RECT 103.7000 72.4000 104.1000 72.8000 ;
	    RECT 106.2000 71.1000 106.6000 73.5000 ;
	    RECT 108.7000 72.8000 109.0000 73.9000 ;
	    RECT 111.5000 73.8000 111.9000 73.9000 ;
	    RECT 115.0000 73.6000 115.4000 75.3000 ;
	    RECT 115.8000 74.8000 116.3000 75.2000 ;
	    RECT 115.9000 74.4000 116.3000 74.8000 ;
	    RECT 116.8000 74.9000 117.1000 75.9000 ;
	    RECT 116.8000 74.5000 117.3000 74.9000 ;
	    RECT 116.8000 73.7000 117.1000 74.5000 ;
	    RECT 117.6000 74.2000 117.9000 75.9000 ;
	    RECT 119.0000 75.7000 119.4000 79.9000 ;
	    RECT 121.2000 78.2000 121.6000 79.9000 ;
	    RECT 120.6000 77.9000 121.6000 78.2000 ;
	    RECT 123.4000 77.9000 123.8000 79.9000 ;
	    RECT 125.5000 77.9000 126.1000 79.9000 ;
	    RECT 120.6000 77.5000 121.0000 77.9000 ;
	    RECT 123.4000 77.6000 123.7000 77.9000 ;
	    RECT 122.3000 77.3000 124.1000 77.6000 ;
	    RECT 125.4000 77.5000 125.8000 77.9000 ;
	    RECT 122.3000 77.2000 122.7000 77.3000 ;
	    RECT 123.7000 77.2000 124.1000 77.3000 ;
	    RECT 120.6000 76.5000 121.0000 76.6000 ;
	    RECT 122.9000 76.5000 123.3000 76.6000 ;
	    RECT 120.6000 76.2000 123.3000 76.5000 ;
	    RECT 123.6000 76.5000 124.7000 76.8000 ;
	    RECT 123.6000 75.9000 123.9000 76.5000 ;
	    RECT 124.3000 76.4000 124.7000 76.5000 ;
	    RECT 125.5000 76.6000 126.2000 77.0000 ;
	    RECT 125.5000 76.1000 125.8000 76.6000 ;
	    RECT 121.5000 75.7000 123.9000 75.9000 ;
	    RECT 119.0000 75.6000 123.9000 75.7000 ;
	    RECT 124.6000 75.8000 125.8000 76.1000 ;
	    RECT 119.0000 75.5000 121.9000 75.6000 ;
	    RECT 119.0000 75.4000 121.8000 75.5000 ;
	    RECT 124.6000 75.2000 124.9000 75.8000 ;
	    RECT 127.8000 75.6000 128.2000 79.9000 ;
	    RECT 126.1000 75.3000 128.2000 75.6000 ;
	    RECT 126.1000 75.2000 126.5000 75.3000 ;
	    RECT 122.2000 75.1000 122.6000 75.2000 ;
	    RECT 120.1000 74.8000 122.6000 75.1000 ;
	    RECT 124.6000 74.8000 125.0000 75.2000 ;
	    RECT 126.9000 74.9000 127.3000 75.0000 ;
	    RECT 120.1000 74.7000 120.5000 74.8000 ;
	    RECT 121.4000 74.7000 121.8000 74.8000 ;
	    RECT 120.9000 74.2000 121.3000 74.3000 ;
	    RECT 124.6000 74.2000 124.9000 74.8000 ;
	    RECT 125.4000 74.6000 127.3000 74.9000 ;
	    RECT 125.4000 74.5000 125.8000 74.6000 ;
	    RECT 117.4000 73.8000 117.9000 74.2000 ;
	    RECT 118.2000 74.1000 118.6000 74.2000 ;
	    RECT 119.4000 74.1000 124.9000 74.2000 ;
	    RECT 118.2000 73.9000 124.9000 74.1000 ;
	    RECT 118.2000 73.8000 120.2000 73.9000 ;
	    RECT 113.5000 73.3000 115.4000 73.6000 ;
	    RECT 113.5000 73.2000 113.9000 73.3000 ;
	    RECT 107.8000 72.1000 108.2000 72.5000 ;
	    RECT 108.6000 72.4000 109.0000 72.8000 ;
	    RECT 109.5000 72.7000 109.9000 72.8000 ;
	    RECT 109.5000 72.4000 110.9000 72.7000 ;
	    RECT 110.6000 72.1000 110.9000 72.4000 ;
	    RECT 112.6000 72.1000 113.0000 72.5000 ;
	    RECT 107.8000 71.8000 108.8000 72.1000 ;
	    RECT 108.4000 71.1000 108.8000 71.8000 ;
	    RECT 110.6000 71.1000 111.0000 72.1000 ;
	    RECT 112.6000 71.8000 113.3000 72.1000 ;
	    RECT 112.7000 71.1000 113.3000 71.8000 ;
	    RECT 115.0000 71.1000 115.4000 73.3000 ;
	    RECT 115.8000 73.4000 117.1000 73.7000 ;
	    RECT 115.8000 71.1000 116.2000 73.4000 ;
	    RECT 117.6000 73.1000 117.9000 73.8000 ;
	    RECT 117.4000 72.8000 117.9000 73.1000 ;
	    RECT 117.4000 71.1000 117.8000 72.8000 ;
	    RECT 119.0000 71.1000 119.4000 73.5000 ;
	    RECT 121.5000 72.8000 121.8000 73.9000 ;
	    RECT 124.3000 73.8000 124.7000 73.9000 ;
	    RECT 127.8000 73.6000 128.2000 75.3000 ;
	    RECT 126.3000 73.3000 128.2000 73.6000 ;
	    RECT 126.3000 73.2000 126.7000 73.3000 ;
	    RECT 120.6000 72.1000 121.0000 72.5000 ;
	    RECT 121.4000 72.4000 121.8000 72.8000 ;
	    RECT 122.3000 72.7000 122.7000 72.8000 ;
	    RECT 122.3000 72.4000 123.7000 72.7000 ;
	    RECT 123.4000 72.1000 123.7000 72.4000 ;
	    RECT 125.4000 72.1000 125.8000 72.5000 ;
	    RECT 120.6000 71.8000 121.6000 72.1000 ;
	    RECT 121.2000 71.1000 121.6000 71.8000 ;
	    RECT 123.4000 71.1000 123.8000 72.1000 ;
	    RECT 125.4000 71.8000 126.1000 72.1000 ;
	    RECT 125.5000 71.1000 126.1000 71.8000 ;
	    RECT 127.8000 71.1000 128.2000 73.3000 ;
	    RECT 128.6000 75.6000 129.0000 79.9000 ;
	    RECT 130.7000 77.9000 131.3000 79.9000 ;
	    RECT 133.0000 77.9000 133.4000 79.9000 ;
	    RECT 135.2000 78.2000 135.6000 79.9000 ;
	    RECT 135.2000 77.9000 136.2000 78.2000 ;
	    RECT 131.0000 77.5000 131.4000 77.9000 ;
	    RECT 133.1000 77.6000 133.4000 77.9000 ;
	    RECT 132.7000 77.3000 134.5000 77.6000 ;
	    RECT 135.8000 77.5000 136.2000 77.9000 ;
	    RECT 132.7000 77.2000 133.1000 77.3000 ;
	    RECT 134.1000 77.2000 134.5000 77.3000 ;
	    RECT 130.6000 76.6000 131.3000 77.0000 ;
	    RECT 131.0000 76.1000 131.3000 76.6000 ;
	    RECT 132.1000 76.5000 133.2000 76.8000 ;
	    RECT 132.1000 76.4000 132.5000 76.5000 ;
	    RECT 131.0000 75.8000 132.2000 76.1000 ;
	    RECT 128.6000 75.3000 130.7000 75.6000 ;
	    RECT 128.6000 73.6000 129.0000 75.3000 ;
	    RECT 130.3000 75.2000 130.7000 75.3000 ;
	    RECT 129.5000 74.9000 129.9000 75.0000 ;
	    RECT 129.5000 74.6000 131.4000 74.9000 ;
	    RECT 131.0000 74.5000 131.4000 74.6000 ;
	    RECT 131.9000 74.2000 132.2000 75.8000 ;
	    RECT 132.9000 75.9000 133.2000 76.5000 ;
	    RECT 133.5000 76.5000 133.9000 76.6000 ;
	    RECT 135.8000 76.5000 136.2000 76.6000 ;
	    RECT 133.5000 76.2000 136.2000 76.5000 ;
	    RECT 132.9000 75.7000 135.3000 75.9000 ;
	    RECT 137.4000 75.7000 137.8000 79.9000 ;
	    RECT 138.2000 76.2000 138.6000 79.9000 ;
	    RECT 139.8000 76.4000 140.2000 79.9000 ;
	    RECT 142.7000 79.2000 143.1000 79.9000 ;
	    RECT 142.2000 78.8000 143.1000 79.2000 ;
	    RECT 138.2000 75.9000 139.5000 76.2000 ;
	    RECT 139.8000 75.9000 140.3000 76.4000 ;
	    RECT 142.7000 76.2000 143.1000 78.8000 ;
	    RECT 143.4000 76.8000 143.8000 77.2000 ;
	    RECT 143.5000 76.2000 143.8000 76.8000 ;
	    RECT 142.7000 75.9000 143.2000 76.2000 ;
	    RECT 143.5000 75.9000 144.2000 76.2000 ;
	    RECT 132.9000 75.6000 137.8000 75.7000 ;
	    RECT 134.9000 75.5000 137.8000 75.6000 ;
	    RECT 135.0000 75.4000 137.8000 75.5000 ;
	    RECT 134.2000 75.1000 134.6000 75.2000 ;
	    RECT 134.2000 74.8000 136.7000 75.1000 ;
	    RECT 138.2000 74.8000 138.7000 75.2000 ;
	    RECT 135.0000 74.7000 135.4000 74.8000 ;
	    RECT 136.3000 74.7000 136.7000 74.8000 ;
	    RECT 138.3000 74.4000 138.7000 74.8000 ;
	    RECT 139.2000 74.9000 139.5000 75.9000 ;
	    RECT 139.2000 74.5000 139.7000 74.9000 ;
	    RECT 135.5000 74.2000 135.9000 74.3000 ;
	    RECT 131.9000 73.9000 137.4000 74.2000 ;
	    RECT 132.1000 73.8000 132.5000 73.9000 ;
	    RECT 128.6000 73.3000 130.5000 73.6000 ;
	    RECT 128.6000 71.1000 129.0000 73.3000 ;
	    RECT 130.1000 73.2000 130.5000 73.3000 ;
	    RECT 135.0000 72.8000 135.3000 73.9000 ;
	    RECT 136.6000 73.8000 137.4000 73.9000 ;
	    RECT 139.2000 73.7000 139.5000 74.5000 ;
	    RECT 140.0000 74.2000 140.3000 75.9000 ;
	    RECT 142.9000 74.2000 143.2000 75.9000 ;
	    RECT 143.8000 75.8000 144.2000 75.9000 ;
	    RECT 145.4000 75.6000 145.8000 79.9000 ;
	    RECT 147.0000 75.6000 147.4000 79.9000 ;
	    RECT 148.6000 75.6000 149.0000 79.9000 ;
	    RECT 150.2000 75.6000 150.6000 79.9000 ;
	    RECT 152.6000 75.6000 153.0000 79.9000 ;
	    RECT 154.2000 75.6000 154.6000 79.9000 ;
	    RECT 155.8000 75.6000 156.2000 79.9000 ;
	    RECT 157.4000 75.6000 157.8000 79.9000 ;
	    RECT 161.4000 77.9000 161.8000 79.9000 ;
	    RECT 144.6000 75.2000 145.8000 75.6000 ;
	    RECT 146.3000 75.2000 147.4000 75.6000 ;
	    RECT 147.9000 75.2000 149.0000 75.6000 ;
	    RECT 149.7000 75.2000 150.6000 75.6000 ;
	    RECT 151.8000 75.2000 153.0000 75.6000 ;
	    RECT 153.5000 75.2000 154.6000 75.6000 ;
	    RECT 155.1000 75.2000 156.2000 75.6000 ;
	    RECT 156.9000 75.2000 157.8000 75.6000 ;
	    RECT 161.5000 75.8000 161.8000 77.9000 ;
	    RECT 163.0000 75.9000 163.4000 79.9000 ;
	    RECT 161.5000 75.5000 162.7000 75.8000 ;
	    RECT 139.8000 74.1000 140.3000 74.2000 ;
	    RECT 141.4000 74.1000 141.8000 74.2000 ;
	    RECT 139.8000 73.8000 142.2000 74.1000 ;
	    RECT 142.9000 73.8000 144.2000 74.2000 ;
	    RECT 144.6000 73.8000 145.0000 75.2000 ;
	    RECT 146.3000 74.5000 146.7000 75.2000 ;
	    RECT 147.9000 74.5000 148.3000 75.2000 ;
	    RECT 149.7000 74.5000 150.1000 75.2000 ;
	    RECT 145.4000 74.1000 146.7000 74.5000 ;
	    RECT 147.1000 74.1000 148.3000 74.5000 ;
	    RECT 148.8000 74.1000 150.1000 74.5000 ;
	    RECT 146.3000 73.8000 146.7000 74.1000 ;
	    RECT 147.9000 73.8000 148.3000 74.1000 ;
	    RECT 149.7000 73.8000 150.1000 74.1000 ;
	    RECT 151.8000 73.8000 152.2000 75.2000 ;
	    RECT 153.5000 74.5000 153.9000 75.2000 ;
	    RECT 155.1000 74.5000 155.5000 75.2000 ;
	    RECT 156.9000 74.5000 157.3000 75.2000 ;
	    RECT 161.4000 74.8000 161.8000 75.2000 ;
	    RECT 152.6000 74.1000 153.9000 74.5000 ;
	    RECT 154.3000 74.1000 155.5000 74.5000 ;
	    RECT 156.0000 74.1000 157.3000 74.5000 ;
	    RECT 153.5000 73.8000 153.9000 74.1000 ;
	    RECT 155.1000 73.8000 155.5000 74.1000 ;
	    RECT 156.9000 73.8000 157.3000 74.1000 ;
	    RECT 160.6000 73.8000 161.0000 74.6000 ;
	    RECT 161.5000 74.4000 161.8000 74.8000 ;
	    RECT 161.5000 74.1000 162.0000 74.4000 ;
	    RECT 161.6000 74.0000 162.0000 74.1000 ;
	    RECT 162.4000 73.8000 162.7000 75.5000 ;
	    RECT 163.1000 75.2000 163.4000 75.9000 ;
	    RECT 163.0000 74.8000 163.4000 75.2000 ;
	    RECT 134.1000 72.7000 134.5000 72.8000 ;
	    RECT 131.0000 72.1000 131.4000 72.5000 ;
	    RECT 133.1000 72.4000 134.5000 72.7000 ;
	    RECT 135.0000 72.4000 135.4000 72.8000 ;
	    RECT 133.1000 72.1000 133.4000 72.4000 ;
	    RECT 135.8000 72.1000 136.2000 72.5000 ;
	    RECT 130.7000 71.8000 131.4000 72.1000 ;
	    RECT 130.7000 71.1000 131.3000 71.8000 ;
	    RECT 133.0000 71.1000 133.4000 72.1000 ;
	    RECT 135.2000 71.8000 136.2000 72.1000 ;
	    RECT 135.2000 71.1000 135.6000 71.8000 ;
	    RECT 137.4000 71.1000 137.8000 73.5000 ;
	    RECT 138.2000 73.4000 139.5000 73.7000 ;
	    RECT 138.2000 71.1000 138.6000 73.4000 ;
	    RECT 140.0000 73.1000 140.3000 73.8000 ;
	    RECT 141.8000 73.6000 142.2000 73.8000 ;
	    RECT 141.5000 73.1000 143.3000 73.3000 ;
	    RECT 143.8000 73.1000 144.1000 73.8000 ;
	    RECT 144.6000 73.4000 145.8000 73.8000 ;
	    RECT 146.3000 73.4000 147.4000 73.8000 ;
	    RECT 147.9000 73.4000 149.0000 73.8000 ;
	    RECT 149.7000 73.4000 150.6000 73.8000 ;
	    RECT 151.8000 73.4000 153.0000 73.8000 ;
	    RECT 153.5000 73.4000 154.6000 73.8000 ;
	    RECT 155.1000 73.4000 156.2000 73.8000 ;
	    RECT 156.9000 73.4000 157.8000 73.8000 ;
	    RECT 162.4000 73.7000 162.8000 73.8000 ;
	    RECT 161.3000 73.5000 162.8000 73.7000 ;
	    RECT 139.8000 72.8000 140.3000 73.1000 ;
	    RECT 141.4000 73.0000 143.4000 73.1000 ;
	    RECT 139.8000 71.1000 140.2000 72.8000 ;
	    RECT 141.4000 71.1000 141.8000 73.0000 ;
	    RECT 143.0000 71.1000 143.4000 73.0000 ;
	    RECT 143.8000 71.1000 144.2000 73.1000 ;
	    RECT 145.4000 71.1000 145.8000 73.4000 ;
	    RECT 147.0000 71.1000 147.4000 73.4000 ;
	    RECT 148.6000 71.1000 149.0000 73.4000 ;
	    RECT 150.2000 71.1000 150.6000 73.4000 ;
	    RECT 152.6000 71.1000 153.0000 73.4000 ;
	    RECT 154.2000 71.1000 154.6000 73.4000 ;
	    RECT 155.8000 71.1000 156.2000 73.4000 ;
	    RECT 157.4000 71.1000 157.8000 73.4000 ;
	    RECT 160.7000 73.4000 162.8000 73.5000 ;
	    RECT 160.7000 73.2000 161.6000 73.4000 ;
	    RECT 160.7000 73.1000 161.0000 73.2000 ;
	    RECT 163.1000 73.1000 163.4000 74.8000 ;
	    RECT 163.8000 73.4000 164.2000 74.2000 ;
	    RECT 160.6000 71.1000 161.0000 73.1000 ;
	    RECT 162.7000 72.6000 163.4000 73.1000 ;
	    RECT 164.6000 73.1000 165.0000 79.9000 ;
	    RECT 165.4000 76.1000 165.8000 76.6000 ;
	    RECT 166.2000 76.1000 166.6000 79.9000 ;
	    RECT 165.4000 75.8000 166.6000 76.1000 ;
	    RECT 164.6000 72.8000 165.5000 73.1000 ;
	    RECT 162.7000 72.2000 163.1000 72.6000 ;
	    RECT 165.1000 72.2000 165.5000 72.8000 ;
	    RECT 162.7000 71.8000 163.4000 72.2000 ;
	    RECT 164.6000 71.8000 165.5000 72.2000 ;
	    RECT 162.7000 71.1000 163.1000 71.8000 ;
	    RECT 165.1000 71.1000 165.5000 71.8000 ;
	    RECT 166.2000 71.1000 166.6000 75.8000 ;
	    RECT 167.8000 75.7000 168.2000 79.9000 ;
	    RECT 170.0000 78.2000 170.4000 79.9000 ;
	    RECT 169.4000 77.9000 170.4000 78.2000 ;
	    RECT 172.2000 77.9000 172.6000 79.9000 ;
	    RECT 174.3000 77.9000 174.9000 79.9000 ;
	    RECT 169.4000 77.5000 169.8000 77.9000 ;
	    RECT 172.2000 77.6000 172.5000 77.9000 ;
	    RECT 171.1000 77.3000 172.9000 77.6000 ;
	    RECT 174.2000 77.5000 174.6000 77.9000 ;
	    RECT 171.1000 77.2000 171.5000 77.3000 ;
	    RECT 172.5000 77.2000 172.9000 77.3000 ;
	    RECT 169.4000 76.5000 169.8000 76.6000 ;
	    RECT 171.7000 76.5000 172.1000 76.6000 ;
	    RECT 169.4000 76.2000 172.1000 76.5000 ;
	    RECT 172.4000 76.5000 173.5000 76.8000 ;
	    RECT 172.4000 75.9000 172.7000 76.5000 ;
	    RECT 173.1000 76.4000 173.5000 76.5000 ;
	    RECT 174.3000 76.6000 175.0000 77.0000 ;
	    RECT 174.3000 76.1000 174.6000 76.6000 ;
	    RECT 170.3000 75.7000 172.7000 75.9000 ;
	    RECT 167.8000 75.6000 172.7000 75.7000 ;
	    RECT 173.4000 75.8000 174.6000 76.1000 ;
	    RECT 167.8000 75.5000 170.7000 75.6000 ;
	    RECT 167.8000 75.4000 170.6000 75.5000 ;
	    RECT 173.4000 75.2000 173.7000 75.8000 ;
	    RECT 176.6000 75.6000 177.0000 79.9000 ;
	    RECT 177.4000 75.8000 177.8000 76.6000 ;
	    RECT 174.9000 75.3000 177.0000 75.6000 ;
	    RECT 174.9000 75.2000 175.3000 75.3000 ;
	    RECT 171.0000 75.1000 171.4000 75.2000 ;
	    RECT 168.9000 74.8000 171.4000 75.1000 ;
	    RECT 173.4000 74.8000 173.8000 75.2000 ;
	    RECT 175.7000 74.9000 176.1000 75.0000 ;
	    RECT 168.9000 74.7000 169.3000 74.8000 ;
	    RECT 169.7000 74.2000 170.1000 74.3000 ;
	    RECT 173.4000 74.2000 173.7000 74.8000 ;
	    RECT 174.2000 74.6000 176.1000 74.9000 ;
	    RECT 174.2000 74.5000 174.6000 74.6000 ;
	    RECT 168.2000 73.9000 173.7000 74.2000 ;
	    RECT 168.2000 73.8000 169.0000 73.9000 ;
	    RECT 167.0000 72.4000 167.4000 73.2000 ;
	    RECT 167.8000 71.1000 168.2000 73.5000 ;
	    RECT 170.3000 72.8000 170.6000 73.9000 ;
	    RECT 173.1000 73.8000 173.5000 73.9000 ;
	    RECT 176.6000 73.6000 177.0000 75.3000 ;
	    RECT 175.1000 73.3000 177.0000 73.6000 ;
	    RECT 175.1000 73.2000 175.5000 73.3000 ;
	    RECT 169.4000 72.1000 169.8000 72.5000 ;
	    RECT 170.2000 72.4000 170.6000 72.8000 ;
	    RECT 171.1000 72.7000 171.5000 72.8000 ;
	    RECT 171.1000 72.4000 172.5000 72.7000 ;
	    RECT 172.2000 72.1000 172.5000 72.4000 ;
	    RECT 174.2000 72.1000 174.6000 72.5000 ;
	    RECT 169.4000 71.8000 170.4000 72.1000 ;
	    RECT 170.0000 71.1000 170.4000 71.8000 ;
	    RECT 172.2000 71.1000 172.6000 72.1000 ;
	    RECT 174.2000 71.8000 174.9000 72.1000 ;
	    RECT 174.3000 71.1000 174.9000 71.8000 ;
	    RECT 176.6000 71.1000 177.0000 73.3000 ;
	    RECT 178.2000 73.1000 178.6000 79.9000 ;
	    RECT 179.8000 75.9000 180.2000 79.9000 ;
	    RECT 180.6000 76.2000 181.0000 79.9000 ;
	    RECT 182.2000 76.2000 182.6000 79.9000 ;
	    RECT 183.0000 77.9000 183.4000 79.9000 ;
	    RECT 183.1000 77.8000 183.4000 77.9000 ;
	    RECT 184.6000 77.9000 185.0000 79.9000 ;
	    RECT 184.6000 77.8000 184.9000 77.9000 ;
	    RECT 183.1000 77.5000 184.9000 77.8000 ;
	    RECT 183.1000 76.2000 183.4000 77.5000 ;
	    RECT 183.8000 76.4000 184.2000 77.2000 ;
	    RECT 186.5000 76.3000 186.9000 79.9000 ;
	    RECT 180.6000 75.9000 182.6000 76.2000 ;
	    RECT 179.9000 75.2000 180.2000 75.9000 ;
	    RECT 183.0000 75.8000 183.4000 76.2000 ;
	    RECT 181.8000 75.2000 182.2000 75.4000 ;
	    RECT 179.8000 74.9000 181.0000 75.2000 ;
	    RECT 181.8000 74.9000 182.6000 75.2000 ;
	    RECT 179.8000 74.8000 180.2000 74.9000 ;
	    RECT 179.0000 74.1000 179.4000 74.2000 ;
	    RECT 179.8000 74.1000 180.2000 74.2000 ;
	    RECT 179.0000 73.8000 180.2000 74.1000 ;
	    RECT 179.0000 73.4000 179.4000 73.8000 ;
	    RECT 177.7000 72.8000 178.6000 73.1000 ;
	    RECT 179.8000 72.8000 180.2000 73.2000 ;
	    RECT 180.7000 73.1000 181.0000 74.9000 ;
	    RECT 182.2000 74.8000 182.6000 74.9000 ;
	    RECT 181.4000 73.8000 181.8000 74.6000 ;
	    RECT 183.1000 74.2000 183.4000 75.8000 ;
	    RECT 185.4000 75.4000 185.8000 76.2000 ;
	    RECT 186.5000 75.9000 187.4000 76.3000 ;
	    RECT 184.2000 74.8000 185.0000 75.2000 ;
	    RECT 186.2000 74.8000 186.6000 75.6000 ;
	    RECT 187.0000 74.2000 187.3000 75.9000 ;
	    RECT 188.6000 75.8000 189.0000 76.6000 ;
	    RECT 183.1000 74.1000 183.9000 74.2000 ;
	    RECT 183.1000 73.9000 184.9000 74.1000 ;
	    RECT 183.6000 73.8000 184.9000 73.9000 ;
	    RECT 177.7000 71.1000 178.1000 72.8000 ;
	    RECT 179.9000 72.4000 180.3000 72.8000 ;
	    RECT 180.6000 71.1000 181.0000 73.1000 ;
	    RECT 183.6000 71.1000 184.0000 73.8000 ;
	    RECT 184.6000 73.2000 184.9000 73.8000 ;
	    RECT 187.0000 73.8000 187.4000 74.2000 ;
	    RECT 184.6000 72.8000 185.0000 73.2000 ;
	    RECT 187.0000 72.2000 187.3000 73.8000 ;
	    RECT 187.8000 73.1000 188.2000 73.2000 ;
	    RECT 189.4000 73.1000 189.8000 79.9000 ;
	    RECT 191.0000 75.6000 191.4000 79.9000 ;
	    RECT 193.1000 76.2000 193.5000 79.9000 ;
	    RECT 194.6000 76.8000 195.0000 77.2000 ;
	    RECT 194.6000 76.2000 194.9000 76.8000 ;
	    RECT 195.3000 76.2000 195.7000 79.9000 ;
	    RECT 197.7000 76.2000 198.1000 79.9000 ;
	    RECT 193.1000 75.9000 193.8000 76.2000 ;
	    RECT 191.0000 75.4000 193.0000 75.6000 ;
	    RECT 191.0000 75.3000 193.1000 75.4000 ;
	    RECT 192.7000 75.0000 193.1000 75.3000 ;
	    RECT 193.5000 75.2000 193.8000 75.9000 ;
	    RECT 194.2000 75.9000 194.9000 76.2000 ;
	    RECT 195.2000 75.9000 195.7000 76.2000 ;
	    RECT 197.4000 75.9000 198.1000 76.2000 ;
	    RECT 194.2000 75.8000 194.6000 75.9000 ;
	    RECT 192.0000 74.2000 192.4000 74.6000 ;
	    RECT 190.2000 73.4000 190.6000 74.2000 ;
	    RECT 191.8000 73.8000 192.3000 74.2000 ;
	    RECT 192.8000 73.5000 193.1000 75.0000 ;
	    RECT 193.4000 74.8000 193.8000 75.2000 ;
	    RECT 193.5000 74.2000 193.8000 74.8000 ;
	    RECT 195.2000 74.2000 195.5000 75.9000 ;
	    RECT 197.4000 75.2000 197.7000 75.9000 ;
	    RECT 199.8000 75.6000 200.2000 79.9000 ;
	    RECT 200.9000 76.3000 201.3000 79.9000 ;
	    RECT 200.9000 75.9000 201.8000 76.3000 ;
	    RECT 201.4000 75.8000 201.8000 75.9000 ;
	    RECT 203.0000 75.8000 203.4000 76.6000 ;
	    RECT 198.2000 75.4000 200.2000 75.6000 ;
	    RECT 198.1000 75.3000 200.2000 75.4000 ;
	    RECT 195.8000 74.4000 196.2000 75.2000 ;
	    RECT 197.4000 74.8000 197.8000 75.2000 ;
	    RECT 198.1000 75.0000 198.5000 75.3000 ;
	    RECT 193.4000 73.8000 193.8000 74.2000 ;
	    RECT 194.2000 73.8000 195.5000 74.2000 ;
	    RECT 196.6000 74.1000 197.0000 74.2000 ;
	    RECT 197.4000 74.1000 197.7000 74.8000 ;
	    RECT 196.2000 73.8000 197.7000 74.1000 ;
	    RECT 191.9000 73.2000 193.1000 73.5000 ;
	    RECT 187.8000 72.8000 189.8000 73.1000 ;
	    RECT 187.8000 72.4000 188.2000 72.8000 ;
	    RECT 187.0000 71.1000 187.4000 72.2000 ;
	    RECT 188.9000 71.1000 189.3000 72.8000 ;
	    RECT 191.0000 72.4000 191.4000 73.2000 ;
	    RECT 191.9000 72.1000 192.2000 73.2000 ;
	    RECT 193.5000 73.1000 193.8000 73.8000 ;
	    RECT 194.3000 73.1000 194.6000 73.8000 ;
	    RECT 196.2000 73.6000 196.6000 73.8000 ;
	    RECT 195.1000 73.1000 196.9000 73.3000 ;
	    RECT 197.4000 73.1000 197.7000 73.8000 ;
	    RECT 198.1000 73.5000 198.4000 75.0000 ;
	    RECT 200.6000 74.8000 201.0000 75.6000 ;
	    RECT 198.8000 74.2000 199.2000 74.6000 ;
	    RECT 201.4000 74.2000 201.7000 75.8000 ;
	    RECT 198.9000 73.8000 199.4000 74.2000 ;
	    RECT 201.4000 73.8000 201.8000 74.2000 ;
	    RECT 198.1000 73.2000 199.3000 73.5000 ;
	    RECT 191.8000 71.1000 192.2000 72.1000 ;
	    RECT 193.4000 71.1000 193.8000 73.1000 ;
	    RECT 194.2000 71.1000 194.6000 73.1000 ;
	    RECT 195.0000 73.0000 197.0000 73.1000 ;
	    RECT 195.0000 71.1000 195.4000 73.0000 ;
	    RECT 196.6000 71.1000 197.0000 73.0000 ;
	    RECT 197.4000 71.1000 197.8000 73.1000 ;
	    RECT 199.0000 72.1000 199.3000 73.2000 ;
	    RECT 199.8000 72.4000 200.2000 73.2000 ;
	    RECT 201.4000 72.1000 201.7000 73.8000 ;
	    RECT 202.2000 72.4000 202.6000 73.2000 ;
	    RECT 203.8000 73.1000 204.2000 79.9000 ;
	    RECT 205.4000 75.9000 205.8000 79.9000 ;
	    RECT 206.2000 76.2000 206.6000 79.9000 ;
	    RECT 207.8000 76.2000 208.2000 79.9000 ;
	    RECT 206.2000 75.9000 208.2000 76.2000 ;
	    RECT 205.5000 75.2000 205.8000 75.9000 ;
	    RECT 210.2000 75.7000 210.6000 79.9000 ;
	    RECT 212.4000 78.2000 212.8000 79.9000 ;
	    RECT 211.8000 77.9000 212.8000 78.2000 ;
	    RECT 214.6000 77.9000 215.0000 79.9000 ;
	    RECT 216.7000 77.9000 217.3000 79.9000 ;
	    RECT 211.8000 77.5000 212.2000 77.9000 ;
	    RECT 214.6000 77.6000 214.9000 77.9000 ;
	    RECT 213.5000 77.3000 215.3000 77.6000 ;
	    RECT 216.6000 77.5000 217.0000 77.9000 ;
	    RECT 213.5000 77.2000 213.9000 77.3000 ;
	    RECT 214.9000 77.2000 215.3000 77.3000 ;
	    RECT 211.8000 76.5000 212.2000 76.6000 ;
	    RECT 214.1000 76.5000 214.5000 76.6000 ;
	    RECT 211.8000 76.2000 214.5000 76.5000 ;
	    RECT 214.8000 76.5000 215.9000 76.8000 ;
	    RECT 214.8000 75.9000 215.1000 76.5000 ;
	    RECT 215.5000 76.4000 215.9000 76.5000 ;
	    RECT 216.7000 76.6000 217.4000 77.0000 ;
	    RECT 216.7000 76.1000 217.0000 76.6000 ;
	    RECT 212.7000 75.7000 215.1000 75.9000 ;
	    RECT 210.2000 75.6000 215.1000 75.7000 ;
	    RECT 215.8000 75.8000 217.0000 76.1000 ;
	    RECT 210.2000 75.5000 213.1000 75.6000 ;
	    RECT 210.2000 75.4000 213.0000 75.5000 ;
	    RECT 207.4000 75.2000 207.8000 75.4000 ;
	    RECT 205.4000 74.9000 206.6000 75.2000 ;
	    RECT 207.4000 74.9000 208.2000 75.2000 ;
	    RECT 213.4000 75.1000 213.8000 75.2000 ;
	    RECT 205.4000 74.8000 205.8000 74.9000 ;
	    RECT 206.2000 74.8000 206.6000 74.9000 ;
	    RECT 207.8000 74.8000 208.2000 74.9000 ;
	    RECT 211.3000 74.8000 213.8000 75.1000 ;
	    RECT 204.6000 73.4000 205.0000 74.2000 ;
	    RECT 203.3000 72.8000 204.2000 73.1000 ;
	    RECT 205.4000 72.8000 205.8000 73.2000 ;
	    RECT 206.3000 73.1000 206.6000 74.8000 ;
	    RECT 211.3000 74.7000 211.7000 74.8000 ;
	    RECT 212.6000 74.7000 213.0000 74.8000 ;
	    RECT 207.0000 73.8000 207.4000 74.6000 ;
	    RECT 212.1000 74.2000 212.5000 74.3000 ;
	    RECT 215.8000 74.2000 216.1000 75.8000 ;
	    RECT 219.0000 75.6000 219.4000 79.9000 ;
	    RECT 217.3000 75.3000 219.4000 75.6000 ;
	    RECT 217.3000 75.2000 217.7000 75.3000 ;
	    RECT 218.1000 74.9000 218.5000 75.0000 ;
	    RECT 216.6000 74.6000 218.5000 74.9000 ;
	    RECT 216.6000 74.5000 217.0000 74.6000 ;
	    RECT 210.6000 73.9000 216.1000 74.2000 ;
	    RECT 210.6000 73.8000 211.4000 73.9000 ;
	    RECT 199.0000 71.1000 199.4000 72.1000 ;
	    RECT 201.4000 71.1000 201.8000 72.1000 ;
	    RECT 203.3000 71.1000 203.7000 72.8000 ;
	    RECT 205.5000 72.4000 205.9000 72.8000 ;
	    RECT 206.2000 71.1000 206.6000 73.1000 ;
	    RECT 210.2000 71.1000 210.6000 73.5000 ;
	    RECT 212.7000 72.8000 213.0000 73.9000 ;
	    RECT 215.5000 73.8000 215.9000 73.9000 ;
	    RECT 219.0000 73.6000 219.4000 75.3000 ;
	    RECT 217.5000 73.3000 219.4000 73.6000 ;
	    RECT 217.5000 73.2000 217.9000 73.3000 ;
	    RECT 211.8000 72.1000 212.2000 72.5000 ;
	    RECT 212.6000 72.4000 213.0000 72.8000 ;
	    RECT 213.5000 72.7000 213.9000 72.8000 ;
	    RECT 213.5000 72.4000 214.9000 72.7000 ;
	    RECT 214.6000 72.1000 214.9000 72.4000 ;
	    RECT 216.6000 72.1000 217.0000 72.5000 ;
	    RECT 211.8000 71.8000 212.8000 72.1000 ;
	    RECT 212.4000 71.1000 212.8000 71.8000 ;
	    RECT 214.6000 71.1000 215.0000 72.1000 ;
	    RECT 216.6000 71.8000 217.3000 72.1000 ;
	    RECT 216.7000 71.1000 217.3000 71.8000 ;
	    RECT 219.0000 71.1000 219.4000 73.3000 ;
	    RECT 219.8000 71.1000 220.2000 79.9000 ;
	    RECT 220.6000 73.1000 221.0000 73.2000 ;
	    RECT 221.4000 73.1000 221.8000 73.2000 ;
	    RECT 220.6000 72.8000 221.8000 73.1000 ;
	    RECT 220.6000 72.4000 221.0000 72.8000 ;
	    RECT 221.4000 72.4000 221.8000 72.8000 ;
	    RECT 222.2000 71.1000 222.6000 79.9000 ;
	    RECT 223.0000 77.1000 223.4000 79.9000 ;
	    RECT 223.8000 77.1000 224.2000 77.2000 ;
	    RECT 223.0000 76.8000 224.2000 77.1000 ;
	    RECT 223.0000 71.1000 223.4000 76.8000 ;
	    RECT 225.9000 76.2000 226.3000 79.9000 ;
	    RECT 228.6000 77.8000 229.0000 79.9000 ;
	    RECT 230.2000 77.9000 230.6000 79.9000 ;
	    RECT 232.3000 79.2000 232.7000 79.9000 ;
	    RECT 231.8000 78.8000 232.7000 79.2000 ;
	    RECT 230.2000 77.8000 230.5000 77.9000 ;
	    RECT 228.6000 77.5000 230.5000 77.8000 ;
	    RECT 226.6000 77.1000 227.0000 77.2000 ;
	    RECT 228.6000 77.1000 228.9000 77.5000 ;
	    RECT 226.6000 76.8000 228.9000 77.1000 ;
	    RECT 226.7000 76.2000 227.0000 76.8000 ;
	    RECT 229.4000 76.4000 229.8000 77.2000 ;
	    RECT 230.2000 76.2000 230.5000 77.5000 ;
	    RECT 232.3000 76.2000 232.7000 78.8000 ;
	    RECT 233.0000 76.8000 233.4000 77.2000 ;
	    RECT 233.1000 76.2000 233.4000 76.8000 ;
	    RECT 234.6000 76.8000 235.0000 77.2000 ;
	    RECT 234.6000 76.2000 234.9000 76.8000 ;
	    RECT 235.3000 76.2000 235.7000 79.9000 ;
	    RECT 238.7000 76.3000 239.1000 79.9000 ;
	    RECT 225.9000 75.9000 226.4000 76.2000 ;
	    RECT 226.7000 75.9000 227.4000 76.2000 ;
	    RECT 225.4000 74.4000 225.8000 75.2000 ;
	    RECT 226.1000 74.2000 226.4000 75.9000 ;
	    RECT 227.0000 75.8000 227.4000 75.9000 ;
	    RECT 227.8000 75.4000 228.2000 76.2000 ;
	    RECT 230.2000 75.8000 230.6000 76.2000 ;
	    RECT 232.3000 75.9000 232.8000 76.2000 ;
	    RECT 233.1000 75.9000 233.8000 76.2000 ;
	    RECT 227.0000 74.8000 227.4000 75.2000 ;
	    RECT 228.6000 74.8000 229.4000 75.2000 ;
	    RECT 227.0000 74.2000 227.3000 74.8000 ;
	    RECT 230.2000 74.2000 230.5000 75.8000 ;
	    RECT 231.8000 74.4000 232.2000 75.2000 ;
	    RECT 232.5000 74.2000 232.8000 75.9000 ;
	    RECT 233.4000 75.8000 233.8000 75.9000 ;
	    RECT 234.2000 75.9000 234.9000 76.2000 ;
	    RECT 235.2000 75.9000 235.7000 76.2000 ;
	    RECT 238.2000 75.9000 239.1000 76.3000 ;
	    RECT 234.2000 75.8000 234.6000 75.9000 ;
	    RECT 233.4000 75.1000 233.7000 75.8000 ;
	    RECT 235.2000 75.1000 235.5000 75.9000 ;
	    RECT 233.4000 74.8000 235.5000 75.1000 ;
	    RECT 235.2000 74.2000 235.5000 74.8000 ;
	    RECT 235.8000 75.1000 236.2000 75.2000 ;
	    RECT 238.3000 75.1000 238.6000 75.9000 ;
	    RECT 235.8000 74.8000 238.6000 75.1000 ;
	    RECT 235.8000 74.4000 236.2000 74.8000 ;
	    RECT 238.3000 74.2000 238.6000 74.8000 ;
	    RECT 223.8000 74.1000 224.2000 74.2000 ;
	    RECT 224.6000 74.1000 225.0000 74.2000 ;
	    RECT 223.8000 73.8000 225.4000 74.1000 ;
	    RECT 226.1000 73.8000 227.4000 74.2000 ;
	    RECT 229.7000 74.1000 230.5000 74.2000 ;
	    RECT 229.6000 73.9000 230.5000 74.1000 ;
	    RECT 231.0000 74.1000 231.4000 74.2000 ;
	    RECT 225.0000 73.6000 225.4000 73.8000 ;
	    RECT 223.8000 72.4000 224.2000 73.2000 ;
	    RECT 224.7000 73.1000 226.5000 73.3000 ;
	    RECT 227.0000 73.1000 227.3000 73.8000 ;
	    RECT 224.6000 73.0000 226.6000 73.1000 ;
	    RECT 224.6000 71.1000 225.0000 73.0000 ;
	    RECT 226.2000 71.1000 226.6000 73.0000 ;
	    RECT 227.0000 71.1000 227.4000 73.1000 ;
	    RECT 229.6000 71.1000 230.0000 73.9000 ;
	    RECT 231.0000 73.8000 231.8000 74.1000 ;
	    RECT 232.5000 73.8000 233.8000 74.2000 ;
	    RECT 234.2000 73.8000 235.5000 74.2000 ;
	    RECT 236.6000 74.1000 237.0000 74.2000 ;
	    RECT 236.2000 73.8000 237.0000 74.1000 ;
	    RECT 238.2000 73.8000 238.6000 74.2000 ;
	    RECT 239.0000 74.8000 239.4000 75.6000 ;
	    RECT 239.0000 74.2000 239.3000 74.8000 ;
	    RECT 239.0000 73.8000 239.4000 74.2000 ;
	    RECT 231.4000 73.6000 231.8000 73.8000 ;
	    RECT 231.1000 73.1000 232.9000 73.3000 ;
	    RECT 233.4000 73.1000 233.7000 73.8000 ;
	    RECT 234.3000 73.1000 234.6000 73.8000 ;
	    RECT 236.2000 73.6000 236.6000 73.8000 ;
	    RECT 235.1000 73.1000 236.9000 73.3000 ;
	    RECT 231.0000 73.0000 233.0000 73.1000 ;
	    RECT 231.0000 71.1000 231.4000 73.0000 ;
	    RECT 232.6000 71.1000 233.0000 73.0000 ;
	    RECT 233.4000 71.1000 233.8000 73.1000 ;
	    RECT 234.2000 71.1000 234.6000 73.1000 ;
	    RECT 235.0000 73.0000 237.0000 73.1000 ;
	    RECT 235.0000 71.1000 235.4000 73.0000 ;
	    RECT 236.6000 71.1000 237.0000 73.0000 ;
	    RECT 237.4000 72.4000 237.8000 73.2000 ;
	    RECT 238.3000 72.1000 238.6000 73.8000 ;
	    RECT 238.2000 71.1000 238.6000 72.1000 ;
	    RECT 239.8000 71.1000 240.2000 79.9000 ;
	    RECT 240.6000 74.8000 241.0000 75.2000 ;
	    RECT 240.6000 74.1000 240.9000 74.8000 ;
	    RECT 241.4000 74.1000 241.8000 74.2000 ;
	    RECT 240.6000 73.8000 241.8000 74.1000 ;
	    RECT 241.4000 73.4000 241.8000 73.8000 ;
	    RECT 240.6000 72.4000 241.0000 73.2000 ;
	    RECT 242.2000 73.1000 242.6000 79.9000 ;
	    RECT 243.0000 75.8000 243.4000 76.6000 ;
	    RECT 245.1000 76.3000 245.5000 79.9000 ;
	    RECT 244.6000 75.9000 245.5000 76.3000 ;
	    RECT 246.2000 76.2000 246.6000 79.9000 ;
	    RECT 247.1000 76.2000 247.5000 76.3000 ;
	    RECT 246.2000 75.9000 247.5000 76.2000 ;
	    RECT 248.4000 75.9000 249.2000 79.9000 ;
	    RECT 250.2000 76.2000 250.6000 76.3000 ;
	    RECT 251.0000 76.2000 251.4000 79.9000 ;
	    RECT 251.8000 77.9000 252.2000 79.9000 ;
	    RECT 251.9000 77.8000 252.2000 77.9000 ;
	    RECT 253.4000 77.9000 253.8000 79.9000 ;
	    RECT 253.4000 77.8000 253.7000 77.9000 ;
	    RECT 251.9000 77.5000 253.7000 77.8000 ;
	    RECT 251.9000 76.2000 252.2000 77.5000 ;
	    RECT 252.6000 76.4000 253.0000 77.2000 ;
	    RECT 250.2000 75.9000 251.4000 76.2000 ;
	    RECT 244.7000 74.2000 245.0000 75.9000 ;
	    RECT 247.7000 75.2000 248.1000 75.3000 ;
	    RECT 248.7000 75.2000 249.0000 75.9000 ;
	    RECT 251.8000 75.8000 252.2000 76.2000 ;
	    RECT 247.3000 74.9000 248.1000 75.2000 ;
	    RECT 247.3000 74.8000 247.7000 74.9000 ;
	    RECT 248.6000 74.8000 249.0000 75.2000 ;
	    RECT 248.0000 74.3000 248.4000 74.4000 ;
	    RECT 247.0000 74.2000 248.4000 74.3000 ;
	    RECT 244.6000 74.1000 245.0000 74.2000 ;
	    RECT 246.2000 74.1000 248.4000 74.2000 ;
	    RECT 244.6000 74.0000 248.4000 74.1000 ;
	    RECT 248.7000 74.2000 249.0000 74.8000 ;
	    RECT 251.9000 74.2000 252.2000 75.8000 ;
	    RECT 253.0000 74.8000 253.8000 75.2000 ;
	    RECT 254.2000 75.1000 254.6000 76.2000 ;
	    RECT 255.0000 75.8000 255.4000 76.6000 ;
	    RECT 255.8000 75.1000 256.2000 79.9000 ;
	    RECT 257.8000 76.8000 258.2000 77.2000 ;
	    RECT 257.8000 76.2000 258.1000 76.8000 ;
	    RECT 258.5000 76.2000 258.9000 79.9000 ;
	    RECT 261.7000 79.2000 262.1000 79.9000 ;
	    RECT 261.7000 78.8000 262.6000 79.2000 ;
	    RECT 261.0000 76.8000 261.4000 77.2000 ;
	    RECT 261.0000 76.2000 261.3000 76.8000 ;
	    RECT 261.7000 76.2000 262.1000 78.8000 ;
	    RECT 265.1000 76.3000 265.5000 79.9000 ;
	    RECT 257.4000 75.9000 258.1000 76.2000 ;
	    RECT 258.4000 75.9000 258.9000 76.2000 ;
	    RECT 260.6000 75.9000 261.3000 76.2000 ;
	    RECT 261.6000 75.9000 262.1000 76.2000 ;
	    RECT 264.6000 75.9000 265.5000 76.3000 ;
	    RECT 257.4000 75.8000 257.8000 75.9000 ;
	    RECT 254.2000 74.8000 256.2000 75.1000 ;
	    RECT 256.6000 75.1000 257.0000 75.2000 ;
	    RECT 258.4000 75.1000 258.7000 75.9000 ;
	    RECT 260.6000 75.8000 261.0000 75.9000 ;
	    RECT 256.6000 74.8000 258.7000 75.1000 ;
	    RECT 244.6000 73.9000 247.3000 74.0000 ;
	    RECT 248.7000 73.9000 249.2000 74.2000 ;
	    RECT 244.6000 73.8000 247.0000 73.9000 ;
	    RECT 242.2000 72.8000 243.1000 73.1000 ;
	    RECT 242.7000 72.2000 243.1000 72.8000 ;
	    RECT 243.8000 72.4000 244.2000 73.2000 ;
	    RECT 242.2000 71.8000 243.1000 72.2000 ;
	    RECT 244.7000 72.1000 245.0000 73.8000 ;
	    RECT 247.1000 73.4000 247.5000 73.5000 ;
	    RECT 242.7000 71.1000 243.1000 71.8000 ;
	    RECT 244.6000 71.1000 245.0000 72.1000 ;
	    RECT 246.2000 73.1000 247.5000 73.4000 ;
	    RECT 247.8000 73.2000 248.6000 73.6000 ;
	    RECT 246.2000 71.1000 246.6000 73.1000 ;
	    RECT 248.9000 72.9000 249.2000 73.9000 ;
	    RECT 249.6000 73.8000 250.0000 74.2000 ;
	    RECT 251.9000 74.1000 252.7000 74.2000 ;
	    RECT 251.9000 73.9000 252.8000 74.1000 ;
	    RECT 249.6000 73.6000 249.9000 73.8000 ;
	    RECT 249.5000 73.2000 249.9000 73.6000 ;
	    RECT 250.2000 73.4000 250.6000 73.5000 ;
	    RECT 250.2000 73.1000 251.4000 73.4000 ;
	    RECT 248.4000 72.2000 249.2000 72.9000 ;
	    RECT 247.8000 71.8000 249.2000 72.2000 ;
	    RECT 248.4000 71.1000 249.2000 71.8000 ;
	    RECT 251.0000 71.1000 251.4000 73.1000 ;
	    RECT 252.4000 71.1000 252.8000 73.9000 ;
	    RECT 255.8000 73.1000 256.2000 74.8000 ;
	    RECT 258.4000 74.2000 258.7000 74.8000 ;
	    RECT 259.0000 74.4000 259.4000 75.2000 ;
	    RECT 261.6000 74.2000 261.9000 75.9000 ;
	    RECT 262.2000 75.1000 262.6000 75.2000 ;
	    RECT 264.7000 75.1000 265.0000 75.9000 ;
	    RECT 262.2000 74.8000 265.0000 75.1000 ;
	    RECT 265.4000 74.8000 265.8000 75.6000 ;
	    RECT 262.2000 74.4000 262.6000 74.8000 ;
	    RECT 264.7000 74.2000 265.0000 74.8000 ;
	    RECT 257.4000 73.8000 258.7000 74.2000 ;
	    RECT 259.8000 74.1000 260.2000 74.2000 ;
	    RECT 259.4000 73.8000 260.2000 74.1000 ;
	    RECT 260.6000 73.8000 261.9000 74.2000 ;
	    RECT 263.0000 74.1000 263.4000 74.2000 ;
	    RECT 262.6000 73.8000 263.4000 74.1000 ;
	    RECT 264.6000 73.8000 265.0000 74.2000 ;
	    RECT 257.5000 73.1000 257.8000 73.8000 ;
	    RECT 259.4000 73.6000 259.8000 73.8000 ;
	    RECT 258.3000 73.1000 260.1000 73.3000 ;
	    RECT 260.7000 73.1000 261.0000 73.8000 ;
	    RECT 262.6000 73.6000 263.0000 73.8000 ;
	    RECT 261.5000 73.1000 263.3000 73.3000 ;
	    RECT 255.3000 72.8000 256.2000 73.1000 ;
	    RECT 255.3000 71.1000 255.7000 72.8000 ;
	    RECT 257.4000 71.1000 257.8000 73.1000 ;
	    RECT 258.2000 73.0000 260.2000 73.1000 ;
	    RECT 258.2000 71.1000 258.6000 73.0000 ;
	    RECT 259.8000 71.1000 260.2000 73.0000 ;
	    RECT 260.6000 71.1000 261.0000 73.1000 ;
	    RECT 261.4000 73.0000 263.4000 73.1000 ;
	    RECT 261.4000 71.1000 261.8000 73.0000 ;
	    RECT 263.0000 71.1000 263.4000 73.0000 ;
	    RECT 264.7000 72.1000 265.0000 73.8000 ;
	    RECT 267.0000 73.1000 267.4000 79.9000 ;
	    RECT 267.8000 75.8000 268.2000 76.6000 ;
	    RECT 267.0000 72.8000 267.9000 73.1000 ;
	    RECT 264.6000 71.1000 265.0000 72.1000 ;
	    RECT 267.5000 72.2000 267.9000 72.8000 ;
	    RECT 267.5000 71.8000 268.2000 72.2000 ;
	    RECT 267.5000 71.1000 267.9000 71.8000 ;
	    RECT 268.6000 71.1000 269.0000 79.9000 ;
	    RECT 269.4000 72.4000 269.8000 73.2000 ;
	    RECT 1.4000 65.1000 1.8000 69.9000 ;
	    RECT 3.5000 68.2000 3.9000 69.9000 ;
	    RECT 3.0000 67.9000 3.9000 68.2000 ;
	    RECT 5.4000 68.9000 5.8000 69.9000 ;
	    RECT 3.0000 67.1000 3.4000 67.9000 ;
	    RECT 5.4000 67.2000 5.7000 68.9000 ;
	    RECT 7.1000 68.2000 7.5000 68.6000 ;
	    RECT 7.0000 67.8000 7.4000 68.2000 ;
	    RECT 7.8000 67.9000 8.2000 69.9000 ;
	    RECT 10.2000 67.9000 10.6000 69.9000 ;
	    RECT 11.0000 68.0000 11.4000 69.9000 ;
	    RECT 12.6000 68.0000 13.0000 69.9000 ;
	    RECT 11.0000 67.9000 13.0000 68.0000 ;
	    RECT 14.2000 68.8000 14.6000 69.9000 ;
	    RECT 4.6000 67.1000 5.0000 67.2000 ;
	    RECT 3.0000 66.8000 5.0000 67.1000 ;
	    RECT 5.4000 67.1000 5.8000 67.2000 ;
	    RECT 7.0000 67.1000 7.3000 67.8000 ;
	    RECT 5.4000 66.8000 7.3000 67.1000 ;
	    RECT 2.2000 65.8000 2.6000 66.2000 ;
	    RECT 2.2000 65.1000 2.5000 65.8000 ;
	    RECT 1.4000 64.8000 2.5000 65.1000 ;
	    RECT 1.4000 61.1000 1.8000 64.8000 ;
	    RECT 3.0000 61.1000 3.4000 66.8000 ;
	    RECT 3.8000 66.1000 4.2000 66.2000 ;
	    RECT 4.6000 66.1000 5.0000 66.2000 ;
	    RECT 3.8000 65.8000 5.0000 66.1000 ;
	    RECT 4.6000 65.4000 5.0000 65.8000 ;
	    RECT 3.8000 64.4000 4.2000 65.2000 ;
	    RECT 5.4000 65.1000 5.7000 66.8000 ;
	    RECT 7.9000 66.2000 8.2000 67.9000 ;
	    RECT 10.3000 67.2000 10.6000 67.9000 ;
	    RECT 11.1000 67.7000 12.9000 67.9000 ;
	    RECT 12.2000 67.2000 12.6000 67.4000 ;
	    RECT 14.2000 67.2000 14.5000 68.8000 ;
	    RECT 15.0000 67.8000 15.4000 68.6000 ;
	    RECT 17.4000 67.9000 17.8000 69.9000 ;
	    RECT 18.1000 68.2000 18.5000 68.6000 ;
	    RECT 19.3000 68.2000 19.7000 69.9000 ;
	    RECT 8.6000 66.4000 9.0000 67.2000 ;
	    RECT 10.2000 66.8000 11.5000 67.2000 ;
	    RECT 12.2000 66.9000 13.0000 67.2000 ;
	    RECT 12.6000 66.8000 13.0000 66.9000 ;
	    RECT 14.2000 66.8000 14.6000 67.2000 ;
	    RECT 7.0000 66.1000 7.4000 66.2000 ;
	    RECT 7.8000 66.1000 8.2000 66.2000 ;
	    RECT 9.4000 66.1000 9.8000 66.2000 ;
	    RECT 7.0000 65.8000 8.2000 66.1000 ;
	    RECT 9.0000 65.8000 9.8000 66.1000 ;
	    RECT 7.1000 65.1000 7.4000 65.8000 ;
	    RECT 9.0000 65.6000 9.4000 65.8000 ;
	    RECT 10.2000 65.1000 10.6000 65.2000 ;
	    RECT 11.2000 65.1000 11.5000 66.8000 ;
	    RECT 11.8000 65.8000 12.2000 66.6000 ;
	    RECT 12.6000 66.1000 13.0000 66.2000 ;
	    RECT 13.4000 66.1000 13.8000 66.2000 ;
	    RECT 12.6000 65.8000 13.8000 66.1000 ;
	    RECT 13.4000 65.4000 13.8000 65.8000 ;
	    RECT 14.2000 65.1000 14.5000 66.8000 ;
	    RECT 16.6000 66.4000 17.0000 67.2000 ;
	    RECT 15.8000 66.1000 16.2000 66.2000 ;
	    RECT 17.4000 66.1000 17.7000 67.9000 ;
	    RECT 18.2000 67.8000 18.6000 68.2000 ;
	    RECT 19.3000 67.9000 20.2000 68.2000 ;
	    RECT 19.0000 67.1000 19.4000 67.2000 ;
	    RECT 19.8000 67.1000 20.2000 67.9000 ;
	    RECT 23.0000 67.9000 23.4000 69.9000 ;
	    RECT 25.4000 68.9000 25.8000 69.9000 ;
	    RECT 23.7000 68.2000 24.1000 68.6000 ;
	    RECT 19.0000 66.8000 20.2000 67.1000 ;
	    RECT 20.6000 67.1000 21.0000 67.6000 ;
	    RECT 21.4000 67.1000 21.8000 67.2000 ;
	    RECT 20.6000 66.8000 21.8000 67.1000 ;
	    RECT 18.2000 66.1000 18.6000 66.2000 ;
	    RECT 15.8000 65.8000 16.6000 66.1000 ;
	    RECT 17.4000 65.8000 18.6000 66.1000 ;
	    RECT 16.2000 65.6000 16.6000 65.8000 ;
	    RECT 18.2000 65.1000 18.5000 65.8000 ;
	    RECT 4.9000 64.7000 5.8000 65.1000 ;
	    RECT 4.9000 61.1000 5.3000 64.7000 ;
	    RECT 7.0000 61.1000 7.4000 65.1000 ;
	    RECT 7.8000 64.8000 9.8000 65.1000 ;
	    RECT 10.2000 64.8000 10.9000 65.1000 ;
	    RECT 11.2000 64.8000 11.7000 65.1000 ;
	    RECT 7.8000 61.1000 8.2000 64.8000 ;
	    RECT 9.4000 61.1000 9.8000 64.8000 ;
	    RECT 10.6000 64.2000 10.9000 64.8000 ;
	    RECT 10.6000 63.8000 11.0000 64.2000 ;
	    RECT 11.3000 61.1000 11.7000 64.8000 ;
	    RECT 13.7000 64.7000 14.6000 65.1000 ;
	    RECT 15.8000 64.8000 17.8000 65.1000 ;
	    RECT 13.7000 61.1000 14.1000 64.7000 ;
	    RECT 15.8000 61.1000 16.2000 64.8000 ;
	    RECT 17.4000 61.1000 17.8000 64.8000 ;
	    RECT 18.2000 61.1000 18.6000 65.1000 ;
	    RECT 19.0000 64.4000 19.4000 65.2000 ;
	    RECT 19.8000 61.1000 20.2000 66.8000 ;
	    RECT 22.2000 66.4000 22.6000 67.2000 ;
	    RECT 20.6000 66.1000 21.0000 66.2000 ;
	    RECT 21.4000 66.1000 21.8000 66.2000 ;
	    RECT 23.0000 66.1000 23.3000 67.9000 ;
	    RECT 23.8000 67.8000 24.2000 68.2000 ;
	    RECT 24.6000 67.8000 25.0000 68.6000 ;
	    RECT 25.5000 67.2000 25.8000 68.9000 ;
	    RECT 27.1000 68.2000 27.5000 68.6000 ;
	    RECT 27.0000 67.8000 27.4000 68.2000 ;
	    RECT 27.8000 67.9000 28.2000 69.9000 ;
	    RECT 31.5000 69.2000 31.9000 69.9000 ;
	    RECT 31.0000 68.8000 31.9000 69.2000 ;
	    RECT 31.5000 68.2000 31.9000 68.8000 ;
	    RECT 25.4000 66.8000 25.8000 67.2000 ;
	    RECT 23.8000 66.1000 24.2000 66.2000 ;
	    RECT 20.6000 65.8000 22.2000 66.1000 ;
	    RECT 23.0000 65.8000 24.2000 66.1000 ;
	    RECT 24.6000 66.1000 25.0000 66.2000 ;
	    RECT 25.5000 66.1000 25.8000 66.8000 ;
	    RECT 24.6000 65.8000 25.8000 66.1000 ;
	    RECT 21.8000 65.6000 22.2000 65.8000 ;
	    RECT 23.8000 65.1000 24.1000 65.8000 ;
	    RECT 25.5000 65.1000 25.8000 65.8000 ;
	    RECT 26.2000 65.4000 26.6000 66.2000 ;
	    RECT 27.0000 66.1000 27.4000 66.2000 ;
	    RECT 27.9000 66.1000 28.2000 67.9000 ;
	    RECT 31.0000 67.9000 31.9000 68.2000 ;
	    RECT 28.6000 66.4000 29.0000 67.2000 ;
	    RECT 30.2000 67.1000 30.6000 67.6000 ;
	    RECT 29.4000 66.8000 30.6000 67.1000 ;
	    RECT 29.4000 66.2000 29.7000 66.8000 ;
	    RECT 29.4000 66.1000 29.8000 66.2000 ;
	    RECT 27.0000 65.8000 28.2000 66.1000 ;
	    RECT 29.0000 65.8000 29.8000 66.1000 ;
	    RECT 27.1000 65.1000 27.4000 65.8000 ;
	    RECT 29.0000 65.6000 29.4000 65.8000 ;
	    RECT 21.4000 64.8000 23.4000 65.1000 ;
	    RECT 21.4000 61.1000 21.8000 64.8000 ;
	    RECT 23.0000 61.1000 23.4000 64.8000 ;
	    RECT 23.8000 61.1000 24.2000 65.1000 ;
	    RECT 25.4000 64.7000 26.3000 65.1000 ;
	    RECT 25.9000 61.1000 26.3000 64.7000 ;
	    RECT 27.0000 61.1000 27.4000 65.1000 ;
	    RECT 27.8000 64.8000 29.8000 65.1000 ;
	    RECT 27.8000 61.1000 28.2000 64.8000 ;
	    RECT 29.4000 61.1000 29.8000 64.8000 ;
	    RECT 31.0000 61.1000 31.4000 67.9000 ;
	    RECT 32.6000 67.1000 33.0000 69.9000 ;
	    RECT 33.4000 67.8000 33.8000 68.6000 ;
	    RECT 34.5000 68.2000 34.9000 69.9000 ;
	    RECT 36.6000 69.6000 38.6000 69.9000 ;
	    RECT 34.5000 67.9000 35.4000 68.2000 ;
	    RECT 36.6000 67.9000 37.0000 69.6000 ;
	    RECT 37.4000 67.9000 37.8000 69.3000 ;
	    RECT 38.2000 68.0000 38.6000 69.6000 ;
	    RECT 39.8000 68.0000 40.2000 69.9000 ;
	    RECT 38.2000 67.9000 40.2000 68.0000 ;
	    RECT 32.6000 66.8000 34.5000 67.1000 ;
	    RECT 31.8000 64.4000 32.2000 65.2000 ;
	    RECT 32.6000 65.1000 33.0000 66.8000 ;
	    RECT 34.2000 66.2000 34.5000 66.8000 ;
	    RECT 34.2000 65.8000 34.6000 66.2000 ;
	    RECT 34.2000 65.1000 34.6000 65.2000 ;
	    RECT 32.6000 64.8000 34.6000 65.1000 ;
	    RECT 32.6000 61.1000 33.0000 64.8000 ;
	    RECT 34.2000 64.4000 34.6000 64.8000 ;
	    RECT 35.0000 65.1000 35.4000 67.9000 ;
	    RECT 35.8000 66.8000 36.2000 67.6000 ;
	    RECT 37.4000 67.2000 37.7000 67.9000 ;
	    RECT 38.3000 67.7000 40.1000 67.9000 ;
	    RECT 39.4000 67.2000 39.8000 67.4000 ;
	    RECT 41.2000 67.2000 41.6000 69.9000 ;
	    RECT 44.1000 68.2000 44.5000 69.9000 ;
	    RECT 42.2000 67.8000 42.6000 68.2000 ;
	    RECT 44.1000 67.9000 45.0000 68.2000 ;
	    RECT 36.6000 66.4000 37.0000 67.2000 ;
	    RECT 37.4000 66.9000 38.6000 67.2000 ;
	    RECT 39.4000 66.9000 40.2000 67.2000 ;
	    RECT 41.2000 67.1000 41.8000 67.2000 ;
	    RECT 42.2000 67.1000 42.5000 67.8000 ;
	    RECT 38.2000 66.8000 38.6000 66.9000 ;
	    RECT 39.8000 66.8000 40.2000 66.9000 ;
	    RECT 40.7000 66.8000 42.5000 67.1000 ;
	    RECT 37.4000 65.8000 37.8000 66.6000 ;
	    RECT 38.3000 65.1000 38.6000 66.8000 ;
	    RECT 39.0000 65.8000 39.4000 66.6000 ;
	    RECT 40.7000 65.2000 41.0000 66.8000 ;
	    RECT 41.8000 65.8000 42.6000 66.2000 ;
	    RECT 44.6000 66.1000 45.0000 67.9000 ;
	    RECT 45.4000 66.8000 45.8000 67.6000 ;
	    RECT 43.0000 65.8000 45.0000 66.1000 ;
	    RECT 35.0000 64.8000 36.1000 65.1000 ;
	    RECT 35.0000 61.1000 35.4000 64.8000 ;
	    RECT 35.8000 64.2000 36.1000 64.8000 ;
	    RECT 35.8000 63.8000 36.2000 64.2000 ;
	    RECT 37.9000 61.1000 38.9000 65.1000 ;
	    RECT 40.6000 64.8000 41.0000 65.2000 ;
	    RECT 43.0000 64.8000 43.4000 65.8000 ;
	    RECT 40.7000 63.5000 41.0000 64.8000 ;
	    RECT 41.4000 64.1000 41.8000 64.6000 ;
	    RECT 43.8000 64.4000 44.2000 65.2000 ;
	    RECT 43.0000 64.1000 43.4000 64.2000 ;
	    RECT 41.4000 63.8000 43.4000 64.1000 ;
	    RECT 40.7000 63.2000 42.5000 63.5000 ;
	    RECT 40.7000 63.1000 41.0000 63.2000 ;
	    RECT 40.6000 61.1000 41.0000 63.1000 ;
	    RECT 42.2000 63.1000 42.5000 63.2000 ;
	    RECT 42.2000 61.1000 42.6000 63.1000 ;
	    RECT 44.6000 61.1000 45.0000 65.8000 ;
	    RECT 45.4000 65.8000 45.8000 66.2000 ;
	    RECT 45.4000 65.1000 45.7000 65.8000 ;
	    RECT 46.2000 65.1000 46.6000 69.9000 ;
	    RECT 48.6000 68.9000 49.0000 69.9000 ;
	    RECT 47.0000 67.8000 47.4000 68.6000 ;
	    RECT 47.8000 67.8000 48.2000 68.6000 ;
	    RECT 48.7000 67.2000 49.0000 68.9000 ;
	    RECT 50.2000 67.5000 50.6000 69.9000 ;
	    RECT 52.4000 69.2000 52.8000 69.9000 ;
	    RECT 51.8000 68.9000 52.8000 69.2000 ;
	    RECT 54.6000 68.9000 55.0000 69.9000 ;
	    RECT 56.7000 69.2000 57.3000 69.9000 ;
	    RECT 56.6000 68.9000 57.3000 69.2000 ;
	    RECT 51.8000 68.5000 52.2000 68.9000 ;
	    RECT 54.6000 68.6000 54.9000 68.9000 ;
	    RECT 52.6000 67.8000 53.0000 68.6000 ;
	    RECT 53.5000 68.3000 54.9000 68.6000 ;
	    RECT 56.6000 68.5000 57.0000 68.9000 ;
	    RECT 53.5000 68.2000 53.9000 68.3000 ;
	    RECT 48.6000 66.8000 49.0000 67.2000 ;
	    RECT 50.6000 67.1000 51.4000 67.2000 ;
	    RECT 52.7000 67.1000 53.0000 67.8000 ;
	    RECT 57.5000 67.7000 57.9000 67.8000 ;
	    RECT 59.0000 67.7000 59.4000 69.9000 ;
	    RECT 62.2000 68.9000 62.6000 69.9000 ;
	    RECT 61.4000 67.8000 61.8000 68.6000 ;
	    RECT 57.5000 67.4000 59.4000 67.7000 ;
	    RECT 55.5000 67.1000 55.9000 67.2000 ;
	    RECT 50.6000 66.8000 56.1000 67.1000 ;
	    RECT 48.7000 65.1000 49.0000 66.8000 ;
	    RECT 52.1000 66.7000 52.5000 66.8000 ;
	    RECT 51.3000 66.2000 51.7000 66.3000 ;
	    RECT 55.8000 66.2000 56.1000 66.8000 ;
	    RECT 56.6000 66.4000 57.0000 66.5000 ;
	    RECT 49.4000 65.4000 49.8000 66.2000 ;
	    RECT 51.3000 65.9000 53.8000 66.2000 ;
	    RECT 53.4000 65.8000 53.8000 65.9000 ;
	    RECT 55.8000 65.8000 56.2000 66.2000 ;
	    RECT 56.6000 66.1000 58.5000 66.4000 ;
	    RECT 58.1000 66.0000 58.5000 66.1000 ;
	    RECT 50.2000 65.5000 53.0000 65.6000 ;
	    RECT 50.2000 65.4000 53.1000 65.5000 ;
	    RECT 50.2000 65.3000 55.1000 65.4000 ;
	    RECT 45.4000 64.8000 46.6000 65.1000 ;
	    RECT 46.2000 61.1000 46.6000 64.8000 ;
	    RECT 48.6000 64.7000 49.5000 65.1000 ;
	    RECT 49.1000 62.2000 49.5000 64.7000 ;
	    RECT 49.1000 61.8000 49.8000 62.2000 ;
	    RECT 49.1000 61.1000 49.5000 61.8000 ;
	    RECT 50.2000 61.1000 50.6000 65.3000 ;
	    RECT 52.7000 65.1000 55.1000 65.3000 ;
	    RECT 51.8000 64.5000 54.5000 64.8000 ;
	    RECT 51.8000 64.4000 52.2000 64.5000 ;
	    RECT 54.1000 64.4000 54.5000 64.5000 ;
	    RECT 54.8000 64.5000 55.1000 65.1000 ;
	    RECT 55.8000 65.2000 56.1000 65.8000 ;
	    RECT 57.3000 65.7000 57.7000 65.8000 ;
	    RECT 59.0000 65.7000 59.4000 67.4000 ;
	    RECT 62.3000 67.2000 62.6000 68.9000 ;
	    RECT 60.6000 67.1000 61.0000 67.2000 ;
	    RECT 62.2000 67.1000 62.6000 67.2000 ;
	    RECT 60.6000 66.8000 62.6000 67.1000 ;
	    RECT 65.6000 67.1000 66.0000 69.9000 ;
	    RECT 67.0000 68.0000 67.4000 69.9000 ;
	    RECT 68.6000 68.0000 69.0000 69.9000 ;
	    RECT 67.0000 67.9000 69.0000 68.0000 ;
	    RECT 69.4000 67.9000 69.8000 69.9000 ;
	    RECT 71.0000 68.9000 71.4000 69.9000 ;
	    RECT 67.1000 67.7000 68.9000 67.9000 ;
	    RECT 67.4000 67.2000 67.8000 67.4000 ;
	    RECT 69.4000 67.2000 69.7000 67.9000 ;
	    RECT 71.0000 67.2000 71.3000 68.9000 ;
	    RECT 71.8000 67.8000 72.2000 68.6000 ;
	    RECT 72.6000 67.5000 73.0000 69.9000 ;
	    RECT 74.8000 69.2000 75.2000 69.9000 ;
	    RECT 74.2000 68.9000 75.2000 69.2000 ;
	    RECT 77.0000 68.9000 77.4000 69.9000 ;
	    RECT 79.1000 69.2000 79.7000 69.9000 ;
	    RECT 79.0000 68.9000 79.7000 69.2000 ;
	    RECT 74.2000 68.5000 74.6000 68.9000 ;
	    RECT 77.0000 68.6000 77.3000 68.9000 ;
	    RECT 75.0000 68.2000 75.4000 68.6000 ;
	    RECT 75.9000 68.3000 77.3000 68.6000 ;
	    RECT 79.0000 68.5000 79.4000 68.9000 ;
	    RECT 75.9000 68.2000 76.3000 68.3000 ;
	    RECT 65.6000 66.9000 66.5000 67.1000 ;
	    RECT 65.7000 66.8000 66.5000 66.9000 ;
	    RECT 67.0000 66.9000 67.8000 67.2000 ;
	    RECT 67.0000 66.8000 67.4000 66.9000 ;
	    RECT 68.5000 66.8000 69.8000 67.2000 ;
	    RECT 71.0000 66.8000 71.4000 67.2000 ;
	    RECT 73.0000 67.1000 73.8000 67.2000 ;
	    RECT 75.1000 67.1000 75.4000 68.2000 ;
	    RECT 79.9000 67.7000 80.3000 67.8000 ;
	    RECT 81.4000 67.7000 81.8000 69.9000 ;
	    RECT 82.2000 67.9000 82.6000 69.9000 ;
	    RECT 83.0000 68.0000 83.4000 69.9000 ;
	    RECT 84.6000 68.0000 85.0000 69.9000 ;
	    RECT 85.5000 68.2000 85.9000 68.6000 ;
	    RECT 83.0000 67.9000 85.0000 68.0000 ;
	    RECT 79.9000 67.4000 81.8000 67.7000 ;
	    RECT 77.9000 67.1000 78.3000 67.2000 ;
	    RECT 73.0000 66.8000 78.5000 67.1000 ;
	    RECT 57.3000 65.4000 59.4000 65.7000 ;
	    RECT 55.8000 64.9000 57.0000 65.2000 ;
	    RECT 55.5000 64.5000 55.9000 64.6000 ;
	    RECT 54.8000 64.2000 55.9000 64.5000 ;
	    RECT 56.7000 64.4000 57.0000 64.9000 ;
	    RECT 56.7000 64.0000 57.4000 64.4000 ;
	    RECT 53.5000 63.7000 53.9000 63.8000 ;
	    RECT 54.9000 63.7000 55.3000 63.8000 ;
	    RECT 51.8000 63.1000 52.2000 63.5000 ;
	    RECT 53.5000 63.4000 55.3000 63.7000 ;
	    RECT 54.6000 63.1000 54.9000 63.4000 ;
	    RECT 56.6000 63.1000 57.0000 63.5000 ;
	    RECT 51.8000 62.8000 52.8000 63.1000 ;
	    RECT 52.4000 61.1000 52.8000 62.8000 ;
	    RECT 54.6000 61.1000 55.0000 63.1000 ;
	    RECT 56.7000 61.1000 57.3000 63.1000 ;
	    RECT 59.0000 61.1000 59.4000 65.4000 ;
	    RECT 62.3000 65.1000 62.6000 66.8000 ;
	    RECT 63.0000 65.4000 63.4000 66.2000 ;
	    RECT 64.6000 65.8000 65.4000 66.2000 ;
	    RECT 62.2000 64.7000 63.1000 65.1000 ;
	    RECT 63.8000 64.8000 64.2000 65.6000 ;
	    RECT 66.2000 65.2000 66.5000 66.8000 ;
	    RECT 67.8000 65.8000 68.2000 66.6000 ;
	    RECT 68.5000 66.1000 68.8000 66.8000 ;
	    RECT 70.2000 66.1000 70.6000 66.2000 ;
	    RECT 68.5000 65.8000 70.6000 66.1000 ;
	    RECT 66.2000 64.8000 66.6000 65.2000 ;
	    RECT 68.5000 65.1000 68.8000 65.8000 ;
	    RECT 70.2000 65.4000 70.6000 65.8000 ;
	    RECT 69.4000 65.1000 69.8000 65.2000 ;
	    RECT 71.0000 65.1000 71.3000 66.8000 ;
	    RECT 74.5000 66.7000 74.9000 66.8000 ;
	    RECT 73.7000 66.2000 74.1000 66.3000 ;
	    RECT 75.0000 66.2000 75.4000 66.3000 ;
	    RECT 78.2000 66.2000 78.5000 66.8000 ;
	    RECT 79.0000 66.4000 79.4000 66.5000 ;
	    RECT 73.7000 65.9000 76.2000 66.2000 ;
	    RECT 75.8000 65.8000 76.2000 65.9000 ;
	    RECT 78.2000 65.8000 78.6000 66.2000 ;
	    RECT 79.0000 66.1000 80.9000 66.4000 ;
	    RECT 80.5000 66.0000 80.9000 66.1000 ;
	    RECT 72.6000 65.5000 75.4000 65.6000 ;
	    RECT 72.6000 65.4000 75.5000 65.5000 ;
	    RECT 72.6000 65.3000 77.5000 65.4000 ;
	    RECT 68.3000 64.8000 68.8000 65.1000 ;
	    RECT 69.1000 64.8000 69.8000 65.1000 ;
	    RECT 62.7000 61.1000 63.1000 64.7000 ;
	    RECT 65.4000 63.8000 65.8000 64.6000 ;
	    RECT 66.2000 63.5000 66.5000 64.8000 ;
	    RECT 64.7000 63.2000 66.5000 63.5000 ;
	    RECT 64.7000 63.1000 65.0000 63.2000 ;
	    RECT 64.6000 61.1000 65.0000 63.1000 ;
	    RECT 66.2000 63.1000 66.5000 63.2000 ;
	    RECT 66.2000 61.1000 66.6000 63.1000 ;
	    RECT 68.3000 61.1000 68.7000 64.8000 ;
	    RECT 69.1000 64.2000 69.4000 64.8000 ;
	    RECT 69.0000 63.8000 69.4000 64.2000 ;
	    RECT 70.5000 64.7000 71.4000 65.1000 ;
	    RECT 70.5000 63.2000 70.9000 64.7000 ;
	    RECT 70.5000 62.8000 71.4000 63.2000 ;
	    RECT 70.5000 61.1000 70.9000 62.8000 ;
	    RECT 72.6000 61.1000 73.0000 65.3000 ;
	    RECT 75.1000 65.1000 77.5000 65.3000 ;
	    RECT 74.2000 64.5000 76.9000 64.8000 ;
	    RECT 74.2000 64.4000 74.6000 64.5000 ;
	    RECT 76.5000 64.4000 76.9000 64.5000 ;
	    RECT 77.2000 64.5000 77.5000 65.1000 ;
	    RECT 78.2000 65.2000 78.5000 65.8000 ;
	    RECT 79.7000 65.7000 80.1000 65.8000 ;
	    RECT 81.4000 65.7000 81.8000 67.4000 ;
	    RECT 82.3000 67.2000 82.6000 67.9000 ;
	    RECT 83.1000 67.7000 84.9000 67.9000 ;
	    RECT 85.4000 67.8000 85.8000 68.2000 ;
	    RECT 86.2000 67.9000 86.6000 69.9000 ;
	    RECT 84.2000 67.2000 84.6000 67.4000 ;
	    RECT 82.2000 66.8000 83.5000 67.2000 ;
	    RECT 84.2000 66.9000 85.0000 67.2000 ;
	    RECT 84.6000 66.8000 85.0000 66.9000 ;
	    RECT 79.7000 65.4000 81.8000 65.7000 ;
	    RECT 78.2000 64.9000 79.4000 65.2000 ;
	    RECT 77.9000 64.5000 78.3000 64.6000 ;
	    RECT 77.2000 64.2000 78.3000 64.5000 ;
	    RECT 79.1000 64.4000 79.4000 64.9000 ;
	    RECT 79.1000 64.0000 79.8000 64.4000 ;
	    RECT 75.9000 63.7000 76.3000 63.8000 ;
	    RECT 77.3000 63.7000 77.7000 63.8000 ;
	    RECT 74.2000 63.1000 74.6000 63.5000 ;
	    RECT 75.9000 63.4000 77.7000 63.7000 ;
	    RECT 77.0000 63.1000 77.3000 63.4000 ;
	    RECT 79.0000 63.1000 79.4000 63.5000 ;
	    RECT 74.2000 62.8000 75.2000 63.1000 ;
	    RECT 74.8000 61.1000 75.2000 62.8000 ;
	    RECT 77.0000 61.1000 77.4000 63.1000 ;
	    RECT 79.1000 61.1000 79.7000 63.1000 ;
	    RECT 81.4000 61.1000 81.8000 65.4000 ;
	    RECT 83.2000 65.2000 83.5000 66.8000 ;
	    RECT 83.8000 65.8000 84.2000 66.6000 ;
	    RECT 85.4000 66.1000 85.8000 66.2000 ;
	    RECT 86.3000 66.1000 86.6000 67.9000 ;
	    RECT 90.4000 67.2000 90.8000 69.9000 ;
	    RECT 92.6000 68.2000 93.0000 69.9000 ;
	    RECT 87.0000 66.4000 87.4000 67.2000 ;
	    RECT 90.2000 67.1000 90.8000 67.2000 ;
	    RECT 92.5000 67.9000 93.0000 68.2000 ;
	    RECT 92.5000 67.2000 92.8000 67.9000 ;
	    RECT 94.2000 67.6000 94.6000 69.9000 ;
	    RECT 95.8000 68.2000 96.2000 69.9000 ;
	    RECT 93.3000 67.3000 94.6000 67.6000 ;
	    RECT 95.7000 67.9000 96.2000 68.2000 ;
	    RECT 90.2000 66.8000 91.3000 67.1000 ;
	    RECT 87.8000 66.1000 88.2000 66.2000 ;
	    RECT 85.4000 65.8000 86.6000 66.1000 ;
	    RECT 87.4000 65.8000 88.2000 66.1000 ;
	    RECT 89.4000 65.8000 90.2000 66.2000 ;
	    RECT 82.2000 65.1000 82.6000 65.2000 ;
	    RECT 82.2000 64.8000 82.9000 65.1000 ;
	    RECT 83.2000 64.8000 84.2000 65.2000 ;
	    RECT 85.5000 65.1000 85.8000 65.8000 ;
	    RECT 87.4000 65.6000 87.8000 65.8000 ;
	    RECT 82.6000 64.2000 82.9000 64.8000 ;
	    RECT 82.6000 63.8000 83.0000 64.2000 ;
	    RECT 83.3000 61.1000 83.7000 64.8000 ;
	    RECT 85.4000 61.1000 85.8000 65.1000 ;
	    RECT 86.2000 64.8000 88.2000 65.1000 ;
	    RECT 88.6000 64.8000 89.0000 65.6000 ;
	    RECT 91.0000 65.2000 91.3000 66.8000 ;
	    RECT 92.5000 66.8000 93.0000 67.2000 ;
	    RECT 91.0000 64.8000 91.4000 65.2000 ;
	    RECT 92.5000 65.1000 92.8000 66.8000 ;
	    RECT 93.3000 66.5000 93.6000 67.3000 ;
	    RECT 95.7000 67.2000 96.0000 67.9000 ;
	    RECT 97.4000 67.6000 97.8000 69.9000 ;
	    RECT 99.0000 68.2000 99.4000 69.9000 ;
	    RECT 96.5000 67.3000 97.8000 67.6000 ;
	    RECT 98.9000 67.9000 99.4000 68.2000 ;
	    RECT 95.7000 66.8000 96.2000 67.2000 ;
	    RECT 93.1000 66.1000 93.6000 66.5000 ;
	    RECT 93.3000 65.1000 93.6000 66.1000 ;
	    RECT 94.1000 66.2000 94.5000 66.6000 ;
	    RECT 94.1000 65.8000 94.6000 66.2000 ;
	    RECT 95.7000 65.1000 96.0000 66.8000 ;
	    RECT 96.5000 66.5000 96.8000 67.3000 ;
	    RECT 98.9000 67.2000 99.2000 67.9000 ;
	    RECT 100.6000 67.6000 101.0000 69.9000 ;
	    RECT 102.2000 68.2000 102.6000 69.9000 ;
	    RECT 99.7000 67.3000 101.0000 67.6000 ;
	    RECT 102.1000 67.9000 102.6000 68.2000 ;
	    RECT 98.2000 67.1000 98.6000 67.2000 ;
	    RECT 98.9000 67.1000 99.4000 67.2000 ;
	    RECT 98.2000 66.8000 99.4000 67.1000 ;
	    RECT 96.3000 66.1000 96.8000 66.5000 ;
	    RECT 96.5000 65.1000 96.8000 66.1000 ;
	    RECT 97.3000 66.2000 97.7000 66.6000 ;
	    RECT 97.3000 65.8000 97.8000 66.2000 ;
	    RECT 98.9000 65.1000 99.2000 66.8000 ;
	    RECT 99.7000 66.5000 100.0000 67.3000 ;
	    RECT 102.1000 67.2000 102.4000 67.9000 ;
	    RECT 103.8000 67.6000 104.2000 69.9000 ;
	    RECT 105.4000 68.2000 105.8000 69.9000 ;
	    RECT 102.9000 67.3000 104.2000 67.6000 ;
	    RECT 105.3000 67.9000 105.8000 68.2000 ;
	    RECT 102.1000 67.1000 102.6000 67.2000 ;
	    RECT 101.4000 66.8000 102.6000 67.1000 ;
	    RECT 99.5000 66.1000 100.0000 66.5000 ;
	    RECT 99.7000 65.1000 100.0000 66.1000 ;
	    RECT 100.5000 66.2000 100.9000 66.6000 ;
	    RECT 101.4000 66.2000 101.7000 66.8000 ;
	    RECT 100.5000 65.8000 101.0000 66.2000 ;
	    RECT 101.4000 65.8000 101.8000 66.2000 ;
	    RECT 102.1000 65.1000 102.4000 66.8000 ;
	    RECT 102.9000 66.5000 103.2000 67.3000 ;
	    RECT 105.3000 67.2000 105.6000 67.9000 ;
	    RECT 107.0000 67.6000 107.4000 69.9000 ;
	    RECT 106.1000 67.3000 107.4000 67.6000 ;
	    RECT 109.4000 67.6000 109.8000 69.9000 ;
	    RECT 111.0000 68.2000 111.4000 69.9000 ;
	    RECT 111.0000 67.9000 111.5000 68.2000 ;
	    RECT 109.4000 67.3000 110.7000 67.6000 ;
	    RECT 105.3000 66.8000 105.8000 67.2000 ;
	    RECT 102.7000 66.1000 103.2000 66.5000 ;
	    RECT 102.9000 65.1000 103.2000 66.1000 ;
	    RECT 103.7000 66.2000 104.1000 66.6000 ;
	    RECT 103.7000 66.1000 104.2000 66.2000 ;
	    RECT 104.6000 66.1000 105.0000 66.2000 ;
	    RECT 103.7000 65.8000 105.0000 66.1000 ;
	    RECT 105.3000 65.1000 105.6000 66.8000 ;
	    RECT 106.1000 66.5000 106.4000 67.3000 ;
	    RECT 105.9000 66.1000 106.4000 66.5000 ;
	    RECT 106.1000 65.1000 106.4000 66.1000 ;
	    RECT 106.9000 66.2000 107.3000 66.6000 ;
	    RECT 109.5000 66.2000 109.9000 66.6000 ;
	    RECT 106.9000 65.8000 107.4000 66.2000 ;
	    RECT 107.8000 66.1000 108.2000 66.2000 ;
	    RECT 109.4000 66.1000 109.9000 66.2000 ;
	    RECT 107.8000 65.8000 109.9000 66.1000 ;
	    RECT 110.4000 66.5000 110.7000 67.3000 ;
	    RECT 111.2000 67.2000 111.5000 67.9000 ;
	    RECT 112.6000 67.6000 113.0000 69.9000 ;
	    RECT 114.2000 68.2000 114.6000 69.9000 ;
	    RECT 114.2000 67.9000 114.7000 68.2000 ;
	    RECT 112.6000 67.3000 113.9000 67.6000 ;
	    RECT 111.0000 67.1000 111.5000 67.2000 ;
	    RECT 111.0000 66.8000 112.1000 67.1000 ;
	    RECT 110.4000 66.1000 110.9000 66.5000 ;
	    RECT 110.4000 65.1000 110.7000 66.1000 ;
	    RECT 111.2000 65.1000 111.5000 66.8000 ;
	    RECT 111.8000 66.2000 112.1000 66.8000 ;
	    RECT 112.7000 66.2000 113.1000 66.6000 ;
	    RECT 111.8000 65.8000 112.2000 66.2000 ;
	    RECT 112.6000 65.8000 113.1000 66.2000 ;
	    RECT 113.6000 66.5000 113.9000 67.3000 ;
	    RECT 114.4000 67.2000 114.7000 67.9000 ;
	    RECT 114.2000 66.8000 114.7000 67.2000 ;
	    RECT 117.6000 67.1000 118.0000 69.9000 ;
	    RECT 119.1000 68.2000 119.5000 68.6000 ;
	    RECT 119.0000 67.8000 119.4000 68.2000 ;
	    RECT 119.8000 67.9000 120.2000 69.9000 ;
	    RECT 122.2000 67.9000 122.6000 69.9000 ;
	    RECT 123.0000 68.0000 123.4000 69.9000 ;
	    RECT 124.6000 68.0000 125.0000 69.9000 ;
	    RECT 123.0000 67.9000 125.0000 68.0000 ;
	    RECT 125.4000 67.9000 125.8000 69.9000 ;
	    RECT 126.2000 68.0000 126.6000 69.9000 ;
	    RECT 127.8000 68.0000 128.2000 69.9000 ;
	    RECT 126.2000 67.9000 128.2000 68.0000 ;
	    RECT 117.6000 66.9000 118.5000 67.1000 ;
	    RECT 117.7000 66.8000 118.5000 66.9000 ;
	    RECT 113.6000 66.1000 114.1000 66.5000 ;
	    RECT 113.6000 65.1000 113.9000 66.1000 ;
	    RECT 114.4000 65.1000 114.7000 66.8000 ;
	    RECT 118.2000 66.2000 118.5000 66.8000 ;
	    RECT 115.0000 66.1000 115.4000 66.2000 ;
	    RECT 115.0000 65.8000 116.2000 66.1000 ;
	    RECT 116.6000 65.8000 117.4000 66.2000 ;
	    RECT 118.2000 65.8000 118.6000 66.2000 ;
	    RECT 119.0000 66.1000 119.4000 66.2000 ;
	    RECT 119.9000 66.1000 120.2000 67.9000 ;
	    RECT 122.3000 67.2000 122.6000 67.9000 ;
	    RECT 123.1000 67.7000 124.9000 67.9000 ;
	    RECT 124.2000 67.2000 124.6000 67.4000 ;
	    RECT 125.5000 67.2000 125.8000 67.9000 ;
	    RECT 126.3000 67.7000 128.1000 67.9000 ;
	    RECT 128.6000 67.6000 129.0000 69.9000 ;
	    RECT 130.2000 68.2000 130.6000 69.9000 ;
	    RECT 130.2000 67.9000 130.7000 68.2000 ;
	    RECT 127.4000 67.2000 127.8000 67.4000 ;
	    RECT 128.6000 67.3000 129.9000 67.6000 ;
	    RECT 120.6000 66.4000 121.0000 67.2000 ;
	    RECT 122.2000 66.8000 123.5000 67.2000 ;
	    RECT 124.2000 66.9000 125.0000 67.2000 ;
	    RECT 124.6000 66.8000 125.0000 66.9000 ;
	    RECT 125.4000 66.8000 126.7000 67.2000 ;
	    RECT 127.4000 66.9000 128.2000 67.2000 ;
	    RECT 127.8000 66.8000 128.2000 66.9000 ;
	    RECT 121.4000 66.1000 121.8000 66.2000 ;
	    RECT 119.0000 65.8000 120.2000 66.1000 ;
	    RECT 121.0000 65.8000 121.8000 66.1000 ;
	    RECT 86.2000 61.1000 86.6000 64.8000 ;
	    RECT 87.8000 61.1000 88.2000 64.8000 ;
	    RECT 90.2000 63.8000 90.6000 64.6000 ;
	    RECT 91.0000 63.5000 91.3000 64.8000 ;
	    RECT 92.5000 64.6000 93.0000 65.1000 ;
	    RECT 93.3000 64.8000 94.6000 65.1000 ;
	    RECT 89.5000 63.2000 91.3000 63.5000 ;
	    RECT 89.5000 63.1000 89.8000 63.2000 ;
	    RECT 89.4000 61.1000 89.8000 63.1000 ;
	    RECT 91.0000 63.1000 91.3000 63.2000 ;
	    RECT 91.0000 61.1000 91.4000 63.1000 ;
	    RECT 92.6000 61.1000 93.0000 64.6000 ;
	    RECT 94.2000 61.1000 94.6000 64.8000 ;
	    RECT 95.7000 64.6000 96.2000 65.1000 ;
	    RECT 96.5000 64.8000 97.8000 65.1000 ;
	    RECT 95.8000 61.1000 96.2000 64.6000 ;
	    RECT 97.4000 61.1000 97.8000 64.8000 ;
	    RECT 98.9000 64.6000 99.4000 65.1000 ;
	    RECT 99.7000 64.8000 101.0000 65.1000 ;
	    RECT 99.0000 61.1000 99.4000 64.6000 ;
	    RECT 100.6000 61.1000 101.0000 64.8000 ;
	    RECT 102.1000 64.6000 102.6000 65.1000 ;
	    RECT 102.9000 64.8000 104.2000 65.1000 ;
	    RECT 102.2000 61.1000 102.6000 64.6000 ;
	    RECT 103.8000 61.1000 104.2000 64.8000 ;
	    RECT 105.3000 64.6000 105.8000 65.1000 ;
	    RECT 106.1000 64.8000 107.4000 65.1000 ;
	    RECT 105.4000 61.1000 105.8000 64.6000 ;
	    RECT 107.0000 61.1000 107.4000 64.8000 ;
	    RECT 109.4000 64.8000 110.7000 65.1000 ;
	    RECT 109.4000 61.1000 109.8000 64.8000 ;
	    RECT 111.0000 64.6000 111.5000 65.1000 ;
	    RECT 112.6000 64.8000 113.9000 65.1000 ;
	    RECT 111.0000 61.1000 111.4000 64.6000 ;
	    RECT 112.6000 61.1000 113.0000 64.8000 ;
	    RECT 114.2000 64.6000 114.7000 65.1000 ;
	    RECT 115.8000 64.8000 116.2000 65.8000 ;
	    RECT 118.2000 65.2000 118.5000 65.8000 ;
	    RECT 118.2000 64.8000 118.6000 65.2000 ;
	    RECT 119.1000 65.1000 119.4000 65.8000 ;
	    RECT 121.0000 65.6000 121.4000 65.8000 ;
	    RECT 122.2000 65.1000 122.6000 65.2000 ;
	    RECT 123.2000 65.1000 123.5000 66.8000 ;
	    RECT 123.8000 65.8000 124.2000 66.6000 ;
	    RECT 125.4000 65.1000 125.8000 65.2000 ;
	    RECT 126.4000 65.1000 126.7000 66.8000 ;
	    RECT 127.0000 65.8000 127.4000 66.6000 ;
	    RECT 128.7000 66.2000 129.1000 66.6000 ;
	    RECT 127.8000 66.1000 128.2000 66.2000 ;
	    RECT 128.6000 66.1000 129.1000 66.2000 ;
	    RECT 127.8000 65.8000 129.1000 66.1000 ;
	    RECT 129.6000 66.5000 129.9000 67.3000 ;
	    RECT 130.4000 67.2000 130.7000 67.9000 ;
	    RECT 131.8000 67.6000 132.2000 69.9000 ;
	    RECT 133.4000 68.2000 133.8000 69.9000 ;
	    RECT 133.4000 67.9000 133.9000 68.2000 ;
	    RECT 131.8000 67.3000 133.1000 67.6000 ;
	    RECT 130.2000 66.8000 130.7000 67.2000 ;
	    RECT 129.6000 66.1000 130.1000 66.5000 ;
	    RECT 129.6000 65.1000 129.9000 66.1000 ;
	    RECT 130.4000 65.1000 130.7000 66.8000 ;
	    RECT 131.9000 66.2000 132.3000 66.6000 ;
	    RECT 131.8000 65.8000 132.3000 66.2000 ;
	    RECT 132.8000 66.5000 133.1000 67.3000 ;
	    RECT 133.6000 67.2000 133.9000 67.9000 ;
	    RECT 135.8000 67.6000 136.2000 69.9000 ;
	    RECT 137.4000 67.6000 137.8000 69.9000 ;
	    RECT 139.0000 67.9000 139.4000 69.9000 ;
	    RECT 139.8000 68.0000 140.2000 69.9000 ;
	    RECT 141.4000 68.0000 141.8000 69.9000 ;
	    RECT 139.8000 67.9000 141.8000 68.0000 ;
	    RECT 143.8000 67.9000 144.2000 69.9000 ;
	    RECT 144.5000 68.2000 144.9000 68.6000 ;
	    RECT 133.4000 67.1000 133.9000 67.2000 ;
	    RECT 134.2000 67.1000 134.6000 67.2000 ;
	    RECT 133.4000 66.8000 134.6000 67.1000 ;
	    RECT 135.0000 66.8000 135.4000 67.6000 ;
	    RECT 135.8000 67.2000 137.8000 67.6000 ;
	    RECT 139.1000 67.2000 139.4000 67.9000 ;
	    RECT 139.9000 67.7000 141.7000 67.9000 ;
	    RECT 141.0000 67.2000 141.4000 67.4000 ;
	    RECT 132.8000 66.1000 133.3000 66.5000 ;
	    RECT 132.8000 65.1000 133.1000 66.1000 ;
	    RECT 133.6000 65.1000 133.9000 66.8000 ;
	    RECT 137.4000 65.8000 137.8000 67.2000 ;
	    RECT 139.0000 66.8000 140.3000 67.2000 ;
	    RECT 141.0000 66.9000 141.8000 67.2000 ;
	    RECT 141.4000 66.8000 141.8000 66.9000 ;
	    RECT 142.2000 67.1000 142.6000 67.2000 ;
	    RECT 143.0000 67.1000 143.4000 67.2000 ;
	    RECT 142.2000 66.8000 143.4000 67.1000 ;
	    RECT 114.2000 61.1000 114.6000 64.6000 ;
	    RECT 117.4000 63.8000 117.8000 64.6000 ;
	    RECT 118.2000 63.5000 118.5000 64.8000 ;
	    RECT 116.7000 63.2000 118.5000 63.5000 ;
	    RECT 116.7000 63.1000 117.0000 63.2000 ;
	    RECT 116.6000 61.1000 117.0000 63.1000 ;
	    RECT 118.2000 63.1000 118.5000 63.2000 ;
	    RECT 118.2000 61.1000 118.6000 63.1000 ;
	    RECT 119.0000 61.1000 119.4000 65.1000 ;
	    RECT 119.8000 64.8000 121.8000 65.1000 ;
	    RECT 122.2000 64.8000 122.9000 65.1000 ;
	    RECT 123.2000 64.8000 123.7000 65.1000 ;
	    RECT 125.4000 64.8000 126.1000 65.1000 ;
	    RECT 126.4000 64.8000 126.9000 65.1000 ;
	    RECT 119.8000 61.1000 120.2000 64.8000 ;
	    RECT 121.4000 61.1000 121.8000 64.8000 ;
	    RECT 122.6000 64.2000 122.9000 64.8000 ;
	    RECT 122.2000 63.8000 123.0000 64.2000 ;
	    RECT 123.3000 62.2000 123.7000 64.8000 ;
	    RECT 125.8000 64.2000 126.1000 64.8000 ;
	    RECT 125.8000 63.8000 126.2000 64.2000 ;
	    RECT 123.3000 61.8000 124.2000 62.2000 ;
	    RECT 123.3000 61.1000 123.7000 61.8000 ;
	    RECT 126.5000 61.1000 126.9000 64.8000 ;
	    RECT 128.6000 64.8000 129.9000 65.1000 ;
	    RECT 128.6000 61.1000 129.0000 64.8000 ;
	    RECT 130.2000 64.6000 130.7000 65.1000 ;
	    RECT 131.8000 64.8000 133.1000 65.1000 ;
	    RECT 130.2000 61.1000 130.6000 64.6000 ;
	    RECT 131.8000 61.1000 132.2000 64.8000 ;
	    RECT 133.4000 64.6000 133.9000 65.1000 ;
	    RECT 135.8000 65.4000 137.8000 65.8000 ;
	    RECT 133.4000 61.1000 133.8000 64.6000 ;
	    RECT 135.8000 61.1000 136.2000 65.4000 ;
	    RECT 137.4000 61.1000 137.8000 65.4000 ;
	    RECT 139.0000 65.1000 139.4000 65.2000 ;
	    RECT 140.0000 65.1000 140.3000 66.8000 ;
	    RECT 140.6000 65.8000 141.0000 66.6000 ;
	    RECT 143.0000 66.4000 143.4000 66.8000 ;
	    RECT 142.2000 66.1000 142.6000 66.2000 ;
	    RECT 143.8000 66.1000 144.1000 67.9000 ;
	    RECT 144.6000 67.8000 145.0000 68.2000 ;
	    RECT 145.4000 68.0000 145.8000 69.9000 ;
	    RECT 147.0000 68.0000 147.4000 69.9000 ;
	    RECT 145.4000 67.9000 147.4000 68.0000 ;
	    RECT 147.8000 67.9000 148.2000 69.9000 ;
	    RECT 150.2000 67.9000 150.6000 69.9000 ;
	    RECT 150.9000 68.2000 151.3000 68.6000 ;
	    RECT 145.5000 67.7000 147.3000 67.9000 ;
	    RECT 145.8000 67.2000 146.2000 67.4000 ;
	    RECT 147.8000 67.2000 148.1000 67.9000 ;
	    RECT 145.4000 66.9000 146.2000 67.2000 ;
	    RECT 146.9000 67.1000 148.2000 67.2000 ;
	    RECT 149.4000 67.1000 149.8000 67.2000 ;
	    RECT 145.4000 66.8000 145.8000 66.9000 ;
	    RECT 146.9000 66.8000 149.8000 67.1000 ;
	    RECT 144.6000 66.1000 145.0000 66.2000 ;
	    RECT 142.2000 65.8000 143.0000 66.1000 ;
	    RECT 143.8000 65.8000 145.0000 66.1000 ;
	    RECT 146.2000 65.8000 146.6000 66.6000 ;
	    RECT 142.6000 65.6000 143.0000 65.8000 ;
	    RECT 144.6000 65.1000 144.9000 65.8000 ;
	    RECT 146.9000 65.1000 147.2000 66.8000 ;
	    RECT 149.4000 66.4000 149.8000 66.8000 ;
	    RECT 148.6000 66.1000 149.0000 66.2000 ;
	    RECT 150.2000 66.1000 150.5000 67.9000 ;
	    RECT 151.0000 67.8000 151.4000 68.2000 ;
	    RECT 151.8000 67.7000 152.2000 69.9000 ;
	    RECT 153.9000 69.2000 154.5000 69.9000 ;
	    RECT 153.9000 68.9000 154.6000 69.2000 ;
	    RECT 156.2000 68.9000 156.6000 69.9000 ;
	    RECT 158.4000 69.2000 158.8000 69.9000 ;
	    RECT 158.4000 68.9000 159.4000 69.2000 ;
	    RECT 154.2000 68.5000 154.6000 68.9000 ;
	    RECT 156.3000 68.6000 156.6000 68.9000 ;
	    RECT 156.3000 68.3000 157.7000 68.6000 ;
	    RECT 157.3000 68.2000 157.7000 68.3000 ;
	    RECT 158.2000 68.2000 158.6000 68.6000 ;
	    RECT 159.0000 68.5000 159.4000 68.9000 ;
	    RECT 153.3000 67.7000 153.7000 67.8000 ;
	    RECT 151.8000 67.4000 153.7000 67.7000 ;
	    RECT 151.0000 66.8000 151.4000 67.2000 ;
	    RECT 151.0000 66.2000 151.3000 66.8000 ;
	    RECT 151.0000 66.1000 151.4000 66.2000 ;
	    RECT 148.6000 65.8000 149.4000 66.1000 ;
	    RECT 150.2000 65.8000 151.4000 66.1000 ;
	    RECT 149.0000 65.6000 149.4000 65.8000 ;
	    RECT 147.8000 65.1000 148.2000 65.2000 ;
	    RECT 151.0000 65.1000 151.3000 65.8000 ;
	    RECT 151.8000 65.7000 152.2000 67.4000 ;
	    RECT 155.3000 67.1000 155.7000 67.2000 ;
	    RECT 158.2000 67.1000 158.5000 68.2000 ;
	    RECT 160.6000 67.5000 161.0000 69.9000 ;
	    RECT 164.3000 68.2000 164.7000 69.9000 ;
	    RECT 163.8000 67.9000 164.7000 68.2000 ;
	    RECT 159.8000 67.1000 160.6000 67.2000 ;
	    RECT 161.4000 67.1000 161.8000 67.2000 ;
	    RECT 155.1000 66.8000 161.8000 67.1000 ;
	    RECT 162.2000 67.1000 162.6000 67.2000 ;
	    RECT 163.0000 67.1000 163.4000 67.6000 ;
	    RECT 162.2000 66.8000 163.4000 67.1000 ;
	    RECT 154.2000 66.4000 154.6000 66.5000 ;
	    RECT 152.7000 66.1000 154.6000 66.4000 ;
	    RECT 155.1000 66.2000 155.4000 66.8000 ;
	    RECT 158.7000 66.7000 159.1000 66.8000 ;
	    RECT 159.5000 66.2000 159.9000 66.3000 ;
	    RECT 152.7000 66.0000 153.1000 66.1000 ;
	    RECT 155.0000 65.8000 155.4000 66.2000 ;
	    RECT 155.8000 66.1000 156.2000 66.2000 ;
	    RECT 157.4000 66.1000 159.9000 66.2000 ;
	    RECT 155.8000 65.9000 159.9000 66.1000 ;
	    RECT 155.8000 65.8000 157.8000 65.9000 ;
	    RECT 153.5000 65.7000 153.9000 65.8000 ;
	    RECT 151.8000 65.4000 153.9000 65.7000 ;
	    RECT 139.0000 64.8000 139.7000 65.1000 ;
	    RECT 140.0000 64.8000 140.5000 65.1000 ;
	    RECT 139.4000 64.2000 139.7000 64.8000 ;
	    RECT 139.4000 63.8000 139.8000 64.2000 ;
	    RECT 140.1000 61.1000 140.5000 64.8000 ;
	    RECT 142.2000 64.8000 144.2000 65.1000 ;
	    RECT 142.2000 61.1000 142.6000 64.8000 ;
	    RECT 143.8000 61.1000 144.2000 64.8000 ;
	    RECT 144.6000 61.1000 145.0000 65.1000 ;
	    RECT 146.7000 64.8000 147.2000 65.1000 ;
	    RECT 147.5000 64.8000 148.2000 65.1000 ;
	    RECT 148.6000 64.8000 150.6000 65.1000 ;
	    RECT 146.7000 61.1000 147.1000 64.8000 ;
	    RECT 147.5000 64.2000 147.8000 64.8000 ;
	    RECT 147.4000 63.8000 148.2000 64.2000 ;
	    RECT 148.6000 61.1000 149.0000 64.8000 ;
	    RECT 150.2000 61.1000 150.6000 64.8000 ;
	    RECT 151.0000 61.1000 151.4000 65.1000 ;
	    RECT 151.8000 61.1000 152.2000 65.4000 ;
	    RECT 155.1000 65.2000 155.4000 65.8000 ;
	    RECT 158.2000 65.5000 161.0000 65.6000 ;
	    RECT 158.1000 65.4000 161.0000 65.5000 ;
	    RECT 154.2000 64.9000 155.4000 65.2000 ;
	    RECT 156.1000 65.3000 161.0000 65.4000 ;
	    RECT 156.1000 65.1000 158.5000 65.3000 ;
	    RECT 154.2000 64.4000 154.5000 64.9000 ;
	    RECT 153.8000 64.0000 154.5000 64.4000 ;
	    RECT 155.3000 64.5000 155.7000 64.6000 ;
	    RECT 156.1000 64.5000 156.4000 65.1000 ;
	    RECT 155.3000 64.2000 156.4000 64.5000 ;
	    RECT 156.7000 64.5000 159.4000 64.8000 ;
	    RECT 156.7000 64.4000 157.1000 64.5000 ;
	    RECT 159.0000 64.4000 159.4000 64.5000 ;
	    RECT 155.9000 63.7000 156.3000 63.8000 ;
	    RECT 157.3000 63.7000 157.7000 63.8000 ;
	    RECT 154.2000 63.1000 154.6000 63.5000 ;
	    RECT 155.9000 63.4000 157.7000 63.7000 ;
	    RECT 156.3000 63.1000 156.6000 63.4000 ;
	    RECT 159.0000 63.1000 159.4000 63.5000 ;
	    RECT 153.9000 61.1000 154.5000 63.1000 ;
	    RECT 156.2000 61.1000 156.6000 63.1000 ;
	    RECT 158.4000 62.8000 159.4000 63.1000 ;
	    RECT 158.4000 61.1000 158.8000 62.8000 ;
	    RECT 160.6000 61.1000 161.0000 65.3000 ;
	    RECT 163.8000 61.1000 164.2000 67.9000 ;
	    RECT 164.6000 65.1000 165.0000 65.2000 ;
	    RECT 165.4000 65.1000 165.8000 69.9000 ;
	    RECT 166.2000 67.8000 166.6000 68.6000 ;
	    RECT 167.8000 68.2000 168.2000 69.9000 ;
	    RECT 167.7000 67.9000 168.2000 68.2000 ;
	    RECT 164.6000 64.8000 165.8000 65.1000 ;
	    RECT 164.6000 64.4000 165.0000 64.8000 ;
	    RECT 165.4000 61.1000 165.8000 64.8000 ;
	    RECT 167.7000 67.2000 168.0000 67.9000 ;
	    RECT 169.4000 67.6000 169.8000 69.9000 ;
	    RECT 168.5000 67.3000 169.8000 67.6000 ;
	    RECT 170.2000 67.6000 170.6000 69.9000 ;
	    RECT 171.8000 68.2000 172.2000 69.9000 ;
	    RECT 171.8000 67.9000 172.3000 68.2000 ;
	    RECT 170.2000 67.3000 171.5000 67.6000 ;
	    RECT 167.7000 66.8000 168.2000 67.2000 ;
	    RECT 167.7000 65.1000 168.0000 66.8000 ;
	    RECT 168.5000 66.5000 168.8000 67.3000 ;
	    RECT 168.3000 66.1000 168.8000 66.5000 ;
	    RECT 168.5000 65.1000 168.8000 66.1000 ;
	    RECT 171.2000 66.5000 171.5000 67.3000 ;
	    RECT 172.0000 67.2000 172.3000 67.9000 ;
	    RECT 171.8000 66.8000 172.3000 67.2000 ;
	    RECT 171.2000 66.1000 171.7000 66.5000 ;
	    RECT 171.2000 65.1000 171.5000 66.1000 ;
	    RECT 172.0000 65.1000 172.3000 66.8000 ;
	    RECT 172.6000 66.1000 173.0000 66.2000 ;
	    RECT 173.4000 66.1000 173.8000 69.9000 ;
	    RECT 174.2000 67.8000 174.6000 68.6000 ;
	    RECT 175.0000 67.8000 175.4000 68.6000 ;
	    RECT 175.0000 67.1000 175.4000 67.2000 ;
	    RECT 175.8000 67.1000 176.2000 69.9000 ;
	    RECT 176.9000 68.2000 177.3000 69.9000 ;
	    RECT 179.0000 68.5000 179.4000 69.5000 ;
	    RECT 175.0000 66.8000 176.2000 67.1000 ;
	    RECT 176.6000 67.8000 177.8000 68.2000 ;
	    RECT 176.6000 67.2000 176.9000 67.8000 ;
	    RECT 176.6000 66.8000 177.0000 67.2000 ;
	    RECT 172.6000 65.8000 173.8000 66.1000 ;
	    RECT 167.7000 64.6000 168.2000 65.1000 ;
	    RECT 168.5000 64.8000 169.8000 65.1000 ;
	    RECT 167.8000 61.1000 168.2000 64.6000 ;
	    RECT 169.4000 61.1000 169.8000 64.8000 ;
	    RECT 170.2000 64.8000 171.5000 65.1000 ;
	    RECT 170.2000 61.1000 170.6000 64.8000 ;
	    RECT 171.8000 64.6000 172.3000 65.1000 ;
	    RECT 171.8000 61.1000 172.2000 64.6000 ;
	    RECT 173.4000 61.1000 173.8000 65.8000 ;
	    RECT 175.8000 61.1000 176.2000 66.8000 ;
	    RECT 176.6000 64.4000 177.0000 65.2000 ;
	    RECT 177.4000 61.1000 177.8000 67.8000 ;
	    RECT 178.2000 66.8000 178.6000 67.6000 ;
	    RECT 179.0000 67.4000 179.3000 68.5000 ;
	    RECT 181.1000 68.0000 181.5000 69.5000 ;
	    RECT 184.6000 68.9000 185.0000 69.9000 ;
	    RECT 187.0000 68.9000 187.4000 69.9000 ;
	    RECT 181.1000 67.7000 181.9000 68.0000 ;
	    RECT 183.8000 67.8000 184.2000 68.6000 ;
	    RECT 181.5000 67.5000 181.9000 67.7000 ;
	    RECT 179.0000 67.1000 181.1000 67.4000 ;
	    RECT 180.6000 66.9000 181.1000 67.1000 ;
	    RECT 181.6000 67.2000 181.9000 67.5000 ;
	    RECT 184.7000 67.2000 185.0000 68.9000 ;
	    RECT 186.2000 67.8000 186.6000 68.6000 ;
	    RECT 187.1000 67.8000 187.4000 68.9000 ;
	    RECT 188.6000 67.9000 189.0000 69.9000 ;
	    RECT 191.3000 68.0000 191.7000 69.5000 ;
	    RECT 193.4000 68.5000 193.8000 69.5000 ;
	    RECT 187.1000 67.5000 188.3000 67.8000 ;
	    RECT 178.2000 66.1000 178.6000 66.2000 ;
	    RECT 179.0000 66.1000 179.4000 66.6000 ;
	    RECT 178.2000 65.8000 179.4000 66.1000 ;
	    RECT 179.8000 65.8000 180.2000 66.6000 ;
	    RECT 180.6000 66.5000 181.3000 66.9000 ;
	    RECT 181.6000 66.8000 182.6000 67.2000 ;
	    RECT 184.6000 67.1000 185.0000 67.2000 ;
	    RECT 185.4000 67.1000 185.8000 67.2000 ;
	    RECT 184.6000 66.8000 185.8000 67.1000 ;
	    RECT 187.0000 66.8000 187.5000 67.2000 ;
	    RECT 180.6000 65.5000 180.9000 66.5000 ;
	    RECT 179.0000 65.2000 180.9000 65.5000 ;
	    RECT 179.0000 63.5000 179.3000 65.2000 ;
	    RECT 181.6000 64.9000 181.9000 66.8000 ;
	    RECT 182.2000 66.1000 182.6000 66.2000 ;
	    RECT 184.7000 66.1000 185.0000 66.8000 ;
	    RECT 187.2000 66.4000 187.6000 66.8000 ;
	    RECT 182.2000 65.8000 185.0000 66.1000 ;
	    RECT 182.2000 65.4000 182.6000 65.8000 ;
	    RECT 184.7000 65.1000 185.0000 65.8000 ;
	    RECT 185.4000 65.4000 185.8000 66.2000 ;
	    RECT 188.0000 66.0000 188.3000 67.5000 ;
	    RECT 188.7000 66.2000 189.0000 67.9000 ;
	    RECT 190.9000 67.7000 191.7000 68.0000 ;
	    RECT 190.9000 67.5000 191.3000 67.7000 ;
	    RECT 190.9000 67.2000 191.2000 67.5000 ;
	    RECT 193.5000 67.4000 193.8000 68.5000 ;
	    RECT 194.2000 67.9000 194.6000 69.9000 ;
	    RECT 196.4000 69.2000 197.2000 69.9000 ;
	    RECT 195.8000 68.8000 197.2000 69.2000 ;
	    RECT 196.4000 68.1000 197.2000 68.8000 ;
	    RECT 194.2000 67.6000 195.4000 67.9000 ;
	    RECT 195.0000 67.5000 195.4000 67.6000 ;
	    RECT 190.2000 66.8000 191.2000 67.2000 ;
	    RECT 191.7000 67.1000 193.8000 67.4000 ;
	    RECT 195.7000 67.4000 196.1000 67.8000 ;
	    RECT 195.7000 67.2000 196.0000 67.4000 ;
	    RECT 191.7000 66.9000 192.2000 67.1000 ;
	    RECT 187.9000 65.7000 188.3000 66.0000 ;
	    RECT 188.6000 66.1000 189.0000 66.2000 ;
	    RECT 189.4000 66.1000 189.8000 66.2000 ;
	    RECT 188.6000 65.8000 189.8000 66.1000 ;
	    RECT 186.2000 65.6000 188.3000 65.7000 ;
	    RECT 186.2000 65.4000 188.2000 65.6000 ;
	    RECT 181.1000 64.6000 181.9000 64.9000 ;
	    RECT 184.6000 64.7000 185.5000 65.1000 ;
	    RECT 179.0000 61.5000 179.4000 63.5000 ;
	    RECT 181.1000 62.2000 181.5000 64.6000 ;
	    RECT 180.6000 61.8000 181.5000 62.2000 ;
	    RECT 181.1000 61.1000 181.5000 61.8000 ;
	    RECT 185.1000 61.1000 185.5000 64.7000 ;
	    RECT 186.2000 61.1000 186.6000 65.4000 ;
	    RECT 188.7000 65.1000 189.0000 65.8000 ;
	    RECT 190.2000 65.4000 190.6000 66.2000 ;
	    RECT 188.3000 64.8000 189.0000 65.1000 ;
	    RECT 190.9000 64.9000 191.2000 66.8000 ;
	    RECT 191.5000 66.5000 192.2000 66.9000 ;
	    RECT 194.2000 66.8000 195.0000 67.2000 ;
	    RECT 195.6000 66.8000 196.0000 67.2000 ;
	    RECT 191.9000 65.5000 192.2000 66.5000 ;
	    RECT 192.6000 65.8000 193.0000 66.6000 ;
	    RECT 193.4000 65.8000 193.8000 66.6000 ;
	    RECT 196.4000 66.4000 196.7000 68.1000 ;
	    RECT 199.0000 67.9000 199.4000 69.9000 ;
	    RECT 197.0000 67.7000 197.8000 67.8000 ;
	    RECT 197.0000 67.4000 198.0000 67.7000 ;
	    RECT 198.3000 67.6000 199.4000 67.9000 ;
	    RECT 198.3000 67.5000 198.7000 67.6000 ;
	    RECT 197.7000 67.2000 198.0000 67.4000 ;
	    RECT 197.0000 66.7000 197.4000 67.1000 ;
	    RECT 197.7000 66.9000 199.4000 67.2000 ;
	    RECT 198.6000 66.8000 199.4000 66.9000 ;
	    RECT 196.2000 66.2000 196.7000 66.4000 ;
	    RECT 195.8000 66.1000 196.7000 66.2000 ;
	    RECT 197.1000 66.4000 197.4000 66.7000 ;
	    RECT 197.1000 66.1000 198.4000 66.4000 ;
	    RECT 195.8000 65.8000 196.5000 66.1000 ;
	    RECT 198.0000 66.0000 198.4000 66.1000 ;
	    RECT 199.8000 66.2000 200.2000 69.9000 ;
	    RECT 201.4000 67.6000 201.8000 69.9000 ;
	    RECT 203.5000 69.2000 203.9000 69.9000 ;
	    RECT 203.5000 68.8000 204.2000 69.2000 ;
	    RECT 203.5000 68.2000 203.9000 68.8000 ;
	    RECT 203.0000 67.9000 203.9000 68.2000 ;
	    RECT 200.7000 67.3000 201.8000 67.6000 ;
	    RECT 191.9000 65.2000 193.8000 65.5000 ;
	    RECT 188.3000 61.1000 188.7000 64.8000 ;
	    RECT 190.9000 64.6000 191.7000 64.9000 ;
	    RECT 191.3000 62.2000 191.7000 64.6000 ;
	    RECT 193.5000 63.5000 193.8000 65.2000 ;
	    RECT 196.2000 65.1000 196.5000 65.8000 ;
	    RECT 196.9000 65.7000 197.3000 65.8000 ;
	    RECT 196.9000 65.4000 198.6000 65.7000 ;
	    RECT 198.3000 65.1000 198.6000 65.4000 ;
	    RECT 199.8000 65.1000 200.1000 66.2000 ;
	    RECT 200.7000 65.8000 201.0000 67.3000 ;
	    RECT 202.2000 66.8000 202.6000 67.6000 ;
	    RECT 200.4000 65.4000 201.0000 65.8000 ;
	    RECT 200.7000 65.1000 201.0000 65.4000 ;
	    RECT 191.0000 61.8000 191.7000 62.2000 ;
	    RECT 191.3000 61.1000 191.7000 61.8000 ;
	    RECT 193.4000 61.5000 193.8000 63.5000 ;
	    RECT 194.2000 64.8000 195.4000 65.1000 ;
	    RECT 196.2000 64.8000 197.2000 65.1000 ;
	    RECT 194.2000 61.1000 194.6000 64.8000 ;
	    RECT 195.0000 64.7000 195.4000 64.8000 ;
	    RECT 196.4000 61.1000 197.2000 64.8000 ;
	    RECT 198.3000 64.8000 199.4000 65.1000 ;
	    RECT 198.3000 64.7000 198.7000 64.8000 ;
	    RECT 199.0000 61.1000 199.4000 64.8000 ;
	    RECT 199.8000 61.1000 200.2000 65.1000 ;
	    RECT 200.7000 64.8000 201.8000 65.1000 ;
	    RECT 201.4000 61.1000 201.8000 64.8000 ;
	    RECT 203.0000 61.1000 203.4000 67.9000 ;
	    RECT 203.8000 65.1000 204.2000 65.2000 ;
	    RECT 204.6000 65.1000 205.0000 69.9000 ;
	    RECT 205.4000 67.8000 205.8000 68.6000 ;
	    RECT 206.2000 67.1000 206.6000 67.2000 ;
	    RECT 207.0000 67.1000 207.4000 69.9000 ;
	    RECT 209.4000 68.9000 209.8000 69.9000 ;
	    RECT 208.6000 67.8000 209.0000 68.6000 ;
	    RECT 206.2000 66.8000 207.4000 67.1000 ;
	    RECT 207.8000 67.1000 208.2000 67.6000 ;
	    RECT 209.5000 67.2000 209.8000 68.9000 ;
	    RECT 209.4000 67.1000 209.8000 67.2000 ;
	    RECT 207.8000 66.8000 209.8000 67.1000 ;
	    RECT 203.8000 64.8000 205.0000 65.1000 ;
	    RECT 203.8000 64.4000 204.2000 64.8000 ;
	    RECT 204.6000 61.1000 205.0000 64.8000 ;
	    RECT 207.0000 61.1000 207.4000 66.8000 ;
	    RECT 209.5000 65.1000 209.8000 66.8000 ;
	    RECT 213.4000 68.9000 213.8000 69.9000 ;
	    RECT 213.4000 67.2000 213.7000 68.9000 ;
	    RECT 214.2000 67.8000 214.6000 68.6000 ;
	    RECT 213.4000 66.8000 213.8000 67.2000 ;
	    RECT 215.6000 67.1000 216.0000 69.9000 ;
	    RECT 219.5000 69.2000 219.9000 69.9000 ;
	    RECT 219.5000 68.8000 220.2000 69.2000 ;
	    RECT 219.5000 68.2000 219.9000 68.8000 ;
	    RECT 220.7000 68.2000 221.1000 68.6000 ;
	    RECT 219.0000 67.9000 219.9000 68.2000 ;
	    RECT 215.1000 66.9000 216.0000 67.1000 ;
	    RECT 215.1000 66.8000 215.9000 66.9000 ;
	    RECT 218.2000 66.8000 218.6000 67.6000 ;
	    RECT 210.2000 65.4000 210.6000 66.2000 ;
	    RECT 212.6000 65.4000 213.0000 66.2000 ;
	    RECT 213.4000 66.1000 213.7000 66.8000 ;
	    RECT 214.2000 66.1000 214.6000 66.2000 ;
	    RECT 213.4000 65.8000 214.6000 66.1000 ;
	    RECT 213.4000 65.1000 213.7000 65.8000 ;
	    RECT 215.1000 65.2000 215.4000 66.8000 ;
	    RECT 216.2000 65.8000 217.0000 66.2000 ;
	    RECT 209.4000 64.7000 210.3000 65.1000 ;
	    RECT 209.9000 64.1000 210.3000 64.7000 ;
	    RECT 212.9000 64.7000 213.8000 65.1000 ;
	    RECT 215.0000 64.8000 215.4000 65.2000 ;
	    RECT 217.4000 65.1000 217.8000 65.6000 ;
	    RECT 218.2000 65.1000 218.6000 65.2000 ;
	    RECT 217.4000 64.8000 218.6000 65.1000 ;
	    RECT 211.0000 64.1000 211.4000 64.2000 ;
	    RECT 209.9000 63.8000 211.4000 64.1000 ;
	    RECT 209.9000 61.1000 210.3000 63.8000 ;
	    RECT 212.9000 61.1000 213.3000 64.7000 ;
	    RECT 215.1000 63.5000 215.4000 64.8000 ;
	    RECT 215.8000 63.8000 216.2000 64.6000 ;
	    RECT 215.1000 63.2000 216.9000 63.5000 ;
	    RECT 215.1000 63.1000 215.4000 63.2000 ;
	    RECT 215.0000 61.1000 215.4000 63.1000 ;
	    RECT 216.6000 63.1000 216.9000 63.2000 ;
	    RECT 216.6000 61.1000 217.0000 63.1000 ;
	    RECT 219.0000 61.1000 219.4000 67.9000 ;
	    RECT 220.6000 67.8000 221.0000 68.2000 ;
	    RECT 221.4000 67.9000 221.8000 69.9000 ;
	    RECT 223.8000 68.0000 224.2000 69.9000 ;
	    RECT 225.4000 68.0000 225.8000 69.9000 ;
	    RECT 223.8000 67.9000 225.8000 68.0000 ;
	    RECT 226.2000 67.9000 226.6000 69.9000 ;
	    RECT 228.3000 69.2000 228.7000 69.9000 ;
	    RECT 227.8000 68.8000 228.7000 69.2000 ;
	    RECT 228.3000 68.2000 228.7000 68.8000 ;
	    RECT 227.8000 67.9000 228.7000 68.2000 ;
	    RECT 229.4000 67.9000 229.8000 69.9000 ;
	    RECT 230.2000 68.0000 230.6000 69.9000 ;
	    RECT 231.8000 68.0000 232.2000 69.9000 ;
	    RECT 230.2000 67.9000 232.2000 68.0000 ;
	    RECT 221.5000 66.2000 221.8000 67.9000 ;
	    RECT 223.9000 67.7000 225.7000 67.9000 ;
	    RECT 224.2000 67.2000 224.6000 67.4000 ;
	    RECT 226.2000 67.2000 226.5000 67.9000 ;
	    RECT 222.2000 66.4000 222.6000 67.2000 ;
	    RECT 223.8000 66.9000 224.6000 67.2000 ;
	    RECT 223.8000 66.8000 224.2000 66.9000 ;
	    RECT 225.3000 66.8000 226.6000 67.2000 ;
	    RECT 227.0000 66.8000 227.4000 67.6000 ;
	    RECT 220.6000 66.1000 221.0000 66.2000 ;
	    RECT 221.4000 66.1000 221.8000 66.2000 ;
	    RECT 223.0000 66.1000 223.4000 66.2000 ;
	    RECT 223.8000 66.1000 224.2000 66.2000 ;
	    RECT 220.6000 65.8000 221.8000 66.1000 ;
	    RECT 222.6000 65.8000 224.2000 66.1000 ;
	    RECT 224.6000 65.8000 225.0000 66.6000 ;
	    RECT 219.8000 64.4000 220.2000 65.2000 ;
	    RECT 220.7000 65.1000 221.0000 65.8000 ;
	    RECT 222.6000 65.6000 223.0000 65.8000 ;
	    RECT 225.3000 65.2000 225.6000 66.8000 ;
	    RECT 220.6000 61.1000 221.0000 65.1000 ;
	    RECT 221.4000 64.8000 223.4000 65.1000 ;
	    RECT 224.6000 64.8000 225.6000 65.2000 ;
	    RECT 226.2000 65.1000 226.6000 65.2000 ;
	    RECT 227.0000 65.1000 227.4000 65.2000 ;
	    RECT 225.9000 64.8000 227.4000 65.1000 ;
	    RECT 221.4000 61.1000 221.8000 64.8000 ;
	    RECT 223.0000 61.1000 223.4000 64.8000 ;
	    RECT 225.1000 61.1000 225.5000 64.8000 ;
	    RECT 225.9000 64.2000 226.2000 64.8000 ;
	    RECT 225.8000 63.8000 226.2000 64.2000 ;
	    RECT 227.8000 61.1000 228.2000 67.9000 ;
	    RECT 229.5000 67.2000 229.8000 67.9000 ;
	    RECT 230.3000 67.7000 232.1000 67.9000 ;
	    RECT 232.6000 67.8000 233.0000 68.6000 ;
	    RECT 231.4000 67.2000 231.8000 67.4000 ;
	    RECT 229.4000 66.8000 230.7000 67.2000 ;
	    RECT 231.4000 67.1000 232.2000 67.2000 ;
	    RECT 232.6000 67.1000 233.0000 67.2000 ;
	    RECT 231.4000 66.9000 233.0000 67.1000 ;
	    RECT 231.8000 66.8000 233.0000 66.9000 ;
	    RECT 228.6000 64.4000 229.0000 65.2000 ;
	    RECT 229.4000 65.1000 229.8000 65.2000 ;
	    RECT 230.4000 65.1000 230.7000 66.8000 ;
	    RECT 231.0000 65.8000 231.4000 66.6000 ;
	    RECT 233.4000 65.1000 233.8000 69.9000 ;
	    RECT 234.2000 67.9000 234.6000 69.9000 ;
	    RECT 235.0000 68.0000 235.4000 69.9000 ;
	    RECT 236.6000 68.0000 237.0000 69.9000 ;
	    RECT 235.0000 67.9000 237.0000 68.0000 ;
	    RECT 237.4000 68.0000 237.8000 69.9000 ;
	    RECT 239.0000 68.0000 239.4000 69.9000 ;
	    RECT 237.4000 67.9000 239.4000 68.0000 ;
	    RECT 239.8000 67.9000 240.2000 69.9000 ;
	    RECT 242.2000 67.9000 242.6000 69.9000 ;
	    RECT 242.9000 68.2000 243.3000 68.6000 ;
	    RECT 234.3000 67.2000 234.6000 67.9000 ;
	    RECT 235.1000 67.7000 236.9000 67.9000 ;
	    RECT 237.5000 67.7000 239.3000 67.9000 ;
	    RECT 236.2000 67.2000 236.6000 67.4000 ;
	    RECT 237.8000 67.2000 238.2000 67.4000 ;
	    RECT 239.8000 67.2000 240.1000 67.9000 ;
	    RECT 234.2000 66.8000 235.5000 67.2000 ;
	    RECT 236.2000 66.9000 237.0000 67.2000 ;
	    RECT 236.6000 66.8000 237.0000 66.9000 ;
	    RECT 237.4000 66.9000 238.2000 67.2000 ;
	    RECT 237.4000 66.8000 237.8000 66.9000 ;
	    RECT 238.9000 66.8000 240.2000 67.2000 ;
	    RECT 234.2000 65.1000 234.6000 65.2000 ;
	    RECT 235.2000 65.1000 235.5000 66.8000 ;
	    RECT 235.8000 65.8000 236.2000 66.6000 ;
	    RECT 238.2000 65.8000 238.6000 66.6000 ;
	    RECT 238.9000 66.1000 239.2000 66.8000 ;
	    RECT 241.4000 66.4000 241.8000 67.2000 ;
	    RECT 240.6000 66.1000 241.0000 66.2000 ;
	    RECT 242.2000 66.1000 242.5000 67.9000 ;
	    RECT 243.0000 67.8000 243.4000 68.2000 ;
	    RECT 243.8000 67.8000 244.2000 68.6000 ;
	    RECT 243.0000 66.1000 243.4000 66.2000 ;
	    RECT 238.9000 65.8000 241.4000 66.1000 ;
	    RECT 242.2000 65.8000 243.4000 66.1000 ;
	    RECT 238.9000 65.1000 239.2000 65.8000 ;
	    RECT 241.0000 65.6000 241.4000 65.8000 ;
	    RECT 239.8000 65.1000 240.2000 65.2000 ;
	    RECT 243.0000 65.1000 243.3000 65.8000 ;
	    RECT 229.4000 64.8000 230.1000 65.1000 ;
	    RECT 230.4000 64.8000 230.9000 65.1000 ;
	    RECT 229.8000 64.2000 230.1000 64.8000 ;
	    RECT 229.8000 63.8000 230.2000 64.2000 ;
	    RECT 230.5000 61.1000 230.9000 64.8000 ;
	    RECT 233.4000 64.8000 234.9000 65.1000 ;
	    RECT 235.2000 64.8000 235.7000 65.1000 ;
	    RECT 233.4000 61.1000 233.8000 64.8000 ;
	    RECT 234.6000 64.2000 234.9000 64.8000 ;
	    RECT 234.6000 63.8000 235.0000 64.2000 ;
	    RECT 235.3000 61.1000 235.7000 64.8000 ;
	    RECT 238.7000 64.8000 239.2000 65.1000 ;
	    RECT 239.5000 64.8000 240.2000 65.1000 ;
	    RECT 240.6000 64.8000 242.6000 65.1000 ;
	    RECT 238.7000 61.1000 239.1000 64.8000 ;
	    RECT 239.5000 64.2000 239.8000 64.8000 ;
	    RECT 239.4000 63.8000 239.8000 64.2000 ;
	    RECT 240.6000 61.1000 241.0000 64.8000 ;
	    RECT 242.2000 61.1000 242.6000 64.8000 ;
	    RECT 243.0000 61.1000 243.4000 65.1000 ;
	    RECT 244.6000 61.1000 245.0000 69.9000 ;
	    RECT 245.4000 67.8000 245.8000 68.6000 ;
	    RECT 246.2000 65.1000 246.6000 69.9000 ;
	    RECT 247.8000 67.8000 248.2000 68.2000 ;
	    RECT 247.8000 67.1000 248.1000 67.8000 ;
	    RECT 248.8000 67.1000 249.2000 69.9000 ;
	    RECT 251.0000 68.9000 251.4000 69.9000 ;
	    RECT 251.0000 67.2000 251.3000 68.9000 ;
	    RECT 251.8000 67.8000 252.2000 68.6000 ;
	    RECT 252.6000 68.0000 253.0000 69.9000 ;
	    RECT 254.2000 68.0000 254.6000 69.9000 ;
	    RECT 252.6000 67.9000 254.6000 68.0000 ;
	    RECT 255.0000 67.9000 255.4000 69.9000 ;
	    RECT 252.7000 67.7000 254.5000 67.9000 ;
	    RECT 253.0000 67.2000 253.4000 67.4000 ;
	    RECT 255.0000 67.2000 255.3000 67.9000 ;
	    RECT 247.8000 66.8000 249.7000 67.1000 ;
	    RECT 247.8000 65.8000 248.6000 66.2000 ;
	    RECT 247.0000 65.1000 247.4000 65.6000 ;
	    RECT 246.2000 64.8000 247.4000 65.1000 ;
	    RECT 249.4000 65.2000 249.7000 66.8000 ;
	    RECT 251.0000 66.8000 251.4000 67.2000 ;
	    RECT 252.6000 66.9000 253.4000 67.2000 ;
	    RECT 252.6000 66.8000 253.0000 66.9000 ;
	    RECT 254.1000 66.8000 255.4000 67.2000 ;
	    RECT 251.0000 66.2000 251.3000 66.8000 ;
	    RECT 250.2000 65.4000 250.6000 66.2000 ;
	    RECT 251.0000 65.8000 251.4000 66.2000 ;
	    RECT 251.8000 66.1000 252.2000 66.2000 ;
	    RECT 253.4000 66.1000 253.8000 66.6000 ;
	    RECT 251.8000 65.8000 253.8000 66.1000 ;
	    RECT 249.4000 64.8000 249.8000 65.2000 ;
	    RECT 251.0000 65.1000 251.3000 65.8000 ;
	    RECT 254.1000 65.1000 254.4000 66.8000 ;
	    RECT 255.0000 65.1000 255.4000 65.2000 ;
	    RECT 255.8000 65.1000 256.2000 69.9000 ;
	    RECT 257.4000 67.9000 257.8000 69.9000 ;
	    RECT 259.6000 69.2000 260.4000 69.9000 ;
	    RECT 259.0000 68.8000 260.4000 69.2000 ;
	    RECT 259.6000 68.1000 260.4000 68.8000 ;
	    RECT 257.4000 67.6000 258.5000 67.9000 ;
	    RECT 259.0000 67.7000 259.8000 67.8000 ;
	    RECT 258.1000 67.5000 258.5000 67.6000 ;
	    RECT 258.8000 67.4000 259.8000 67.7000 ;
	    RECT 258.8000 67.2000 259.1000 67.4000 ;
	    RECT 257.4000 66.9000 259.1000 67.2000 ;
	    RECT 257.4000 66.8000 258.2000 66.9000 ;
	    RECT 259.4000 66.7000 259.8000 67.1000 ;
	    RECT 259.4000 66.4000 259.7000 66.7000 ;
	    RECT 258.4000 66.1000 259.7000 66.4000 ;
	    RECT 260.1000 66.4000 260.4000 68.1000 ;
	    RECT 262.2000 67.9000 262.6000 69.9000 ;
	    RECT 263.8000 68.2000 264.2000 69.9000 ;
	    RECT 260.7000 67.4000 261.1000 67.8000 ;
	    RECT 261.4000 67.6000 262.6000 67.9000 ;
	    RECT 263.7000 67.9000 264.2000 68.2000 ;
	    RECT 261.4000 67.5000 261.8000 67.6000 ;
	    RECT 260.8000 67.2000 261.1000 67.4000 ;
	    RECT 263.7000 67.2000 264.0000 67.9000 ;
	    RECT 265.4000 67.6000 265.8000 69.9000 ;
	    RECT 264.5000 67.3000 265.8000 67.6000 ;
	    RECT 266.2000 67.6000 266.6000 69.9000 ;
	    RECT 267.8000 68.2000 268.2000 69.9000 ;
	    RECT 267.8000 67.9000 268.3000 68.2000 ;
	    RECT 266.2000 67.3000 267.5000 67.6000 ;
	    RECT 260.8000 66.8000 261.2000 67.2000 ;
	    RECT 263.7000 67.1000 264.2000 67.2000 ;
	    RECT 263.0000 66.8000 264.2000 67.1000 ;
	    RECT 260.1000 66.2000 260.6000 66.4000 ;
	    RECT 263.0000 66.2000 263.3000 66.8000 ;
	    RECT 260.1000 66.1000 261.0000 66.2000 ;
	    RECT 258.4000 66.0000 258.8000 66.1000 ;
	    RECT 260.3000 65.8000 261.0000 66.1000 ;
	    RECT 263.0000 65.8000 263.4000 66.2000 ;
	    RECT 259.5000 65.7000 259.9000 65.8000 ;
	    RECT 258.2000 65.4000 259.9000 65.7000 ;
	    RECT 258.2000 65.1000 258.5000 65.4000 ;
	    RECT 260.3000 65.1000 260.6000 65.8000 ;
	    RECT 263.7000 65.1000 264.0000 66.8000 ;
	    RECT 264.5000 66.5000 264.8000 67.3000 ;
	    RECT 264.3000 66.1000 264.8000 66.5000 ;
	    RECT 264.5000 65.1000 264.8000 66.1000 ;
	    RECT 265.3000 66.2000 265.7000 66.6000 ;
	    RECT 266.3000 66.2000 266.7000 66.6000 ;
	    RECT 265.3000 66.1000 265.8000 66.2000 ;
	    RECT 266.2000 66.1000 266.7000 66.2000 ;
	    RECT 265.3000 65.8000 266.7000 66.1000 ;
	    RECT 267.2000 66.5000 267.5000 67.3000 ;
	    RECT 268.0000 67.2000 268.3000 67.9000 ;
	    RECT 267.8000 66.8000 268.3000 67.2000 ;
	    RECT 267.2000 66.1000 267.7000 66.5000 ;
	    RECT 267.2000 65.1000 267.5000 66.1000 ;
	    RECT 268.0000 65.1000 268.3000 66.8000 ;
	    RECT 246.2000 61.1000 246.6000 64.8000 ;
	    RECT 248.6000 63.8000 249.0000 64.6000 ;
	    RECT 249.4000 63.5000 249.7000 64.8000 ;
	    RECT 247.9000 63.2000 249.7000 63.5000 ;
	    RECT 247.9000 63.1000 248.2000 63.2000 ;
	    RECT 247.8000 61.1000 248.2000 63.1000 ;
	    RECT 249.4000 63.1000 249.7000 63.2000 ;
	    RECT 250.5000 64.7000 251.4000 65.1000 ;
	    RECT 253.9000 64.8000 254.4000 65.1000 ;
	    RECT 254.7000 64.8000 256.2000 65.1000 ;
	    RECT 249.4000 61.1000 249.8000 63.1000 ;
	    RECT 250.5000 61.1000 250.9000 64.7000 ;
	    RECT 253.9000 61.1000 254.3000 64.8000 ;
	    RECT 254.7000 64.2000 255.0000 64.8000 ;
	    RECT 254.6000 63.8000 255.0000 64.2000 ;
	    RECT 255.8000 61.1000 256.2000 64.8000 ;
	    RECT 257.4000 64.8000 258.5000 65.1000 ;
	    RECT 257.4000 61.1000 257.8000 64.8000 ;
	    RECT 258.1000 64.7000 258.5000 64.8000 ;
	    RECT 259.6000 64.8000 260.6000 65.1000 ;
	    RECT 261.4000 64.8000 262.6000 65.1000 ;
	    RECT 259.6000 61.1000 260.4000 64.8000 ;
	    RECT 261.4000 64.7000 261.8000 64.8000 ;
	    RECT 262.2000 61.1000 262.6000 64.8000 ;
	    RECT 263.7000 64.6000 264.2000 65.1000 ;
	    RECT 264.5000 64.8000 265.8000 65.1000 ;
	    RECT 263.8000 61.1000 264.2000 64.6000 ;
	    RECT 265.4000 61.1000 265.8000 64.8000 ;
	    RECT 266.2000 64.8000 267.5000 65.1000 ;
	    RECT 266.2000 61.1000 266.6000 64.8000 ;
	    RECT 267.8000 64.6000 268.3000 65.1000 ;
	    RECT 267.8000 61.1000 268.2000 64.6000 ;
	    RECT 0.6000 56.2000 1.0000 59.9000 ;
	    RECT 1.3000 56.2000 1.7000 56.3000 ;
	    RECT 0.6000 55.9000 1.7000 56.2000 ;
	    RECT 2.8000 56.2000 3.6000 59.9000 ;
	    RECT 4.6000 56.2000 5.0000 56.3000 ;
	    RECT 5.4000 56.2000 5.8000 59.9000 ;
	    RECT 2.8000 55.9000 4.2000 56.2000 ;
	    RECT 4.6000 55.9000 5.8000 56.2000 ;
	    RECT 1.4000 55.6000 1.7000 55.9000 ;
	    RECT 3.5000 55.8000 4.2000 55.9000 ;
	    RECT 1.4000 55.3000 3.1000 55.6000 ;
	    RECT 2.7000 55.2000 3.1000 55.3000 ;
	    RECT 3.5000 55.2000 3.8000 55.8000 ;
	    RECT 1.6000 54.9000 2.0000 55.0000 ;
	    RECT 3.5000 54.9000 4.2000 55.2000 ;
	    RECT 1.6000 54.6000 2.9000 54.9000 ;
	    RECT 2.6000 54.3000 2.9000 54.6000 ;
	    RECT 3.3000 54.8000 4.2000 54.9000 ;
	    RECT 7.0000 55.1000 7.4000 59.9000 ;
	    RECT 8.1000 59.2000 8.5000 59.9000 ;
	    RECT 8.1000 58.8000 9.0000 59.2000 ;
	    RECT 8.1000 56.3000 8.5000 58.8000 ;
	    RECT 8.1000 55.9000 9.0000 56.3000 ;
	    RECT 7.8000 55.1000 8.2000 55.6000 ;
	    RECT 7.0000 54.8000 8.2000 55.1000 ;
	    RECT 3.3000 54.6000 3.8000 54.8000 ;
	    RECT 2.6000 53.9000 3.0000 54.3000 ;
	    RECT 1.3000 53.4000 1.7000 53.5000 ;
	    RECT 0.6000 53.1000 1.7000 53.4000 ;
	    RECT 0.6000 51.1000 1.0000 53.1000 ;
	    RECT 3.3000 52.9000 3.6000 54.6000 ;
	    RECT 4.6000 53.4000 5.0000 53.5000 ;
	    RECT 4.6000 53.1000 5.8000 53.4000 ;
	    RECT 2.8000 51.1000 3.6000 52.9000 ;
	    RECT 5.4000 51.1000 5.8000 53.1000 ;
	    RECT 7.0000 51.1000 7.4000 54.8000 ;
	    RECT 8.6000 54.2000 8.9000 55.9000 ;
	    RECT 11.0000 55.1000 11.4000 59.9000 ;
	    RECT 12.2000 56.8000 12.6000 57.2000 ;
	    RECT 12.2000 56.2000 12.5000 56.8000 ;
	    RECT 12.9000 56.2000 13.3000 59.9000 ;
	    RECT 11.8000 55.9000 12.5000 56.2000 ;
	    RECT 12.8000 55.9000 13.3000 56.2000 ;
	    RECT 11.8000 55.8000 12.2000 55.9000 ;
	    RECT 12.8000 55.2000 13.1000 55.9000 ;
	    RECT 11.8000 55.1000 12.2000 55.2000 ;
	    RECT 11.0000 54.8000 12.2000 55.1000 ;
	    RECT 12.6000 54.8000 13.1000 55.2000 ;
	    RECT 8.6000 53.8000 9.0000 54.2000 ;
	    RECT 8.6000 52.1000 8.9000 53.8000 ;
	    RECT 10.2000 52.4000 10.6000 53.2000 ;
	    RECT 8.6000 51.1000 9.0000 52.1000 ;
	    RECT 11.0000 51.1000 11.4000 54.8000 ;
	    RECT 12.8000 54.2000 13.1000 54.8000 ;
	    RECT 13.4000 54.4000 13.8000 55.2000 ;
	    RECT 15.8000 55.1000 16.2000 59.9000 ;
	    RECT 17.9000 56.3000 18.3000 59.9000 ;
	    RECT 17.4000 55.9000 18.3000 56.3000 ;
	    RECT 19.0000 55.9000 19.4000 59.9000 ;
	    RECT 19.8000 56.2000 20.2000 59.9000 ;
	    RECT 21.4000 56.2000 21.8000 59.9000 ;
	    RECT 19.8000 55.9000 21.8000 56.2000 ;
	    RECT 15.8000 54.8000 16.9000 55.1000 ;
	    RECT 11.8000 53.8000 13.1000 54.2000 ;
	    RECT 14.2000 54.1000 14.6000 54.2000 ;
	    RECT 13.8000 53.8000 14.6000 54.1000 ;
	    RECT 11.9000 53.1000 12.2000 53.8000 ;
	    RECT 13.8000 53.6000 14.2000 53.8000 ;
	    RECT 12.7000 53.1000 14.5000 53.3000 ;
	    RECT 11.8000 51.1000 12.2000 53.1000 ;
	    RECT 12.6000 53.0000 14.6000 53.1000 ;
	    RECT 12.6000 51.1000 13.0000 53.0000 ;
	    RECT 14.2000 51.1000 14.6000 53.0000 ;
	    RECT 15.8000 51.1000 16.2000 54.8000 ;
	    RECT 16.6000 54.2000 16.9000 54.8000 ;
	    RECT 17.5000 54.2000 17.8000 55.9000 ;
	    RECT 18.2000 54.8000 18.6000 55.6000 ;
	    RECT 19.1000 55.2000 19.4000 55.9000 ;
	    RECT 22.2000 55.8000 22.6000 56.6000 ;
	    RECT 21.0000 55.2000 21.4000 55.4000 ;
	    RECT 19.0000 54.9000 20.2000 55.2000 ;
	    RECT 21.0000 55.1000 21.8000 55.2000 ;
	    RECT 23.0000 55.1000 23.4000 59.9000 ;
	    RECT 24.6000 56.2000 25.0000 59.9000 ;
	    RECT 26.8000 59.2000 27.6000 59.9000 ;
	    RECT 26.2000 58.8000 27.6000 59.2000 ;
	    RECT 25.3000 56.2000 25.7000 56.3000 ;
	    RECT 24.6000 55.9000 25.7000 56.2000 ;
	    RECT 26.8000 56.2000 27.6000 58.8000 ;
	    RECT 28.6000 56.2000 29.0000 56.3000 ;
	    RECT 29.4000 56.2000 29.8000 59.9000 ;
	    RECT 30.6000 56.8000 31.0000 57.2000 ;
	    RECT 30.6000 56.2000 30.9000 56.8000 ;
	    RECT 31.3000 56.2000 31.7000 59.9000 ;
	    RECT 26.8000 55.9000 27.8000 56.2000 ;
	    RECT 28.6000 55.9000 29.8000 56.2000 ;
	    RECT 30.2000 55.9000 30.9000 56.2000 ;
	    RECT 31.2000 55.9000 31.7000 56.2000 ;
	    RECT 34.2000 56.1000 34.6000 59.9000 ;
	    RECT 35.0000 56.1000 35.4000 56.6000 ;
	    RECT 25.4000 55.6000 25.7000 55.9000 ;
	    RECT 25.4000 55.3000 27.1000 55.6000 ;
	    RECT 26.7000 55.2000 27.1000 55.3000 ;
	    RECT 27.5000 55.2000 27.8000 55.9000 ;
	    RECT 30.2000 55.8000 30.6000 55.9000 ;
	    RECT 31.2000 55.2000 31.5000 55.9000 ;
	    RECT 34.2000 55.8000 35.4000 56.1000 ;
	    RECT 21.0000 54.9000 23.4000 55.1000 ;
	    RECT 19.0000 54.8000 19.4000 54.9000 ;
	    RECT 16.6000 53.8000 17.0000 54.2000 ;
	    RECT 17.4000 53.8000 17.8000 54.2000 ;
	    RECT 17.5000 53.1000 17.8000 53.8000 ;
	    RECT 19.0000 53.1000 19.4000 53.2000 ;
	    RECT 19.9000 53.1000 20.2000 54.9000 ;
	    RECT 21.4000 54.8000 23.4000 54.9000 ;
	    RECT 20.6000 53.8000 21.0000 54.6000 ;
	    RECT 23.0000 53.1000 23.4000 54.8000 ;
	    RECT 25.6000 54.9000 26.0000 55.0000 ;
	    RECT 27.5000 54.9000 28.2000 55.2000 ;
	    RECT 25.6000 54.6000 26.9000 54.9000 ;
	    RECT 26.6000 54.3000 26.9000 54.6000 ;
	    RECT 27.3000 54.8000 28.2000 54.9000 ;
	    RECT 31.0000 54.8000 31.5000 55.2000 ;
	    RECT 27.3000 54.6000 27.8000 54.8000 ;
	    RECT 26.6000 53.9000 27.0000 54.3000 ;
	    RECT 25.3000 53.4000 25.7000 53.5000 ;
	    RECT 17.4000 52.8000 19.4000 53.1000 ;
	    RECT 17.5000 52.1000 17.8000 52.8000 ;
	    RECT 19.1000 52.4000 19.5000 52.8000 ;
	    RECT 17.4000 51.1000 17.8000 52.1000 ;
	    RECT 19.8000 51.1000 20.2000 53.1000 ;
	    RECT 22.5000 52.8000 23.4000 53.1000 ;
	    RECT 24.6000 53.1000 25.7000 53.4000 ;
	    RECT 22.5000 51.1000 22.9000 52.8000 ;
	    RECT 24.6000 51.1000 25.0000 53.1000 ;
	    RECT 27.3000 52.9000 27.6000 54.6000 ;
	    RECT 31.2000 54.2000 31.5000 54.8000 ;
	    RECT 31.8000 54.4000 32.2000 55.2000 ;
	    RECT 29.0000 53.8000 29.8000 54.2000 ;
	    RECT 30.2000 53.8000 31.5000 54.2000 ;
	    RECT 32.6000 54.1000 33.0000 54.2000 ;
	    RECT 32.2000 53.8000 33.0000 54.1000 ;
	    RECT 28.6000 53.4000 29.0000 53.5000 ;
	    RECT 28.6000 53.1000 29.8000 53.4000 ;
	    RECT 30.3000 53.1000 30.6000 53.8000 ;
	    RECT 32.2000 53.6000 32.6000 53.8000 ;
	    RECT 31.1000 53.1000 32.9000 53.3000 ;
	    RECT 26.8000 51.1000 27.6000 52.9000 ;
	    RECT 29.4000 51.1000 29.8000 53.1000 ;
	    RECT 30.2000 51.1000 30.6000 53.1000 ;
	    RECT 31.0000 53.0000 33.0000 53.1000 ;
	    RECT 31.0000 51.1000 31.4000 53.0000 ;
	    RECT 32.6000 51.1000 33.0000 53.0000 ;
	    RECT 34.2000 51.1000 34.6000 55.8000 ;
	    RECT 35.8000 53.1000 36.2000 59.9000 ;
	    RECT 37.4000 56.2000 37.8000 59.9000 ;
	    RECT 39.0000 56.2000 39.4000 59.9000 ;
	    RECT 37.4000 55.9000 39.4000 56.2000 ;
	    RECT 39.8000 55.9000 40.2000 59.9000 ;
	    RECT 40.9000 56.3000 41.3000 59.9000 ;
	    RECT 40.9000 55.9000 41.8000 56.3000 ;
	    RECT 37.8000 55.2000 38.2000 55.4000 ;
	    RECT 39.8000 55.2000 40.1000 55.9000 ;
	    RECT 37.4000 54.9000 38.2000 55.2000 ;
	    RECT 39.0000 54.9000 40.2000 55.2000 ;
	    RECT 37.4000 54.8000 37.8000 54.9000 ;
	    RECT 36.6000 53.4000 37.0000 54.2000 ;
	    RECT 38.2000 53.8000 38.6000 54.6000 ;
	    RECT 35.3000 52.8000 36.2000 53.1000 ;
	    RECT 39.0000 53.1000 39.3000 54.9000 ;
	    RECT 39.8000 54.8000 40.2000 54.9000 ;
	    RECT 40.6000 54.8000 41.0000 55.6000 ;
	    RECT 41.4000 54.2000 41.7000 55.9000 ;
	    RECT 43.0000 55.6000 43.4000 59.9000 ;
	    RECT 45.1000 57.9000 45.7000 59.9000 ;
	    RECT 47.4000 57.9000 47.8000 59.9000 ;
	    RECT 49.6000 58.2000 50.0000 59.9000 ;
	    RECT 49.6000 57.9000 50.6000 58.2000 ;
	    RECT 45.4000 57.5000 45.8000 57.9000 ;
	    RECT 47.5000 57.6000 47.8000 57.9000 ;
	    RECT 47.1000 57.3000 48.9000 57.6000 ;
	    RECT 50.2000 57.5000 50.6000 57.9000 ;
	    RECT 47.1000 57.2000 47.5000 57.3000 ;
	    RECT 48.5000 57.2000 48.9000 57.3000 ;
	    RECT 45.0000 56.6000 45.7000 57.0000 ;
	    RECT 45.4000 56.1000 45.7000 56.6000 ;
	    RECT 46.5000 56.5000 47.6000 56.8000 ;
	    RECT 46.5000 56.4000 46.9000 56.5000 ;
	    RECT 45.4000 55.8000 46.6000 56.1000 ;
	    RECT 43.0000 55.3000 45.1000 55.6000 ;
	    RECT 41.4000 53.8000 41.8000 54.2000 ;
	    RECT 39.8000 53.1000 40.2000 53.2000 ;
	    RECT 41.4000 53.1000 41.7000 53.8000 ;
	    RECT 35.3000 51.1000 35.7000 52.8000 ;
	    RECT 39.0000 51.1000 39.4000 53.1000 ;
	    RECT 39.8000 52.8000 41.7000 53.1000 ;
	    RECT 39.7000 52.4000 40.1000 52.8000 ;
	    RECT 41.4000 52.1000 41.7000 52.8000 ;
	    RECT 43.0000 53.6000 43.4000 55.3000 ;
	    RECT 44.7000 55.2000 45.1000 55.3000 ;
	    RECT 43.9000 54.9000 44.3000 55.0000 ;
	    RECT 43.9000 54.6000 45.8000 54.9000 ;
	    RECT 45.4000 54.5000 45.8000 54.6000 ;
	    RECT 46.3000 54.2000 46.6000 55.8000 ;
	    RECT 47.3000 55.9000 47.6000 56.5000 ;
	    RECT 47.9000 56.5000 48.3000 56.6000 ;
	    RECT 50.2000 56.5000 50.6000 56.6000 ;
	    RECT 47.9000 56.2000 50.6000 56.5000 ;
	    RECT 47.3000 55.7000 49.7000 55.9000 ;
	    RECT 51.8000 55.7000 52.2000 59.9000 ;
	    RECT 52.9000 56.2000 53.3000 59.9000 ;
	    RECT 47.3000 55.6000 52.2000 55.7000 ;
	    RECT 49.3000 55.5000 52.2000 55.6000 ;
	    RECT 49.4000 55.4000 52.2000 55.5000 ;
	    RECT 52.6000 55.9000 53.3000 56.2000 ;
	    RECT 52.6000 55.8000 53.0000 55.9000 ;
	    RECT 52.6000 55.2000 52.9000 55.8000 ;
	    RECT 55.0000 55.6000 55.4000 59.9000 ;
	    RECT 53.4000 55.4000 55.4000 55.6000 ;
	    RECT 53.3000 55.3000 55.4000 55.4000 ;
	    RECT 57.4000 55.6000 57.8000 59.9000 ;
	    RECT 59.5000 57.9000 60.1000 59.9000 ;
	    RECT 61.8000 57.9000 62.2000 59.9000 ;
	    RECT 64.0000 58.2000 64.4000 59.9000 ;
	    RECT 64.0000 57.9000 65.0000 58.2000 ;
	    RECT 59.8000 57.5000 60.2000 57.9000 ;
	    RECT 61.9000 57.6000 62.2000 57.9000 ;
	    RECT 61.5000 57.3000 63.3000 57.6000 ;
	    RECT 64.6000 57.5000 65.0000 57.9000 ;
	    RECT 61.5000 57.2000 61.9000 57.3000 ;
	    RECT 62.9000 57.2000 63.3000 57.3000 ;
	    RECT 59.4000 56.6000 60.1000 57.0000 ;
	    RECT 59.8000 56.1000 60.1000 56.6000 ;
	    RECT 60.9000 56.5000 62.0000 56.8000 ;
	    RECT 60.9000 56.4000 61.3000 56.5000 ;
	    RECT 59.8000 55.8000 61.0000 56.1000 ;
	    RECT 57.4000 55.3000 59.5000 55.6000 ;
	    RECT 48.6000 55.1000 49.0000 55.2000 ;
	    RECT 48.6000 54.8000 51.1000 55.1000 ;
	    RECT 49.4000 54.7000 49.8000 54.8000 ;
	    RECT 50.7000 54.7000 51.1000 54.8000 ;
	    RECT 52.6000 54.8000 53.0000 55.2000 ;
	    RECT 53.3000 55.0000 53.7000 55.3000 ;
	    RECT 49.9000 54.2000 50.3000 54.3000 ;
	    RECT 46.3000 53.9000 51.8000 54.2000 ;
	    RECT 46.5000 53.8000 46.9000 53.9000 ;
	    RECT 43.0000 53.3000 44.9000 53.6000 ;
	    RECT 41.4000 51.1000 41.8000 52.1000 ;
	    RECT 43.0000 51.1000 43.4000 53.3000 ;
	    RECT 44.5000 53.2000 44.9000 53.3000 ;
	    RECT 49.4000 52.8000 49.7000 53.9000 ;
	    RECT 51.0000 53.8000 51.8000 53.9000 ;
	    RECT 48.5000 52.7000 48.9000 52.8000 ;
	    RECT 45.4000 52.1000 45.8000 52.5000 ;
	    RECT 47.5000 52.4000 48.9000 52.7000 ;
	    RECT 49.4000 52.4000 49.8000 52.8000 ;
	    RECT 47.5000 52.1000 47.8000 52.4000 ;
	    RECT 50.2000 52.1000 50.6000 52.5000 ;
	    RECT 45.1000 51.8000 45.8000 52.1000 ;
	    RECT 45.1000 51.1000 45.7000 51.8000 ;
	    RECT 47.4000 51.1000 47.8000 52.1000 ;
	    RECT 49.6000 51.8000 50.6000 52.1000 ;
	    RECT 49.6000 51.1000 50.0000 51.8000 ;
	    RECT 51.8000 51.1000 52.2000 53.5000 ;
	    RECT 52.6000 53.1000 52.9000 54.8000 ;
	    RECT 53.3000 53.5000 53.6000 55.0000 ;
	    RECT 54.0000 54.2000 54.4000 54.6000 ;
	    RECT 54.1000 53.8000 54.6000 54.2000 ;
	    RECT 57.4000 53.6000 57.8000 55.3000 ;
	    RECT 59.1000 55.2000 59.5000 55.3000 ;
	    RECT 58.3000 54.9000 58.7000 55.0000 ;
	    RECT 58.3000 54.6000 60.2000 54.9000 ;
	    RECT 59.8000 54.5000 60.2000 54.6000 ;
	    RECT 60.7000 54.2000 61.0000 55.8000 ;
	    RECT 61.7000 55.9000 62.0000 56.5000 ;
	    RECT 62.3000 56.5000 62.7000 56.6000 ;
	    RECT 64.6000 56.5000 65.0000 56.6000 ;
	    RECT 62.3000 56.2000 65.0000 56.5000 ;
	    RECT 61.7000 55.7000 64.1000 55.9000 ;
	    RECT 66.2000 55.7000 66.6000 59.9000 ;
	    RECT 67.0000 55.9000 67.4000 59.9000 ;
	    RECT 67.8000 56.2000 68.2000 59.9000 ;
	    RECT 69.4000 56.2000 69.8000 59.9000 ;
	    RECT 71.3000 59.2000 71.7000 59.9000 ;
	    RECT 71.3000 58.8000 72.2000 59.2000 ;
	    RECT 70.6000 56.8000 71.0000 57.2000 ;
	    RECT 70.6000 56.2000 70.9000 56.8000 ;
	    RECT 71.3000 56.2000 71.7000 58.8000 ;
	    RECT 73.8000 56.8000 74.2000 57.2000 ;
	    RECT 73.8000 56.2000 74.1000 56.8000 ;
	    RECT 74.5000 56.2000 74.9000 59.9000 ;
	    RECT 67.8000 55.9000 69.8000 56.2000 ;
	    RECT 70.2000 55.9000 70.9000 56.2000 ;
	    RECT 71.2000 55.9000 71.7000 56.2000 ;
	    RECT 73.4000 55.9000 74.1000 56.2000 ;
	    RECT 74.4000 55.9000 74.9000 56.2000 ;
	    RECT 76.6000 56.2000 77.0000 59.9000 ;
	    RECT 78.2000 56.2000 78.6000 59.9000 ;
	    RECT 76.6000 55.9000 78.6000 56.2000 ;
	    RECT 79.0000 55.9000 79.4000 59.9000 ;
	    RECT 79.8000 57.9000 80.2000 59.9000 ;
	    RECT 79.9000 57.8000 80.2000 57.9000 ;
	    RECT 81.4000 57.9000 81.8000 59.9000 ;
	    RECT 81.4000 57.8000 81.7000 57.9000 ;
	    RECT 79.9000 57.5000 81.7000 57.8000 ;
	    RECT 79.9000 56.2000 80.2000 57.5000 ;
	    RECT 80.6000 56.4000 81.0000 57.2000 ;
	    RECT 61.7000 55.6000 66.6000 55.7000 ;
	    RECT 63.7000 55.5000 66.6000 55.6000 ;
	    RECT 63.8000 55.4000 66.6000 55.5000 ;
	    RECT 67.1000 55.2000 67.4000 55.9000 ;
	    RECT 70.2000 55.8000 70.6000 55.9000 ;
	    RECT 69.0000 55.2000 69.4000 55.4000 ;
	    RECT 63.0000 55.1000 63.4000 55.2000 ;
	    RECT 63.0000 54.8000 65.5000 55.1000 ;
	    RECT 67.0000 54.9000 68.2000 55.2000 ;
	    RECT 69.0000 54.9000 69.8000 55.2000 ;
	    RECT 67.0000 54.8000 67.4000 54.9000 ;
	    RECT 63.8000 54.7000 64.2000 54.8000 ;
	    RECT 65.1000 54.7000 65.5000 54.8000 ;
	    RECT 64.3000 54.2000 64.7000 54.3000 ;
	    RECT 60.7000 53.9000 66.2000 54.2000 ;
	    RECT 60.9000 53.8000 61.3000 53.9000 ;
	    RECT 62.2000 53.8000 62.6000 53.9000 ;
	    RECT 53.3000 53.2000 54.5000 53.5000 ;
	    RECT 57.4000 53.3000 59.3000 53.6000 ;
	    RECT 52.6000 51.1000 53.0000 53.1000 ;
	    RECT 54.2000 52.1000 54.5000 53.2000 ;
	    RECT 55.0000 52.4000 55.4000 53.2000 ;
	    RECT 54.2000 51.1000 54.6000 52.1000 ;
	    RECT 57.4000 51.1000 57.8000 53.3000 ;
	    RECT 58.9000 53.2000 59.3000 53.3000 ;
	    RECT 63.8000 52.8000 64.1000 53.9000 ;
	    RECT 65.4000 53.8000 66.2000 53.9000 ;
	    RECT 62.9000 52.7000 63.3000 52.8000 ;
	    RECT 59.8000 52.1000 60.2000 52.5000 ;
	    RECT 61.9000 52.4000 63.3000 52.7000 ;
	    RECT 63.8000 52.4000 64.2000 52.8000 ;
	    RECT 61.9000 52.1000 62.2000 52.4000 ;
	    RECT 64.6000 52.1000 65.0000 52.5000 ;
	    RECT 59.5000 51.8000 60.2000 52.1000 ;
	    RECT 59.5000 51.1000 60.1000 51.8000 ;
	    RECT 61.8000 51.1000 62.2000 52.1000 ;
	    RECT 64.0000 51.8000 65.0000 52.1000 ;
	    RECT 64.0000 51.1000 64.4000 51.8000 ;
	    RECT 66.2000 51.1000 66.6000 53.5000 ;
	    RECT 67.0000 52.8000 67.4000 53.2000 ;
	    RECT 67.9000 53.1000 68.2000 54.9000 ;
	    RECT 69.4000 54.8000 69.8000 54.9000 ;
	    RECT 68.6000 53.8000 69.0000 54.6000 ;
	    RECT 71.2000 54.2000 71.5000 55.9000 ;
	    RECT 73.4000 55.8000 73.8000 55.9000 ;
	    RECT 71.8000 55.1000 72.2000 55.2000 ;
	    RECT 73.4000 55.1000 73.7000 55.8000 ;
	    RECT 74.4000 55.2000 74.7000 55.9000 ;
	    RECT 77.0000 55.2000 77.4000 55.4000 ;
	    RECT 79.0000 55.2000 79.3000 55.9000 ;
	    RECT 79.8000 55.8000 80.2000 56.2000 ;
	    RECT 79.9000 55.2000 80.2000 55.8000 ;
	    RECT 71.8000 54.8000 73.7000 55.1000 ;
	    RECT 74.2000 54.8000 74.7000 55.2000 ;
	    RECT 71.8000 54.4000 72.2000 54.8000 ;
	    RECT 74.4000 54.2000 74.7000 54.8000 ;
	    RECT 75.0000 54.4000 75.4000 55.2000 ;
	    RECT 76.6000 54.9000 77.4000 55.2000 ;
	    RECT 78.2000 54.9000 79.4000 55.2000 ;
	    RECT 76.6000 54.8000 77.0000 54.9000 ;
	    RECT 70.2000 53.8000 71.5000 54.2000 ;
	    RECT 72.6000 54.1000 73.0000 54.2000 ;
	    RECT 72.2000 53.8000 73.0000 54.1000 ;
	    RECT 73.4000 53.8000 74.7000 54.2000 ;
	    RECT 75.8000 54.1000 76.2000 54.2000 ;
	    RECT 75.4000 53.8000 76.2000 54.1000 ;
	    RECT 76.6000 54.1000 77.0000 54.2000 ;
	    RECT 77.4000 54.1000 77.8000 54.6000 ;
	    RECT 76.6000 53.8000 77.8000 54.1000 ;
	    RECT 70.3000 53.1000 70.6000 53.8000 ;
	    RECT 72.2000 53.6000 72.6000 53.8000 ;
	    RECT 71.1000 53.1000 72.9000 53.3000 ;
	    RECT 73.5000 53.1000 73.8000 53.8000 ;
	    RECT 75.4000 53.6000 75.8000 53.8000 ;
	    RECT 74.3000 53.1000 76.1000 53.3000 ;
	    RECT 78.2000 53.1000 78.5000 54.9000 ;
	    RECT 79.0000 54.8000 79.4000 54.9000 ;
	    RECT 79.8000 54.8000 80.2000 55.2000 ;
	    RECT 81.0000 54.8000 81.8000 55.2000 ;
	    RECT 82.2000 54.8000 82.6000 56.2000 ;
	    RECT 83.0000 55.6000 83.4000 59.9000 ;
	    RECT 85.1000 57.9000 85.7000 59.9000 ;
	    RECT 87.4000 57.9000 87.8000 59.9000 ;
	    RECT 89.6000 58.2000 90.0000 59.9000 ;
	    RECT 89.6000 57.9000 90.6000 58.2000 ;
	    RECT 85.4000 57.5000 85.8000 57.9000 ;
	    RECT 87.5000 57.6000 87.8000 57.9000 ;
	    RECT 87.1000 57.3000 88.9000 57.6000 ;
	    RECT 90.2000 57.5000 90.6000 57.9000 ;
	    RECT 87.1000 57.2000 87.5000 57.3000 ;
	    RECT 88.5000 57.2000 88.9000 57.3000 ;
	    RECT 84.6000 57.0000 85.3000 57.2000 ;
	    RECT 84.6000 56.8000 85.7000 57.0000 ;
	    RECT 85.0000 56.6000 85.7000 56.8000 ;
	    RECT 85.4000 56.1000 85.7000 56.6000 ;
	    RECT 86.5000 56.5000 87.6000 56.8000 ;
	    RECT 86.5000 56.4000 86.9000 56.5000 ;
	    RECT 85.4000 55.8000 86.6000 56.1000 ;
	    RECT 83.0000 55.3000 85.1000 55.6000 ;
	    RECT 79.9000 54.2000 80.2000 54.8000 ;
	    RECT 79.9000 54.1000 80.7000 54.2000 ;
	    RECT 79.9000 53.9000 80.8000 54.1000 ;
	    RECT 67.1000 52.4000 67.5000 52.8000 ;
	    RECT 67.8000 51.1000 68.2000 53.1000 ;
	    RECT 70.2000 51.1000 70.6000 53.1000 ;
	    RECT 71.0000 53.0000 73.0000 53.1000 ;
	    RECT 71.0000 51.1000 71.4000 53.0000 ;
	    RECT 72.6000 51.1000 73.0000 53.0000 ;
	    RECT 73.4000 51.1000 73.8000 53.1000 ;
	    RECT 74.2000 53.0000 76.2000 53.1000 ;
	    RECT 74.2000 51.1000 74.6000 53.0000 ;
	    RECT 75.8000 51.1000 76.2000 53.0000 ;
	    RECT 78.2000 51.1000 78.6000 53.1000 ;
	    RECT 79.0000 52.8000 79.4000 53.2000 ;
	    RECT 78.9000 52.4000 79.3000 52.8000 ;
	    RECT 80.4000 51.1000 80.8000 53.9000 ;
	    RECT 83.0000 53.6000 83.4000 55.3000 ;
	    RECT 84.7000 55.2000 85.1000 55.3000 ;
	    RECT 83.9000 54.9000 84.3000 55.0000 ;
	    RECT 83.9000 54.6000 85.8000 54.9000 ;
	    RECT 85.4000 54.5000 85.8000 54.6000 ;
	    RECT 86.3000 54.2000 86.6000 55.8000 ;
	    RECT 87.3000 55.9000 87.6000 56.5000 ;
	    RECT 87.9000 56.5000 88.3000 56.6000 ;
	    RECT 90.2000 56.5000 90.6000 56.6000 ;
	    RECT 87.9000 56.2000 90.6000 56.5000 ;
	    RECT 87.3000 55.7000 89.7000 55.9000 ;
	    RECT 91.8000 55.7000 92.2000 59.9000 ;
	    RECT 93.4000 56.4000 93.8000 59.9000 ;
	    RECT 87.3000 55.6000 92.2000 55.7000 ;
	    RECT 89.3000 55.5000 92.2000 55.6000 ;
	    RECT 89.4000 55.4000 92.2000 55.5000 ;
	    RECT 93.3000 55.9000 93.8000 56.4000 ;
	    RECT 95.0000 56.2000 95.4000 59.9000 ;
	    RECT 96.6000 56.4000 97.0000 59.9000 ;
	    RECT 94.1000 55.9000 95.4000 56.2000 ;
	    RECT 96.5000 55.9000 97.0000 56.4000 ;
	    RECT 98.2000 56.2000 98.6000 59.9000 ;
	    RECT 99.8000 57.9000 100.2000 59.9000 ;
	    RECT 97.3000 55.9000 98.6000 56.2000 ;
	    RECT 88.6000 55.1000 89.0000 55.2000 ;
	    RECT 88.6000 54.8000 91.1000 55.1000 ;
	    RECT 89.4000 54.7000 89.8000 54.8000 ;
	    RECT 90.7000 54.7000 91.1000 54.8000 ;
	    RECT 89.9000 54.2000 90.3000 54.3000 ;
	    RECT 93.3000 54.2000 93.6000 55.9000 ;
	    RECT 94.1000 54.9000 94.4000 55.9000 ;
	    RECT 93.9000 54.5000 94.4000 54.9000 ;
	    RECT 86.3000 53.9000 91.8000 54.2000 ;
	    RECT 86.5000 53.8000 86.9000 53.9000 ;
	    RECT 83.0000 53.3000 84.9000 53.6000 ;
	    RECT 83.0000 51.1000 83.4000 53.3000 ;
	    RECT 84.5000 53.2000 84.9000 53.3000 ;
	    RECT 89.4000 52.8000 89.7000 53.9000 ;
	    RECT 91.0000 53.8000 91.8000 53.9000 ;
	    RECT 93.3000 53.8000 93.8000 54.2000 ;
	    RECT 88.5000 52.7000 88.9000 52.8000 ;
	    RECT 85.4000 52.1000 85.8000 52.5000 ;
	    RECT 87.5000 52.4000 88.9000 52.7000 ;
	    RECT 89.4000 52.4000 89.8000 52.8000 ;
	    RECT 87.5000 52.1000 87.8000 52.4000 ;
	    RECT 90.2000 52.1000 90.6000 52.5000 ;
	    RECT 85.1000 51.8000 85.8000 52.1000 ;
	    RECT 85.1000 51.1000 85.7000 51.8000 ;
	    RECT 87.4000 51.1000 87.8000 52.1000 ;
	    RECT 89.6000 51.8000 90.6000 52.1000 ;
	    RECT 89.6000 51.1000 90.0000 51.8000 ;
	    RECT 91.8000 51.1000 92.2000 53.5000 ;
	    RECT 93.3000 53.2000 93.6000 53.8000 ;
	    RECT 94.1000 53.7000 94.4000 54.5000 ;
	    RECT 94.9000 54.8000 95.4000 55.2000 ;
	    RECT 94.9000 54.4000 95.3000 54.8000 ;
	    RECT 96.5000 54.2000 96.8000 55.9000 ;
	    RECT 97.3000 54.9000 97.6000 55.9000 ;
	    RECT 99.9000 55.8000 100.2000 57.9000 ;
	    RECT 101.4000 55.9000 101.8000 59.9000 ;
	    RECT 99.9000 55.5000 101.1000 55.8000 ;
	    RECT 97.1000 54.5000 97.6000 54.9000 ;
	    RECT 96.5000 53.8000 97.0000 54.2000 ;
	    RECT 94.1000 53.4000 95.4000 53.7000 ;
	    RECT 93.3000 52.8000 93.8000 53.2000 ;
	    RECT 93.4000 51.1000 93.8000 52.8000 ;
	    RECT 95.0000 51.1000 95.4000 53.4000 ;
	    RECT 96.5000 53.1000 96.8000 53.8000 ;
	    RECT 97.3000 53.7000 97.6000 54.5000 ;
	    RECT 98.1000 54.8000 98.6000 55.2000 ;
	    RECT 99.8000 54.8000 100.2000 55.2000 ;
	    RECT 98.1000 54.4000 98.5000 54.8000 ;
	    RECT 99.0000 53.8000 99.4000 54.6000 ;
	    RECT 99.9000 54.4000 100.2000 54.8000 ;
	    RECT 99.9000 54.1000 100.4000 54.4000 ;
	    RECT 100.0000 54.0000 100.4000 54.1000 ;
	    RECT 100.8000 53.8000 101.1000 55.5000 ;
	    RECT 101.5000 55.2000 101.8000 55.9000 ;
	    RECT 101.4000 54.8000 101.8000 55.2000 ;
	    RECT 100.8000 53.7000 101.2000 53.8000 ;
	    RECT 97.3000 53.4000 98.6000 53.7000 ;
	    RECT 99.7000 53.5000 101.2000 53.7000 ;
	    RECT 96.5000 52.8000 97.0000 53.1000 ;
	    RECT 96.6000 51.1000 97.0000 52.8000 ;
	    RECT 98.2000 51.1000 98.6000 53.4000 ;
	    RECT 99.1000 53.4000 101.2000 53.5000 ;
	    RECT 99.1000 53.2000 100.0000 53.4000 ;
	    RECT 99.1000 53.1000 99.4000 53.2000 ;
	    RECT 101.5000 53.1000 101.8000 54.8000 ;
	    RECT 102.2000 53.4000 102.6000 54.2000 ;
	    RECT 99.0000 51.1000 99.4000 53.1000 ;
	    RECT 101.1000 52.6000 101.8000 53.1000 ;
	    RECT 103.0000 53.1000 103.4000 59.9000 ;
	    RECT 103.8000 55.8000 104.2000 56.6000 ;
	    RECT 105.4000 56.4000 105.8000 59.9000 ;
	    RECT 105.3000 55.9000 105.8000 56.4000 ;
	    RECT 107.0000 56.2000 107.4000 59.9000 ;
	    RECT 106.1000 55.9000 107.4000 56.2000 ;
	    RECT 105.3000 54.2000 105.6000 55.9000 ;
	    RECT 106.1000 54.9000 106.4000 55.9000 ;
	    RECT 109.4000 55.6000 109.8000 59.9000 ;
	    RECT 111.5000 57.9000 112.1000 59.9000 ;
	    RECT 113.8000 57.9000 114.2000 59.9000 ;
	    RECT 116.0000 58.2000 116.4000 59.9000 ;
	    RECT 116.0000 57.9000 117.0000 58.2000 ;
	    RECT 111.8000 57.5000 112.2000 57.9000 ;
	    RECT 113.9000 57.6000 114.2000 57.9000 ;
	    RECT 113.5000 57.3000 115.3000 57.6000 ;
	    RECT 116.6000 57.5000 117.0000 57.9000 ;
	    RECT 113.5000 57.2000 113.9000 57.3000 ;
	    RECT 114.9000 57.2000 115.3000 57.3000 ;
	    RECT 111.4000 56.6000 112.1000 57.0000 ;
	    RECT 111.8000 56.1000 112.1000 56.6000 ;
	    RECT 112.9000 56.5000 114.0000 56.8000 ;
	    RECT 112.9000 56.4000 113.3000 56.5000 ;
	    RECT 111.8000 55.8000 113.0000 56.1000 ;
	    RECT 109.4000 55.3000 111.5000 55.6000 ;
	    RECT 105.9000 54.5000 106.4000 54.9000 ;
	    RECT 105.3000 53.8000 105.8000 54.2000 ;
	    RECT 105.3000 53.1000 105.6000 53.8000 ;
	    RECT 106.1000 53.7000 106.4000 54.5000 ;
	    RECT 106.9000 55.1000 107.4000 55.2000 ;
	    RECT 108.6000 55.1000 109.0000 55.2000 ;
	    RECT 106.9000 54.8000 109.0000 55.1000 ;
	    RECT 106.9000 54.4000 107.3000 54.8000 ;
	    RECT 106.1000 53.4000 107.4000 53.7000 ;
	    RECT 103.0000 52.8000 103.9000 53.1000 ;
	    RECT 105.3000 52.8000 105.8000 53.1000 ;
	    RECT 101.1000 52.2000 101.5000 52.6000 ;
	    RECT 103.5000 52.2000 103.9000 52.8000 ;
	    RECT 101.1000 51.8000 101.8000 52.2000 ;
	    RECT 103.5000 51.8000 104.2000 52.2000 ;
	    RECT 101.1000 51.1000 101.5000 51.8000 ;
	    RECT 103.5000 51.1000 103.9000 51.8000 ;
	    RECT 105.4000 51.1000 105.8000 52.8000 ;
	    RECT 107.0000 51.1000 107.4000 53.4000 ;
	    RECT 109.4000 53.6000 109.8000 55.3000 ;
	    RECT 111.1000 55.2000 111.5000 55.3000 ;
	    RECT 110.3000 54.9000 110.7000 55.0000 ;
	    RECT 110.3000 54.6000 112.2000 54.9000 ;
	    RECT 111.8000 54.5000 112.2000 54.6000 ;
	    RECT 112.7000 54.2000 113.0000 55.8000 ;
	    RECT 113.7000 55.9000 114.0000 56.5000 ;
	    RECT 114.3000 56.5000 114.7000 56.6000 ;
	    RECT 116.6000 56.5000 117.0000 56.6000 ;
	    RECT 114.3000 56.2000 117.0000 56.5000 ;
	    RECT 113.7000 55.7000 116.1000 55.9000 ;
	    RECT 118.2000 55.7000 118.6000 59.9000 ;
	    RECT 119.0000 55.9000 119.4000 59.9000 ;
	    RECT 119.8000 56.2000 120.2000 59.9000 ;
	    RECT 121.4000 56.2000 121.8000 59.9000 ;
	    RECT 123.0000 57.9000 123.4000 59.9000 ;
	    RECT 123.1000 57.8000 123.4000 57.9000 ;
	    RECT 124.6000 57.9000 125.0000 59.9000 ;
	    RECT 124.6000 57.8000 124.9000 57.9000 ;
	    RECT 123.1000 57.5000 124.9000 57.8000 ;
	    RECT 123.0000 57.1000 123.4000 57.2000 ;
	    RECT 123.8000 57.1000 124.2000 57.2000 ;
	    RECT 123.0000 56.8000 124.2000 57.1000 ;
	    RECT 123.8000 56.4000 124.2000 56.8000 ;
	    RECT 124.6000 56.2000 124.9000 57.5000 ;
	    RECT 119.8000 55.9000 121.8000 56.2000 ;
	    RECT 113.7000 55.6000 118.6000 55.7000 ;
	    RECT 115.7000 55.5000 118.6000 55.6000 ;
	    RECT 115.8000 55.4000 118.6000 55.5000 ;
	    RECT 119.1000 55.2000 119.4000 55.9000 ;
	    RECT 121.0000 55.2000 121.4000 55.4000 ;
	    RECT 115.0000 55.1000 115.4000 55.2000 ;
	    RECT 115.0000 54.8000 117.5000 55.1000 ;
	    RECT 119.0000 54.9000 120.2000 55.2000 ;
	    RECT 121.0000 54.9000 121.8000 55.2000 ;
	    RECT 119.0000 54.8000 119.4000 54.9000 ;
	    RECT 119.8000 54.8000 120.2000 54.9000 ;
	    RECT 121.4000 54.8000 121.8000 54.9000 ;
	    RECT 122.2000 54.8000 122.6000 56.2000 ;
	    RECT 124.6000 55.8000 125.0000 56.2000 ;
	    RECT 123.0000 54.8000 123.8000 55.2000 ;
	    RECT 115.8000 54.7000 116.2000 54.8000 ;
	    RECT 117.1000 54.7000 117.5000 54.8000 ;
	    RECT 116.3000 54.2000 116.7000 54.3000 ;
	    RECT 110.2000 53.6000 110.6000 54.2000 ;
	    RECT 112.6000 53.9000 118.2000 54.2000 ;
	    RECT 112.6000 53.8000 113.3000 53.9000 ;
	    RECT 109.4000 53.3000 111.3000 53.6000 ;
	    RECT 109.4000 51.1000 109.8000 53.3000 ;
	    RECT 110.9000 53.2000 111.3000 53.3000 ;
	    RECT 115.8000 52.8000 116.1000 53.9000 ;
	    RECT 117.4000 53.8000 118.2000 53.9000 ;
	    RECT 114.9000 52.7000 115.3000 52.8000 ;
	    RECT 111.8000 52.1000 112.2000 52.5000 ;
	    RECT 113.9000 52.4000 115.3000 52.7000 ;
	    RECT 115.8000 52.4000 116.2000 52.8000 ;
	    RECT 113.9000 52.1000 114.2000 52.4000 ;
	    RECT 116.6000 52.1000 117.0000 52.5000 ;
	    RECT 111.5000 51.8000 112.2000 52.1000 ;
	    RECT 111.5000 51.1000 112.1000 51.8000 ;
	    RECT 113.8000 51.1000 114.2000 52.1000 ;
	    RECT 116.0000 51.8000 117.0000 52.1000 ;
	    RECT 116.0000 51.1000 116.4000 51.8000 ;
	    RECT 118.2000 51.1000 118.6000 53.5000 ;
	    RECT 119.0000 52.8000 119.4000 53.2000 ;
	    RECT 119.9000 53.1000 120.2000 54.8000 ;
	    RECT 120.6000 53.8000 121.0000 54.6000 ;
	    RECT 124.6000 54.2000 124.9000 55.8000 ;
	    RECT 123.8000 53.9000 124.9000 54.2000 ;
	    RECT 123.8000 53.8000 124.4000 53.9000 ;
	    RECT 119.1000 52.4000 119.5000 52.8000 ;
	    RECT 119.8000 51.1000 120.2000 53.1000 ;
	    RECT 124.0000 51.1000 124.4000 53.8000 ;
	    RECT 125.4000 53.4000 125.8000 54.2000 ;
	    RECT 126.2000 54.1000 126.6000 59.9000 ;
	    RECT 127.0000 57.1000 127.4000 57.2000 ;
	    RECT 127.8000 57.1000 128.2000 59.9000 ;
	    RECT 127.0000 56.8000 128.2000 57.1000 ;
	    RECT 127.0000 54.8000 127.4000 55.2000 ;
	    RECT 127.8000 55.1000 128.2000 56.8000 ;
	    RECT 129.9000 56.2000 130.3000 59.9000 ;
	    RECT 130.6000 56.8000 131.0000 57.2000 ;
	    RECT 130.7000 56.2000 131.0000 56.8000 ;
	    RECT 131.8000 56.2000 132.2000 59.9000 ;
	    RECT 133.4000 56.2000 133.8000 59.9000 ;
	    RECT 129.9000 55.9000 130.4000 56.2000 ;
	    RECT 130.7000 55.9000 131.4000 56.2000 ;
	    RECT 131.8000 55.9000 133.8000 56.2000 ;
	    RECT 134.2000 55.9000 134.6000 59.9000 ;
	    RECT 129.4000 55.1000 129.8000 55.2000 ;
	    RECT 127.8000 54.8000 129.8000 55.1000 ;
	    RECT 127.0000 54.1000 127.3000 54.8000 ;
	    RECT 126.2000 53.8000 127.3000 54.1000 ;
	    RECT 126.2000 51.1000 126.6000 53.8000 ;
	    RECT 127.0000 52.4000 127.4000 53.2000 ;
	    RECT 127.8000 51.1000 128.2000 54.8000 ;
	    RECT 129.4000 54.4000 129.8000 54.8000 ;
	    RECT 130.1000 54.2000 130.4000 55.9000 ;
	    RECT 131.0000 55.8000 131.4000 55.9000 ;
	    RECT 132.2000 55.2000 132.6000 55.4000 ;
	    RECT 134.2000 55.2000 134.5000 55.9000 ;
	    RECT 135.0000 55.7000 135.4000 59.9000 ;
	    RECT 137.2000 58.2000 137.6000 59.9000 ;
	    RECT 136.6000 57.9000 137.6000 58.2000 ;
	    RECT 139.4000 57.9000 139.8000 59.9000 ;
	    RECT 141.5000 57.9000 142.1000 59.9000 ;
	    RECT 136.6000 57.5000 137.0000 57.9000 ;
	    RECT 139.4000 57.6000 139.7000 57.9000 ;
	    RECT 138.3000 57.3000 140.1000 57.6000 ;
	    RECT 141.4000 57.5000 141.8000 57.9000 ;
	    RECT 138.3000 57.2000 138.7000 57.3000 ;
	    RECT 139.7000 57.2000 140.1000 57.3000 ;
	    RECT 136.6000 56.5000 137.0000 56.6000 ;
	    RECT 138.9000 56.5000 139.3000 56.6000 ;
	    RECT 136.6000 56.2000 139.3000 56.5000 ;
	    RECT 139.6000 56.5000 140.7000 56.8000 ;
	    RECT 139.6000 55.9000 139.9000 56.5000 ;
	    RECT 140.3000 56.4000 140.7000 56.5000 ;
	    RECT 141.5000 56.6000 142.2000 57.0000 ;
	    RECT 141.5000 56.1000 141.8000 56.6000 ;
	    RECT 137.5000 55.7000 139.9000 55.9000 ;
	    RECT 135.0000 55.6000 139.9000 55.7000 ;
	    RECT 140.6000 55.8000 141.8000 56.1000 ;
	    RECT 135.0000 55.5000 137.9000 55.6000 ;
	    RECT 135.0000 55.4000 137.8000 55.5000 ;
	    RECT 140.6000 55.2000 140.9000 55.8000 ;
	    RECT 143.8000 55.6000 144.2000 59.9000 ;
	    RECT 144.6000 57.9000 145.0000 59.9000 ;
	    RECT 144.7000 57.8000 145.0000 57.9000 ;
	    RECT 146.2000 57.9000 146.6000 59.9000 ;
	    RECT 148.6000 57.9000 149.0000 59.9000 ;
	    RECT 146.2000 57.8000 146.5000 57.9000 ;
	    RECT 144.7000 57.5000 146.5000 57.8000 ;
	    RECT 148.7000 57.8000 149.0000 57.9000 ;
	    RECT 150.2000 57.9000 150.6000 59.9000 ;
	    RECT 150.2000 57.8000 150.5000 57.9000 ;
	    RECT 148.7000 57.5000 150.5000 57.8000 ;
	    RECT 144.7000 56.2000 145.0000 57.5000 ;
	    RECT 145.4000 57.1000 145.8000 57.2000 ;
	    RECT 149.4000 57.1000 149.8000 57.2000 ;
	    RECT 145.4000 56.8000 149.8000 57.1000 ;
	    RECT 145.4000 56.4000 145.8000 56.8000 ;
	    RECT 149.4000 56.4000 149.8000 56.8000 ;
	    RECT 150.2000 56.2000 150.5000 57.5000 ;
	    RECT 144.6000 55.8000 145.0000 56.2000 ;
	    RECT 142.1000 55.3000 144.2000 55.6000 ;
	    RECT 142.1000 55.2000 142.5000 55.3000 ;
	    RECT 131.8000 54.9000 132.6000 55.2000 ;
	    RECT 133.4000 54.9000 134.6000 55.2000 ;
	    RECT 138.2000 55.1000 138.6000 55.2000 ;
	    RECT 131.8000 54.8000 132.2000 54.9000 ;
	    RECT 128.6000 54.1000 129.0000 54.2000 ;
	    RECT 130.1000 54.1000 131.4000 54.2000 ;
	    RECT 131.8000 54.1000 132.2000 54.2000 ;
	    RECT 128.6000 53.8000 129.4000 54.1000 ;
	    RECT 130.1000 53.8000 132.2000 54.1000 ;
	    RECT 132.6000 53.8000 133.0000 54.6000 ;
	    RECT 129.0000 53.6000 129.4000 53.8000 ;
	    RECT 128.7000 53.1000 130.5000 53.3000 ;
	    RECT 131.0000 53.1000 131.3000 53.8000 ;
	    RECT 133.4000 53.1000 133.7000 54.9000 ;
	    RECT 134.2000 54.8000 134.6000 54.9000 ;
	    RECT 136.1000 54.8000 138.6000 55.1000 ;
	    RECT 140.6000 54.8000 141.0000 55.2000 ;
	    RECT 142.9000 54.9000 143.3000 55.0000 ;
	    RECT 134.2000 54.2000 134.5000 54.8000 ;
	    RECT 136.1000 54.7000 136.5000 54.8000 ;
	    RECT 137.4000 54.7000 137.8000 54.8000 ;
	    RECT 136.9000 54.2000 137.3000 54.3000 ;
	    RECT 140.6000 54.2000 140.9000 54.8000 ;
	    RECT 141.4000 54.6000 143.3000 54.9000 ;
	    RECT 141.4000 54.5000 141.8000 54.6000 ;
	    RECT 134.2000 53.8000 134.6000 54.2000 ;
	    RECT 135.4000 53.9000 140.9000 54.2000 ;
	    RECT 135.4000 53.8000 136.2000 53.9000 ;
	    RECT 128.6000 53.0000 130.6000 53.1000 ;
	    RECT 128.6000 51.1000 129.0000 53.0000 ;
	    RECT 130.2000 51.1000 130.6000 53.0000 ;
	    RECT 131.0000 51.1000 131.4000 53.1000 ;
	    RECT 133.4000 51.1000 133.8000 53.1000 ;
	    RECT 134.2000 52.8000 134.6000 53.2000 ;
	    RECT 134.1000 52.4000 134.5000 52.8000 ;
	    RECT 135.0000 51.1000 135.4000 53.5000 ;
	    RECT 137.5000 52.8000 137.8000 53.9000 ;
	    RECT 140.3000 53.8000 140.7000 53.9000 ;
	    RECT 143.8000 53.6000 144.2000 55.3000 ;
	    RECT 144.7000 54.2000 145.0000 55.8000 ;
	    RECT 147.0000 55.4000 147.4000 56.2000 ;
	    RECT 147.8000 55.4000 148.2000 56.2000 ;
	    RECT 150.2000 55.8000 150.6000 56.2000 ;
	    RECT 151.0000 55.9000 151.4000 59.9000 ;
	    RECT 152.6000 56.2000 153.0000 59.9000 ;
	    RECT 151.9000 55.9000 153.0000 56.2000 ;
	    RECT 153.4000 56.2000 153.8000 59.9000 ;
	    RECT 155.0000 56.2000 155.4000 59.9000 ;
	    RECT 153.4000 55.9000 155.4000 56.2000 ;
	    RECT 155.8000 55.9000 156.2000 59.9000 ;
	    RECT 157.9000 56.2000 158.3000 59.9000 ;
	    RECT 158.6000 56.8000 159.0000 57.2000 ;
	    RECT 158.7000 56.2000 159.0000 56.8000 ;
	    RECT 157.9000 55.9000 158.4000 56.2000 ;
	    RECT 158.7000 55.9000 159.4000 56.2000 ;
	    RECT 145.8000 54.8000 146.6000 55.2000 ;
	    RECT 148.6000 54.8000 149.4000 55.2000 ;
	    RECT 150.2000 54.2000 150.5000 55.8000 ;
	    RECT 144.7000 54.1000 145.5000 54.2000 ;
	    RECT 149.7000 54.1000 150.5000 54.2000 ;
	    RECT 144.7000 53.9000 145.6000 54.1000 ;
	    RECT 142.3000 53.3000 144.2000 53.6000 ;
	    RECT 142.3000 53.2000 142.7000 53.3000 ;
	    RECT 136.6000 52.1000 137.0000 52.5000 ;
	    RECT 137.4000 52.4000 137.8000 52.8000 ;
	    RECT 138.3000 52.7000 138.7000 52.8000 ;
	    RECT 138.3000 52.4000 139.7000 52.7000 ;
	    RECT 139.4000 52.1000 139.7000 52.4000 ;
	    RECT 141.4000 52.1000 141.8000 52.5000 ;
	    RECT 136.6000 51.8000 137.6000 52.1000 ;
	    RECT 137.2000 51.1000 137.6000 51.8000 ;
	    RECT 139.4000 51.1000 139.8000 52.1000 ;
	    RECT 141.4000 51.8000 142.1000 52.1000 ;
	    RECT 141.5000 51.1000 142.1000 51.8000 ;
	    RECT 143.8000 51.1000 144.2000 53.3000 ;
	    RECT 145.2000 51.1000 145.6000 53.9000 ;
	    RECT 149.6000 53.9000 150.5000 54.1000 ;
	    RECT 151.0000 54.8000 151.3000 55.9000 ;
	    RECT 151.9000 55.6000 152.2000 55.9000 ;
	    RECT 151.6000 55.2000 152.2000 55.6000 ;
	    RECT 153.8000 55.2000 154.2000 55.4000 ;
	    RECT 155.8000 55.2000 156.1000 55.9000 ;
	    RECT 149.6000 51.1000 150.0000 53.9000 ;
	    RECT 151.0000 51.1000 151.4000 54.8000 ;
	    RECT 151.9000 53.7000 152.2000 55.2000 ;
	    RECT 153.4000 54.9000 154.2000 55.2000 ;
	    RECT 155.0000 54.9000 156.2000 55.2000 ;
	    RECT 153.4000 54.8000 153.8000 54.9000 ;
	    RECT 154.2000 53.8000 154.6000 54.6000 ;
	    RECT 151.9000 53.4000 153.0000 53.7000 ;
	    RECT 152.6000 51.1000 153.0000 53.4000 ;
	    RECT 155.0000 53.1000 155.3000 54.9000 ;
	    RECT 155.8000 54.8000 156.2000 54.9000 ;
	    RECT 157.4000 54.4000 157.8000 55.2000 ;
	    RECT 158.1000 54.2000 158.4000 55.9000 ;
	    RECT 159.0000 55.8000 159.4000 55.9000 ;
	    RECT 161.4000 55.7000 161.8000 59.9000 ;
	    RECT 163.6000 58.2000 164.0000 59.9000 ;
	    RECT 163.0000 57.9000 164.0000 58.2000 ;
	    RECT 165.8000 57.9000 166.2000 59.9000 ;
	    RECT 167.9000 57.9000 168.5000 59.9000 ;
	    RECT 163.0000 57.5000 163.4000 57.9000 ;
	    RECT 165.8000 57.6000 166.1000 57.9000 ;
	    RECT 164.7000 57.3000 166.5000 57.6000 ;
	    RECT 167.8000 57.5000 168.2000 57.9000 ;
	    RECT 164.7000 57.2000 165.1000 57.3000 ;
	    RECT 166.1000 57.2000 166.5000 57.3000 ;
	    RECT 163.0000 56.5000 163.4000 56.6000 ;
	    RECT 165.3000 56.5000 165.7000 56.6000 ;
	    RECT 163.0000 56.2000 165.7000 56.5000 ;
	    RECT 166.0000 56.5000 167.1000 56.8000 ;
	    RECT 166.0000 55.9000 166.3000 56.5000 ;
	    RECT 166.7000 56.4000 167.1000 56.5000 ;
	    RECT 167.9000 56.6000 168.6000 57.0000 ;
	    RECT 167.9000 56.1000 168.2000 56.6000 ;
	    RECT 163.9000 55.7000 166.3000 55.9000 ;
	    RECT 161.4000 55.6000 166.3000 55.7000 ;
	    RECT 167.0000 55.8000 168.2000 56.1000 ;
	    RECT 161.4000 55.5000 164.3000 55.6000 ;
	    RECT 161.4000 55.4000 164.2000 55.5000 ;
	    RECT 164.6000 55.1000 165.0000 55.2000 ;
	    RECT 162.5000 54.8000 165.0000 55.1000 ;
	    RECT 162.5000 54.7000 162.9000 54.8000 ;
	    RECT 163.8000 54.7000 164.2000 54.8000 ;
	    RECT 163.3000 54.2000 163.7000 54.3000 ;
	    RECT 167.0000 54.2000 167.3000 55.8000 ;
	    RECT 170.2000 55.6000 170.6000 59.9000 ;
	    RECT 168.5000 55.3000 170.6000 55.6000 ;
	    RECT 168.5000 55.2000 168.9000 55.3000 ;
	    RECT 169.3000 54.9000 169.7000 55.0000 ;
	    RECT 167.8000 54.6000 169.7000 54.9000 ;
	    RECT 167.8000 54.5000 168.2000 54.6000 ;
	    RECT 158.1000 53.8000 159.4000 54.2000 ;
	    RECT 161.8000 53.9000 167.3000 54.2000 ;
	    RECT 161.8000 53.8000 162.6000 53.9000 ;
	    RECT 155.0000 51.1000 155.4000 53.1000 ;
	    RECT 155.8000 52.8000 156.2000 53.2000 ;
	    RECT 156.7000 53.1000 158.5000 53.3000 ;
	    RECT 159.0000 53.1000 159.3000 53.8000 ;
	    RECT 156.6000 53.0000 158.6000 53.1000 ;
	    RECT 155.7000 52.4000 156.1000 52.8000 ;
	    RECT 156.6000 51.1000 157.0000 53.0000 ;
	    RECT 158.2000 51.1000 158.6000 53.0000 ;
	    RECT 159.0000 51.1000 159.4000 53.1000 ;
	    RECT 161.4000 51.1000 161.8000 53.5000 ;
	    RECT 163.9000 52.8000 164.2000 53.9000 ;
	    RECT 166.7000 53.8000 167.1000 53.9000 ;
	    RECT 170.2000 53.6000 170.6000 55.3000 ;
	    RECT 168.7000 53.3000 170.6000 53.6000 ;
	    RECT 171.0000 53.4000 171.4000 54.2000 ;
	    RECT 171.8000 54.1000 172.2000 59.9000 ;
	    RECT 172.6000 55.8000 173.0000 56.6000 ;
	    RECT 173.4000 55.9000 173.8000 59.9000 ;
	    RECT 174.2000 56.2000 174.6000 59.9000 ;
	    RECT 175.8000 56.2000 176.2000 59.9000 ;
	    RECT 174.2000 55.9000 176.2000 56.2000 ;
	    RECT 173.5000 55.2000 173.8000 55.9000 ;
	    RECT 175.4000 55.2000 175.8000 55.4000 ;
	    RECT 173.4000 54.9000 174.6000 55.2000 ;
	    RECT 175.4000 54.9000 176.2000 55.2000 ;
	    RECT 173.4000 54.8000 173.8000 54.9000 ;
	    RECT 172.6000 54.1000 173.0000 54.2000 ;
	    RECT 171.8000 53.8000 173.0000 54.1000 ;
	    RECT 168.7000 53.2000 169.1000 53.3000 ;
	    RECT 163.0000 52.1000 163.4000 52.5000 ;
	    RECT 163.8000 52.4000 164.2000 52.8000 ;
	    RECT 164.7000 52.7000 165.1000 52.8000 ;
	    RECT 164.7000 52.4000 166.1000 52.7000 ;
	    RECT 165.8000 52.1000 166.1000 52.4000 ;
	    RECT 167.8000 52.1000 168.2000 52.5000 ;
	    RECT 163.0000 51.8000 164.0000 52.1000 ;
	    RECT 163.6000 51.1000 164.0000 51.8000 ;
	    RECT 165.8000 51.1000 166.2000 52.1000 ;
	    RECT 167.8000 51.8000 168.5000 52.1000 ;
	    RECT 167.9000 51.1000 168.5000 51.8000 ;
	    RECT 170.2000 51.1000 170.6000 53.3000 ;
	    RECT 171.8000 53.1000 172.2000 53.8000 ;
	    RECT 171.8000 52.8000 172.7000 53.1000 ;
	    RECT 173.4000 52.8000 173.8000 53.2000 ;
	    RECT 174.3000 53.1000 174.6000 54.9000 ;
	    RECT 175.8000 54.8000 176.2000 54.9000 ;
	    RECT 175.0000 53.8000 175.4000 54.6000 ;
	    RECT 172.3000 51.1000 172.7000 52.8000 ;
	    RECT 173.5000 52.4000 173.9000 52.8000 ;
	    RECT 174.2000 51.1000 174.6000 53.1000 ;
	    RECT 176.6000 52.4000 177.0000 53.2000 ;
	    RECT 177.4000 51.1000 177.8000 59.9000 ;
	    RECT 178.2000 53.4000 178.6000 54.2000 ;
	    RECT 179.0000 54.1000 179.4000 59.9000 ;
	    RECT 179.8000 55.8000 180.2000 56.6000 ;
	    RECT 180.6000 55.9000 181.0000 59.9000 ;
	    RECT 181.4000 56.2000 181.8000 59.9000 ;
	    RECT 183.0000 56.2000 183.4000 59.9000 ;
	    RECT 181.4000 55.9000 183.4000 56.2000 ;
	    RECT 180.7000 55.2000 181.0000 55.9000 ;
	    RECT 183.8000 55.7000 184.2000 59.9000 ;
	    RECT 186.0000 58.2000 186.4000 59.9000 ;
	    RECT 185.4000 57.9000 186.4000 58.2000 ;
	    RECT 188.2000 57.9000 188.6000 59.9000 ;
	    RECT 190.3000 57.9000 190.9000 59.9000 ;
	    RECT 185.4000 57.5000 185.8000 57.9000 ;
	    RECT 188.2000 57.6000 188.5000 57.9000 ;
	    RECT 187.1000 57.3000 188.9000 57.6000 ;
	    RECT 190.2000 57.5000 190.6000 57.9000 ;
	    RECT 187.1000 57.2000 187.5000 57.3000 ;
	    RECT 188.5000 57.2000 188.9000 57.3000 ;
	    RECT 185.4000 56.5000 185.8000 56.6000 ;
	    RECT 187.7000 56.5000 188.1000 56.6000 ;
	    RECT 185.4000 56.2000 188.1000 56.5000 ;
	    RECT 188.4000 56.5000 189.5000 56.8000 ;
	    RECT 188.4000 55.9000 188.7000 56.5000 ;
	    RECT 189.1000 56.4000 189.5000 56.5000 ;
	    RECT 190.3000 56.6000 191.0000 57.0000 ;
	    RECT 190.3000 56.1000 190.6000 56.6000 ;
	    RECT 186.3000 55.7000 188.7000 55.9000 ;
	    RECT 183.8000 55.6000 188.7000 55.7000 ;
	    RECT 189.4000 55.8000 190.6000 56.1000 ;
	    RECT 183.8000 55.5000 186.7000 55.6000 ;
	    RECT 183.8000 55.4000 186.6000 55.5000 ;
	    RECT 182.6000 55.2000 183.0000 55.4000 ;
	    RECT 189.4000 55.2000 189.7000 55.8000 ;
	    RECT 192.6000 55.6000 193.0000 59.9000 ;
	    RECT 190.9000 55.3000 193.0000 55.6000 ;
	    RECT 190.9000 55.2000 191.3000 55.3000 ;
	    RECT 180.6000 54.9000 181.8000 55.2000 ;
	    RECT 182.6000 54.9000 183.4000 55.2000 ;
	    RECT 187.0000 55.1000 187.4000 55.2000 ;
	    RECT 180.6000 54.8000 181.0000 54.9000 ;
	    RECT 179.8000 54.1000 180.2000 54.2000 ;
	    RECT 179.0000 53.8000 180.2000 54.1000 ;
	    RECT 179.0000 53.1000 179.4000 53.8000 ;
	    RECT 179.0000 52.8000 179.9000 53.1000 ;
	    RECT 180.6000 52.8000 181.0000 53.2000 ;
	    RECT 181.5000 53.1000 181.8000 54.9000 ;
	    RECT 183.0000 54.8000 183.4000 54.9000 ;
	    RECT 184.9000 54.8000 187.4000 55.1000 ;
	    RECT 189.4000 54.8000 189.8000 55.2000 ;
	    RECT 191.7000 54.9000 192.1000 55.0000 ;
	    RECT 184.9000 54.7000 185.3000 54.8000 ;
	    RECT 186.2000 54.7000 186.6000 54.8000 ;
	    RECT 182.2000 53.8000 182.6000 54.6000 ;
	    RECT 185.7000 54.2000 186.1000 54.3000 ;
	    RECT 189.4000 54.2000 189.7000 54.8000 ;
	    RECT 190.2000 54.6000 192.1000 54.9000 ;
	    RECT 190.2000 54.5000 190.6000 54.6000 ;
	    RECT 183.0000 54.1000 183.4000 54.2000 ;
	    RECT 184.2000 54.1000 189.7000 54.2000 ;
	    RECT 183.0000 53.9000 189.7000 54.1000 ;
	    RECT 183.0000 53.8000 185.0000 53.9000 ;
	    RECT 179.5000 51.1000 179.9000 52.8000 ;
	    RECT 180.7000 52.4000 181.1000 52.8000 ;
	    RECT 181.4000 51.1000 181.8000 53.1000 ;
	    RECT 183.8000 51.1000 184.2000 53.5000 ;
	    RECT 186.3000 52.8000 186.6000 53.9000 ;
	    RECT 189.1000 53.8000 189.5000 53.9000 ;
	    RECT 192.6000 53.6000 193.0000 55.3000 ;
	    RECT 191.1000 53.3000 193.0000 53.6000 ;
	    RECT 191.1000 53.2000 191.5000 53.3000 ;
	    RECT 185.4000 52.1000 185.8000 52.5000 ;
	    RECT 186.2000 52.4000 186.6000 52.8000 ;
	    RECT 187.1000 52.7000 187.5000 52.8000 ;
	    RECT 187.1000 52.4000 188.5000 52.7000 ;
	    RECT 188.2000 52.1000 188.5000 52.4000 ;
	    RECT 190.2000 52.1000 190.6000 52.5000 ;
	    RECT 185.4000 51.8000 186.4000 52.1000 ;
	    RECT 186.0000 51.1000 186.4000 51.8000 ;
	    RECT 188.2000 51.1000 188.6000 52.1000 ;
	    RECT 190.2000 51.8000 190.9000 52.1000 ;
	    RECT 190.3000 51.1000 190.9000 51.8000 ;
	    RECT 192.6000 51.1000 193.0000 53.3000 ;
	    RECT 193.4000 51.1000 193.8000 59.9000 ;
	    RECT 195.0000 55.6000 195.4000 59.9000 ;
	    RECT 197.1000 57.9000 197.7000 59.9000 ;
	    RECT 199.4000 57.9000 199.8000 59.9000 ;
	    RECT 201.6000 58.2000 202.0000 59.9000 ;
	    RECT 201.6000 57.9000 202.6000 58.2000 ;
	    RECT 197.4000 57.5000 197.8000 57.9000 ;
	    RECT 199.5000 57.6000 199.8000 57.9000 ;
	    RECT 199.1000 57.3000 200.9000 57.6000 ;
	    RECT 202.2000 57.5000 202.6000 57.9000 ;
	    RECT 199.1000 57.2000 199.5000 57.3000 ;
	    RECT 200.5000 57.2000 200.9000 57.3000 ;
	    RECT 197.0000 56.6000 197.7000 57.0000 ;
	    RECT 197.4000 56.1000 197.7000 56.6000 ;
	    RECT 198.5000 56.5000 199.6000 56.8000 ;
	    RECT 198.5000 56.4000 198.9000 56.5000 ;
	    RECT 197.4000 55.8000 198.6000 56.1000 ;
	    RECT 195.0000 55.3000 197.1000 55.6000 ;
	    RECT 195.0000 53.6000 195.4000 55.3000 ;
	    RECT 196.7000 55.2000 197.1000 55.3000 ;
	    RECT 198.3000 55.2000 198.6000 55.8000 ;
	    RECT 199.3000 55.9000 199.6000 56.5000 ;
	    RECT 199.9000 56.5000 200.3000 56.6000 ;
	    RECT 202.2000 56.5000 202.6000 56.6000 ;
	    RECT 199.9000 56.2000 202.6000 56.5000 ;
	    RECT 199.3000 55.7000 201.7000 55.9000 ;
	    RECT 203.8000 55.7000 204.2000 59.9000 ;
	    RECT 204.6000 55.9000 205.0000 59.9000 ;
	    RECT 205.4000 56.2000 205.8000 59.9000 ;
	    RECT 207.0000 56.2000 207.4000 59.9000 ;
	    RECT 205.4000 55.9000 207.4000 56.2000 ;
	    RECT 199.3000 55.6000 204.2000 55.7000 ;
	    RECT 201.3000 55.5000 204.2000 55.6000 ;
	    RECT 201.4000 55.4000 204.2000 55.5000 ;
	    RECT 204.7000 55.2000 205.0000 55.9000 ;
	    RECT 209.4000 55.7000 209.8000 59.9000 ;
	    RECT 211.6000 58.2000 212.0000 59.9000 ;
	    RECT 211.0000 57.9000 212.0000 58.2000 ;
	    RECT 213.8000 57.9000 214.2000 59.9000 ;
	    RECT 215.9000 57.9000 216.5000 59.9000 ;
	    RECT 211.0000 57.5000 211.4000 57.9000 ;
	    RECT 213.8000 57.6000 214.1000 57.9000 ;
	    RECT 212.7000 57.3000 214.5000 57.6000 ;
	    RECT 215.8000 57.5000 216.2000 57.9000 ;
	    RECT 212.7000 57.2000 213.1000 57.3000 ;
	    RECT 214.1000 57.2000 214.5000 57.3000 ;
	    RECT 211.0000 56.5000 211.4000 56.6000 ;
	    RECT 213.3000 56.5000 213.7000 56.6000 ;
	    RECT 211.0000 56.2000 213.7000 56.5000 ;
	    RECT 214.0000 56.5000 215.1000 56.8000 ;
	    RECT 214.0000 55.9000 214.3000 56.5000 ;
	    RECT 214.7000 56.4000 215.1000 56.5000 ;
	    RECT 215.9000 56.6000 216.6000 57.0000 ;
	    RECT 215.9000 56.1000 216.2000 56.6000 ;
	    RECT 211.9000 55.7000 214.3000 55.9000 ;
	    RECT 209.4000 55.6000 214.3000 55.7000 ;
	    RECT 215.0000 55.8000 216.2000 56.1000 ;
	    RECT 209.4000 55.5000 212.3000 55.6000 ;
	    RECT 209.4000 55.4000 212.2000 55.5000 ;
	    RECT 206.6000 55.2000 207.0000 55.4000 ;
	    RECT 195.9000 54.9000 196.3000 55.0000 ;
	    RECT 195.9000 54.6000 197.8000 54.9000 ;
	    RECT 198.2000 54.8000 198.6000 55.2000 ;
	    RECT 204.6000 54.9000 205.8000 55.2000 ;
	    RECT 206.6000 54.9000 207.4000 55.2000 ;
	    RECT 212.6000 55.1000 213.0000 55.2000 ;
	    RECT 204.6000 54.8000 205.0000 54.9000 ;
	    RECT 197.4000 54.5000 197.8000 54.6000 ;
	    RECT 198.3000 54.2000 198.6000 54.8000 ;
	    RECT 201.9000 54.2000 202.3000 54.3000 ;
	    RECT 198.3000 54.1000 203.8000 54.2000 ;
	    RECT 204.6000 54.1000 205.0000 54.2000 ;
	    RECT 198.3000 53.9000 205.0000 54.1000 ;
	    RECT 198.5000 53.8000 198.9000 53.9000 ;
	    RECT 195.0000 53.3000 196.9000 53.6000 ;
	    RECT 194.2000 53.1000 194.6000 53.2000 ;
	    RECT 195.0000 53.1000 195.4000 53.3000 ;
	    RECT 196.5000 53.2000 196.9000 53.3000 ;
	    RECT 194.2000 52.8000 195.4000 53.1000 ;
	    RECT 201.4000 52.8000 201.7000 53.9000 ;
	    RECT 203.0000 53.8000 205.0000 53.9000 ;
	    RECT 194.2000 52.4000 194.6000 52.8000 ;
	    RECT 195.0000 51.1000 195.4000 52.8000 ;
	    RECT 200.5000 52.7000 200.9000 52.8000 ;
	    RECT 197.4000 52.1000 197.8000 52.5000 ;
	    RECT 199.5000 52.4000 200.9000 52.7000 ;
	    RECT 201.4000 52.4000 201.8000 52.8000 ;
	    RECT 199.5000 52.1000 199.8000 52.4000 ;
	    RECT 202.2000 52.1000 202.6000 52.5000 ;
	    RECT 197.1000 51.8000 197.8000 52.1000 ;
	    RECT 197.1000 51.1000 197.7000 51.8000 ;
	    RECT 199.4000 51.1000 199.8000 52.1000 ;
	    RECT 201.6000 51.8000 202.6000 52.1000 ;
	    RECT 201.6000 51.1000 202.0000 51.8000 ;
	    RECT 203.8000 51.1000 204.2000 53.5000 ;
	    RECT 205.5000 53.2000 205.8000 54.9000 ;
	    RECT 207.0000 54.8000 207.4000 54.9000 ;
	    RECT 210.5000 54.8000 213.0000 55.1000 ;
	    RECT 210.5000 54.7000 210.9000 54.8000 ;
	    RECT 211.8000 54.7000 212.2000 54.8000 ;
	    RECT 206.2000 53.8000 206.6000 54.6000 ;
	    RECT 211.3000 54.2000 211.7000 54.3000 ;
	    RECT 215.0000 54.2000 215.3000 55.8000 ;
	    RECT 218.2000 55.6000 218.6000 59.9000 ;
	    RECT 216.5000 55.3000 218.6000 55.6000 ;
	    RECT 219.0000 55.7000 219.4000 59.9000 ;
	    RECT 221.2000 58.2000 221.6000 59.9000 ;
	    RECT 220.6000 57.9000 221.6000 58.2000 ;
	    RECT 223.4000 57.9000 223.8000 59.9000 ;
	    RECT 225.5000 57.9000 226.1000 59.9000 ;
	    RECT 220.6000 57.5000 221.0000 57.9000 ;
	    RECT 223.4000 57.6000 223.7000 57.9000 ;
	    RECT 222.3000 57.3000 224.1000 57.6000 ;
	    RECT 225.4000 57.5000 225.8000 57.9000 ;
	    RECT 222.3000 57.2000 222.7000 57.3000 ;
	    RECT 223.7000 57.2000 224.1000 57.3000 ;
	    RECT 220.6000 56.5000 221.0000 56.6000 ;
	    RECT 222.9000 56.5000 223.3000 56.6000 ;
	    RECT 220.6000 56.2000 223.3000 56.5000 ;
	    RECT 223.6000 56.5000 224.7000 56.8000 ;
	    RECT 223.6000 55.9000 223.9000 56.5000 ;
	    RECT 224.3000 56.4000 224.7000 56.5000 ;
	    RECT 225.5000 56.6000 226.2000 57.0000 ;
	    RECT 225.5000 56.1000 225.8000 56.6000 ;
	    RECT 221.5000 55.7000 223.9000 55.9000 ;
	    RECT 219.0000 55.6000 223.9000 55.7000 ;
	    RECT 224.6000 55.8000 225.8000 56.1000 ;
	    RECT 219.0000 55.5000 221.9000 55.6000 ;
	    RECT 219.0000 55.4000 221.8000 55.5000 ;
	    RECT 216.5000 55.2000 216.9000 55.3000 ;
	    RECT 217.3000 54.9000 217.7000 55.0000 ;
	    RECT 215.8000 54.6000 217.7000 54.9000 ;
	    RECT 215.8000 54.5000 216.2000 54.6000 ;
	    RECT 209.8000 53.9000 215.3000 54.2000 ;
	    RECT 209.8000 53.8000 210.6000 53.9000 ;
	    RECT 204.6000 52.8000 205.0000 53.2000 ;
	    RECT 204.7000 52.4000 205.1000 52.8000 ;
	    RECT 205.4000 51.1000 205.8000 53.2000 ;
	    RECT 209.4000 51.1000 209.8000 53.5000 ;
	    RECT 211.9000 52.8000 212.2000 53.9000 ;
	    RECT 214.7000 53.8000 215.1000 53.9000 ;
	    RECT 218.2000 53.6000 218.6000 55.3000 ;
	    RECT 222.2000 55.1000 222.6000 55.2000 ;
	    RECT 220.1000 54.8000 222.6000 55.1000 ;
	    RECT 220.1000 54.7000 220.5000 54.8000 ;
	    RECT 221.4000 54.7000 221.8000 54.8000 ;
	    RECT 220.9000 54.2000 221.3000 54.3000 ;
	    RECT 224.6000 54.2000 224.9000 55.8000 ;
	    RECT 227.8000 55.6000 228.2000 59.9000 ;
	    RECT 228.9000 59.2000 229.3000 59.9000 ;
	    RECT 228.9000 58.8000 229.8000 59.2000 ;
	    RECT 228.9000 56.3000 229.3000 58.8000 ;
	    RECT 231.8000 57.9000 232.2000 59.9000 ;
	    RECT 228.9000 55.9000 229.8000 56.3000 ;
	    RECT 226.1000 55.3000 228.2000 55.6000 ;
	    RECT 226.1000 55.2000 226.5000 55.3000 ;
	    RECT 226.9000 54.9000 227.3000 55.0000 ;
	    RECT 225.4000 54.6000 227.3000 54.9000 ;
	    RECT 225.4000 54.5000 225.8000 54.6000 ;
	    RECT 219.4000 53.9000 224.9000 54.2000 ;
	    RECT 219.4000 53.8000 220.2000 53.9000 ;
	    RECT 216.7000 53.3000 218.6000 53.6000 ;
	    RECT 216.7000 53.2000 217.1000 53.3000 ;
	    RECT 211.0000 52.1000 211.4000 52.5000 ;
	    RECT 211.8000 52.4000 212.2000 52.8000 ;
	    RECT 212.7000 52.7000 213.1000 52.8000 ;
	    RECT 212.7000 52.4000 214.1000 52.7000 ;
	    RECT 213.8000 52.1000 214.1000 52.4000 ;
	    RECT 215.8000 52.1000 216.2000 52.5000 ;
	    RECT 211.0000 51.8000 212.0000 52.1000 ;
	    RECT 211.6000 51.1000 212.0000 51.8000 ;
	    RECT 213.8000 51.1000 214.2000 52.1000 ;
	    RECT 215.8000 51.8000 216.5000 52.1000 ;
	    RECT 215.9000 51.1000 216.5000 51.8000 ;
	    RECT 218.2000 51.1000 218.6000 53.3000 ;
	    RECT 219.0000 51.1000 219.4000 53.5000 ;
	    RECT 221.5000 52.8000 221.8000 53.9000 ;
	    RECT 222.2000 53.8000 222.6000 53.9000 ;
	    RECT 224.3000 53.8000 224.7000 53.9000 ;
	    RECT 227.8000 53.6000 228.2000 55.3000 ;
	    RECT 228.6000 54.8000 229.0000 55.6000 ;
	    RECT 228.6000 54.2000 228.9000 54.8000 ;
	    RECT 229.4000 54.2000 229.7000 55.9000 ;
	    RECT 231.9000 55.8000 232.2000 57.9000 ;
	    RECT 233.4000 55.9000 233.8000 59.9000 ;
	    RECT 231.9000 55.5000 233.1000 55.8000 ;
	    RECT 231.8000 54.8000 232.2000 55.2000 ;
	    RECT 228.6000 53.8000 229.0000 54.2000 ;
	    RECT 229.4000 53.8000 229.8000 54.2000 ;
	    RECT 231.0000 54.1000 231.4000 54.6000 ;
	    RECT 231.9000 54.4000 232.2000 54.8000 ;
	    RECT 231.9000 54.1000 232.4000 54.4000 ;
	    RECT 230.2000 53.8000 231.4000 54.1000 ;
	    RECT 232.0000 54.0000 232.4000 54.1000 ;
	    RECT 232.8000 53.8000 233.1000 55.5000 ;
	    RECT 233.5000 55.2000 233.8000 55.9000 ;
	    RECT 233.4000 54.8000 233.8000 55.2000 ;
	    RECT 226.3000 53.3000 228.2000 53.6000 ;
	    RECT 226.3000 53.2000 226.7000 53.3000 ;
	    RECT 220.6000 52.1000 221.0000 52.5000 ;
	    RECT 221.4000 52.4000 221.8000 52.8000 ;
	    RECT 222.3000 52.7000 222.7000 52.8000 ;
	    RECT 222.3000 52.4000 223.7000 52.7000 ;
	    RECT 223.4000 52.1000 223.7000 52.4000 ;
	    RECT 225.4000 52.1000 225.8000 52.5000 ;
	    RECT 220.6000 51.8000 221.6000 52.1000 ;
	    RECT 221.2000 51.1000 221.6000 51.8000 ;
	    RECT 223.4000 51.1000 223.8000 52.1000 ;
	    RECT 225.4000 51.8000 226.1000 52.1000 ;
	    RECT 225.5000 51.1000 226.1000 51.8000 ;
	    RECT 227.8000 51.1000 228.2000 53.3000 ;
	    RECT 229.4000 52.1000 229.7000 53.8000 ;
	    RECT 230.2000 53.2000 230.5000 53.8000 ;
	    RECT 232.8000 53.7000 233.2000 53.8000 ;
	    RECT 231.7000 53.5000 233.2000 53.7000 ;
	    RECT 231.1000 53.4000 233.2000 53.5000 ;
	    RECT 231.1000 53.2000 232.0000 53.4000 ;
	    RECT 230.2000 52.4000 230.6000 53.2000 ;
	    RECT 231.1000 53.1000 231.4000 53.2000 ;
	    RECT 233.5000 53.1000 233.8000 54.8000 ;
	    RECT 229.4000 51.1000 229.8000 52.1000 ;
	    RECT 231.0000 51.1000 231.4000 53.1000 ;
	    RECT 233.1000 52.6000 233.8000 53.1000 ;
	    RECT 234.2000 55.6000 234.6000 59.9000 ;
	    RECT 236.3000 57.9000 236.9000 59.9000 ;
	    RECT 238.6000 57.9000 239.0000 59.9000 ;
	    RECT 240.8000 58.2000 241.2000 59.9000 ;
	    RECT 240.8000 57.9000 241.8000 58.2000 ;
	    RECT 236.6000 57.5000 237.0000 57.9000 ;
	    RECT 238.7000 57.6000 239.0000 57.9000 ;
	    RECT 238.3000 57.3000 240.1000 57.6000 ;
	    RECT 241.4000 57.5000 241.8000 57.9000 ;
	    RECT 238.3000 57.2000 238.7000 57.3000 ;
	    RECT 239.7000 57.2000 240.1000 57.3000 ;
	    RECT 236.2000 56.6000 236.9000 57.0000 ;
	    RECT 236.6000 56.1000 236.9000 56.6000 ;
	    RECT 237.7000 56.5000 238.8000 56.8000 ;
	    RECT 237.7000 56.4000 238.1000 56.5000 ;
	    RECT 236.6000 55.8000 237.8000 56.1000 ;
	    RECT 234.2000 55.3000 236.3000 55.6000 ;
	    RECT 234.2000 53.6000 234.6000 55.3000 ;
	    RECT 235.9000 55.2000 236.3000 55.3000 ;
	    RECT 235.1000 54.9000 235.5000 55.0000 ;
	    RECT 235.1000 54.6000 237.0000 54.9000 ;
	    RECT 236.6000 54.5000 237.0000 54.6000 ;
	    RECT 237.5000 54.2000 237.8000 55.8000 ;
	    RECT 238.5000 55.9000 238.8000 56.5000 ;
	    RECT 239.1000 56.5000 239.5000 56.6000 ;
	    RECT 241.4000 56.5000 241.8000 56.6000 ;
	    RECT 239.1000 56.2000 241.8000 56.5000 ;
	    RECT 238.5000 55.7000 240.9000 55.9000 ;
	    RECT 243.0000 55.7000 243.4000 59.9000 ;
	    RECT 238.5000 55.6000 243.4000 55.7000 ;
	    RECT 240.5000 55.5000 243.4000 55.6000 ;
	    RECT 240.6000 55.4000 243.4000 55.5000 ;
	    RECT 244.6000 56.1000 245.0000 59.9000 ;
	    RECT 246.2000 57.9000 246.6000 59.9000 ;
	    RECT 245.4000 56.1000 245.8000 56.2000 ;
	    RECT 244.6000 55.8000 245.8000 56.1000 ;
	    RECT 246.3000 55.8000 246.6000 57.9000 ;
	    RECT 247.8000 55.9000 248.2000 59.9000 ;
	    RECT 248.6000 56.9000 249.0000 59.9000 ;
	    RECT 248.7000 56.6000 249.0000 56.9000 ;
	    RECT 250.2000 59.6000 252.2000 59.9000 ;
	    RECT 250.2000 56.9000 250.6000 59.6000 ;
	    RECT 251.0000 56.9000 251.4000 59.3000 ;
	    RECT 251.8000 57.0000 252.2000 59.6000 ;
	    RECT 252.7000 59.6000 254.5000 59.9000 ;
	    RECT 252.7000 59.5000 253.0000 59.6000 ;
	    RECT 250.2000 56.6000 250.5000 56.9000 ;
	    RECT 248.7000 56.3000 250.5000 56.6000 ;
	    RECT 251.1000 56.7000 251.4000 56.9000 ;
	    RECT 252.6000 56.7000 253.0000 59.5000 ;
	    RECT 254.2000 59.5000 254.5000 59.6000 ;
	    RECT 251.1000 56.5000 253.0000 56.7000 ;
	    RECT 253.4000 56.5000 253.8000 59.3000 ;
	    RECT 254.2000 56.5000 254.6000 59.5000 ;
	    RECT 251.1000 56.4000 252.9000 56.5000 ;
	    RECT 253.4000 56.2000 253.7000 56.5000 ;
	    RECT 255.3000 56.3000 255.7000 59.9000 ;
	    RECT 253.4000 56.1000 253.8000 56.2000 ;
	    RECT 239.8000 55.1000 240.2000 55.2000 ;
	    RECT 239.8000 54.8000 242.3000 55.1000 ;
	    RECT 240.6000 54.7000 241.0000 54.8000 ;
	    RECT 241.9000 54.7000 242.3000 54.8000 ;
	    RECT 241.1000 54.2000 241.5000 54.3000 ;
	    RECT 237.5000 53.9000 243.0000 54.2000 ;
	    RECT 237.7000 53.8000 238.1000 53.9000 ;
	    RECT 234.2000 53.3000 236.1000 53.6000 ;
	    RECT 233.1000 51.1000 233.5000 52.6000 ;
	    RECT 234.2000 51.1000 234.6000 53.3000 ;
	    RECT 235.7000 53.2000 236.1000 53.3000 ;
	    RECT 240.6000 52.8000 240.9000 53.9000 ;
	    RECT 242.2000 53.8000 243.0000 53.9000 ;
	    RECT 239.7000 52.7000 240.1000 52.8000 ;
	    RECT 236.6000 52.1000 237.0000 52.5000 ;
	    RECT 238.7000 52.4000 240.1000 52.7000 ;
	    RECT 240.6000 52.4000 241.0000 52.8000 ;
	    RECT 238.7000 52.1000 239.0000 52.4000 ;
	    RECT 241.4000 52.1000 241.8000 52.5000 ;
	    RECT 236.3000 51.8000 237.0000 52.1000 ;
	    RECT 236.3000 51.1000 236.9000 51.8000 ;
	    RECT 238.6000 51.1000 239.0000 52.1000 ;
	    RECT 240.8000 51.8000 241.8000 52.1000 ;
	    RECT 240.8000 51.1000 241.2000 51.8000 ;
	    RECT 243.0000 51.1000 243.4000 53.5000 ;
	    RECT 243.8000 52.4000 244.2000 53.2000 ;
	    RECT 244.6000 51.1000 245.0000 55.8000 ;
	    RECT 246.3000 55.5000 247.5000 55.8000 ;
	    RECT 246.2000 54.8000 246.6000 55.2000 ;
	    RECT 245.4000 53.8000 245.8000 54.6000 ;
	    RECT 246.3000 54.4000 246.6000 54.8000 ;
	    RECT 246.3000 54.1000 246.8000 54.4000 ;
	    RECT 246.4000 54.0000 246.8000 54.1000 ;
	    RECT 247.2000 53.8000 247.5000 55.5000 ;
	    RECT 247.9000 55.2000 248.2000 55.9000 ;
	    RECT 252.1000 55.8000 253.8000 56.1000 ;
	    RECT 255.3000 55.9000 256.2000 56.3000 ;
	    RECT 257.4000 55.9000 257.8000 59.9000 ;
	    RECT 258.2000 56.2000 258.6000 59.9000 ;
	    RECT 259.8000 56.2000 260.2000 59.9000 ;
	    RECT 261.9000 56.2000 262.3000 59.9000 ;
	    RECT 258.2000 55.9000 260.2000 56.2000 ;
	    RECT 247.8000 55.1000 248.2000 55.2000 ;
	    RECT 251.0000 55.1000 251.8000 55.2000 ;
	    RECT 247.8000 54.8000 251.8000 55.1000 ;
	    RECT 247.2000 53.7000 247.6000 53.8000 ;
	    RECT 246.1000 53.5000 247.6000 53.7000 ;
	    RECT 245.5000 53.4000 247.6000 53.5000 ;
	    RECT 245.5000 53.2000 246.4000 53.4000 ;
	    RECT 245.5000 53.1000 245.8000 53.2000 ;
	    RECT 247.9000 53.1000 248.2000 54.8000 ;
	    RECT 249.4000 54.1000 249.8000 54.2000 ;
	    RECT 250.2000 54.1000 251.0000 54.2000 ;
	    RECT 249.4000 53.8000 251.0000 54.1000 ;
	    RECT 245.4000 51.1000 245.8000 53.1000 ;
	    RECT 247.5000 52.6000 248.2000 53.1000 ;
	    RECT 249.4000 52.8000 250.6000 53.2000 ;
	    RECT 247.5000 51.1000 247.9000 52.6000 ;
	    RECT 252.1000 52.5000 252.4000 55.8000 ;
	    RECT 255.0000 54.8000 255.4000 55.6000 ;
	    RECT 250.4000 52.2000 252.4000 52.5000 ;
	    RECT 250.2000 51.8000 250.7000 52.2000 ;
	    RECT 251.8000 52.1000 252.4000 52.2000 ;
	    RECT 255.8000 54.2000 256.1000 55.9000 ;
	    RECT 257.5000 55.2000 257.8000 55.9000 ;
	    RECT 261.4000 55.8000 262.4000 56.2000 ;
	    RECT 259.4000 55.2000 259.8000 55.4000 ;
	    RECT 257.4000 54.9000 258.6000 55.2000 ;
	    RECT 259.4000 54.9000 260.2000 55.2000 ;
	    RECT 257.4000 54.8000 257.8000 54.9000 ;
	    RECT 255.8000 53.8000 256.2000 54.2000 ;
	    RECT 255.8000 52.2000 256.1000 53.8000 ;
	    RECT 258.3000 53.2000 258.6000 54.9000 ;
	    RECT 259.8000 54.8000 260.2000 54.9000 ;
	    RECT 259.0000 53.8000 259.4000 54.6000 ;
	    RECT 262.1000 54.2000 262.4000 55.8000 ;
	    RECT 260.6000 54.1000 261.0000 54.2000 ;
	    RECT 260.6000 53.8000 261.4000 54.1000 ;
	    RECT 262.1000 53.8000 263.4000 54.2000 ;
	    RECT 264.6000 54.1000 265.0000 59.9000 ;
	    RECT 265.4000 54.1000 265.8000 54.2000 ;
	    RECT 264.6000 53.8000 265.8000 54.1000 ;
	    RECT 261.0000 53.6000 261.4000 53.8000 ;
	    RECT 256.6000 52.4000 257.0000 53.2000 ;
	    RECT 257.4000 52.8000 257.8000 53.2000 ;
	    RECT 257.5000 52.4000 257.9000 52.8000 ;
	    RECT 250.2000 51.1000 250.6000 51.8000 ;
	    RECT 251.8000 51.1000 252.2000 52.1000 ;
	    RECT 255.8000 51.1000 256.2000 52.2000 ;
	    RECT 258.2000 51.1000 258.6000 53.2000 ;
	    RECT 260.7000 53.1000 262.5000 53.3000 ;
	    RECT 263.0000 53.1000 263.3000 53.8000 ;
	    RECT 260.6000 53.0000 262.6000 53.1000 ;
	    RECT 260.6000 51.1000 261.0000 53.0000 ;
	    RECT 262.2000 51.1000 262.6000 53.0000 ;
	    RECT 263.0000 51.1000 263.4000 53.1000 ;
	    RECT 264.6000 51.1000 265.0000 53.8000 ;
	    RECT 265.4000 53.4000 265.8000 53.8000 ;
	    RECT 266.2000 54.1000 266.6000 59.9000 ;
	    RECT 267.0000 55.8000 267.4000 56.6000 ;
	    RECT 269.1000 56.3000 269.5000 59.9000 ;
	    RECT 268.6000 55.9000 269.5000 56.3000 ;
	    RECT 267.0000 55.1000 267.3000 55.8000 ;
	    RECT 268.7000 55.1000 269.0000 55.9000 ;
	    RECT 267.0000 54.8000 269.0000 55.1000 ;
	    RECT 268.7000 54.2000 269.0000 54.8000 ;
	    RECT 267.0000 54.1000 267.4000 54.2000 ;
	    RECT 266.2000 53.8000 267.4000 54.1000 ;
	    RECT 268.6000 53.8000 269.0000 54.2000 ;
	    RECT 266.2000 53.1000 266.6000 53.8000 ;
	    RECT 266.2000 52.8000 267.1000 53.1000 ;
	    RECT 266.7000 51.1000 267.1000 52.8000 ;
	    RECT 267.8000 52.4000 268.2000 53.2000 ;
	    RECT 268.7000 52.1000 269.0000 53.8000 ;
	    RECT 268.6000 51.1000 269.0000 52.1000 ;
	    RECT 0.6000 47.9000 1.0000 49.9000 ;
	    RECT 2.8000 49.2000 3.6000 49.9000 ;
	    RECT 2.8000 48.8000 4.2000 49.2000 ;
	    RECT 2.8000 48.1000 3.6000 48.8000 ;
	    RECT 0.6000 47.6000 1.8000 47.9000 ;
	    RECT 1.4000 47.5000 1.8000 47.6000 ;
	    RECT 2.1000 47.4000 2.5000 47.8000 ;
	    RECT 2.1000 47.2000 2.4000 47.4000 ;
	    RECT 2.0000 46.8000 2.4000 47.2000 ;
	    RECT 2.8000 47.1000 3.1000 48.1000 ;
	    RECT 5.4000 47.9000 5.8000 49.9000 ;
	    RECT 7.5000 48.2000 7.9000 49.9000 ;
	    RECT 8.7000 48.2000 9.1000 48.6000 ;
	    RECT 3.4000 47.4000 4.2000 47.8000 ;
	    RECT 4.5000 47.6000 5.8000 47.9000 ;
	    RECT 7.0000 47.9000 7.9000 48.2000 ;
	    RECT 4.5000 47.5000 4.9000 47.6000 ;
	    RECT 2.8000 46.8000 3.3000 47.1000 ;
	    RECT 3.0000 46.2000 3.3000 46.8000 ;
	    RECT 3.0000 45.8000 3.4000 46.2000 ;
	    RECT 4.3000 46.1000 4.7000 46.2000 ;
	    RECT 3.9000 45.8000 4.7000 46.1000 ;
	    RECT 6.2000 46.1000 6.6000 46.2000 ;
	    RECT 7.0000 46.1000 7.4000 47.9000 ;
	    RECT 8.6000 47.8000 9.0000 48.2000 ;
	    RECT 9.4000 47.9000 9.8000 49.9000 ;
	    RECT 9.5000 46.2000 9.8000 47.9000 ;
	    RECT 10.2000 46.4000 10.6000 47.2000 ;
	    RECT 6.2000 45.8000 7.4000 46.1000 ;
	    RECT 8.6000 46.1000 9.0000 46.2000 ;
	    RECT 9.4000 46.1000 9.8000 46.2000 ;
	    RECT 11.0000 46.1000 11.4000 46.2000 ;
	    RECT 11.8000 46.1000 12.2000 49.9000 ;
	    RECT 14.2000 48.8000 14.6000 49.9000 ;
	    RECT 16.1000 49.2000 16.5000 49.9000 ;
	    RECT 15.8000 48.8000 16.5000 49.2000 ;
	    RECT 12.6000 48.1000 13.0000 48.6000 ;
	    RECT 14.2000 48.1000 14.5000 48.8000 ;
	    RECT 12.6000 47.8000 14.5000 48.1000 ;
	    RECT 16.1000 48.2000 16.5000 48.8000 ;
	    RECT 16.1000 47.9000 17.0000 48.2000 ;
	    RECT 8.6000 45.8000 9.8000 46.1000 ;
	    RECT 10.6000 45.8000 12.2000 46.1000 ;
	    RECT 3.0000 45.1000 3.3000 45.8000 ;
	    RECT 3.9000 45.7000 4.3000 45.8000 ;
	    RECT 0.6000 44.8000 1.8000 45.1000 ;
	    RECT 0.6000 41.1000 1.0000 44.8000 ;
	    RECT 1.4000 44.7000 1.8000 44.8000 ;
	    RECT 2.8000 41.1000 3.6000 45.1000 ;
	    RECT 4.5000 44.8000 5.8000 45.1000 ;
	    RECT 4.5000 44.7000 4.9000 44.8000 ;
	    RECT 5.4000 41.1000 5.8000 44.8000 ;
	    RECT 7.0000 41.1000 7.4000 45.8000 ;
	    RECT 8.7000 45.1000 9.0000 45.8000 ;
	    RECT 10.6000 45.6000 11.0000 45.8000 ;
	    RECT 8.6000 41.1000 9.0000 45.1000 ;
	    RECT 9.4000 44.8000 11.4000 45.1000 ;
	    RECT 9.4000 41.1000 9.8000 44.8000 ;
	    RECT 11.0000 41.1000 11.4000 44.8000 ;
	    RECT 11.8000 41.1000 12.2000 45.8000 ;
	    RECT 14.2000 47.2000 14.5000 47.8000 ;
	    RECT 14.2000 46.8000 14.6000 47.2000 ;
	    RECT 14.2000 45.1000 14.5000 46.8000 ;
	    RECT 13.7000 44.7000 14.6000 45.1000 ;
	    RECT 13.7000 41.1000 14.1000 44.7000 ;
	    RECT 15.8000 44.4000 16.2000 45.2000 ;
	    RECT 16.6000 41.1000 17.0000 47.9000 ;
	    RECT 18.2000 47.9000 18.6000 49.9000 ;
	    RECT 20.4000 49.2000 21.2000 49.9000 ;
	    RECT 20.4000 48.8000 21.8000 49.2000 ;
	    RECT 20.4000 48.1000 21.2000 48.8000 ;
	    RECT 18.2000 47.6000 19.3000 47.9000 ;
	    RECT 17.4000 46.8000 17.8000 47.6000 ;
	    RECT 18.9000 47.5000 19.3000 47.6000 ;
	    RECT 20.2000 46.7000 20.6000 47.1000 ;
	    RECT 20.2000 46.4000 20.5000 46.7000 ;
	    RECT 19.2000 46.1000 20.5000 46.4000 ;
	    RECT 20.9000 46.4000 21.2000 48.1000 ;
	    RECT 23.0000 47.9000 23.4000 49.9000 ;
	    RECT 22.2000 47.6000 23.4000 47.9000 ;
	    RECT 22.2000 47.5000 22.6000 47.6000 ;
	    RECT 20.9000 46.2000 21.4000 46.4000 ;
	    RECT 20.9000 46.1000 21.8000 46.2000 ;
	    RECT 19.2000 46.0000 19.6000 46.1000 ;
	    RECT 21.1000 45.8000 21.8000 46.1000 ;
	    RECT 20.3000 45.7000 20.7000 45.8000 ;
	    RECT 19.0000 45.4000 20.7000 45.7000 ;
	    RECT 19.0000 45.1000 19.3000 45.4000 ;
	    RECT 21.1000 45.1000 21.4000 45.8000 ;
	    RECT 24.6000 45.1000 25.0000 49.9000 ;
	    RECT 25.7000 49.2000 26.1000 49.9000 ;
	    RECT 25.4000 48.8000 26.1000 49.2000 ;
	    RECT 28.6000 48.9000 29.0000 49.9000 ;
	    RECT 25.7000 48.2000 26.1000 48.8000 ;
	    RECT 25.7000 47.9000 26.6000 48.2000 ;
	    RECT 25.4000 45.1000 25.8000 45.2000 ;
	    RECT 18.2000 44.8000 19.3000 45.1000 ;
	    RECT 18.2000 41.1000 18.6000 44.8000 ;
	    RECT 18.9000 44.7000 19.3000 44.8000 ;
	    RECT 20.4000 44.8000 21.4000 45.1000 ;
	    RECT 22.2000 44.8000 23.4000 45.1000 ;
	    RECT 20.4000 41.1000 21.2000 44.8000 ;
	    RECT 22.2000 44.7000 22.6000 44.8000 ;
	    RECT 23.0000 41.1000 23.4000 44.8000 ;
	    RECT 24.6000 44.8000 25.8000 45.1000 ;
	    RECT 24.6000 41.1000 25.0000 44.8000 ;
	    RECT 25.4000 44.4000 25.8000 44.8000 ;
	    RECT 26.2000 41.1000 26.6000 47.9000 ;
	    RECT 27.0000 46.8000 27.4000 47.6000 ;
	    RECT 28.7000 47.2000 29.0000 48.9000 ;
	    RECT 28.6000 46.8000 29.0000 47.2000 ;
	    RECT 27.0000 46.1000 27.4000 46.2000 ;
	    RECT 28.7000 46.1000 29.0000 46.8000 ;
	    RECT 27.0000 45.8000 29.0000 46.1000 ;
	    RECT 28.7000 45.1000 29.0000 45.8000 ;
	    RECT 29.4000 46.1000 29.8000 46.2000 ;
	    RECT 30.2000 46.1000 30.6000 49.9000 ;
	    RECT 31.0000 47.8000 31.4000 48.6000 ;
	    RECT 31.8000 47.9000 32.2000 49.9000 ;
	    RECT 34.0000 48.1000 34.8000 49.9000 ;
	    RECT 31.8000 47.6000 32.9000 47.9000 ;
	    RECT 32.5000 47.5000 32.9000 47.6000 ;
	    RECT 33.8000 46.7000 34.2000 47.1000 ;
	    RECT 33.8000 46.4000 34.1000 46.7000 ;
	    RECT 29.4000 45.8000 30.6000 46.1000 ;
	    RECT 32.8000 46.1000 34.1000 46.4000 ;
	    RECT 34.5000 46.4000 34.8000 48.1000 ;
	    RECT 36.6000 47.9000 37.0000 49.9000 ;
	    RECT 35.8000 47.6000 37.0000 47.9000 ;
	    RECT 35.8000 47.5000 36.2000 47.6000 ;
	    RECT 36.2000 46.8000 37.0000 47.2000 ;
	    RECT 34.5000 46.2000 35.0000 46.4000 ;
	    RECT 34.5000 46.1000 35.4000 46.2000 ;
	    RECT 32.8000 46.0000 33.2000 46.1000 ;
	    RECT 34.7000 45.8000 35.4000 46.1000 ;
	    RECT 29.4000 45.4000 29.8000 45.8000 ;
	    RECT 28.6000 44.7000 29.5000 45.1000 ;
	    RECT 29.1000 41.1000 29.5000 44.7000 ;
	    RECT 30.2000 41.1000 30.6000 45.8000 ;
	    RECT 33.9000 45.7000 34.3000 45.8000 ;
	    RECT 32.6000 45.4000 34.3000 45.7000 ;
	    RECT 32.6000 45.1000 32.9000 45.4000 ;
	    RECT 34.7000 45.1000 35.0000 45.8000 ;
	    RECT 31.8000 44.8000 32.9000 45.1000 ;
	    RECT 31.8000 41.1000 32.2000 44.8000 ;
	    RECT 32.5000 44.7000 32.9000 44.8000 ;
	    RECT 34.0000 44.8000 35.0000 45.1000 ;
	    RECT 35.8000 44.8000 37.0000 45.1000 ;
	    RECT 34.0000 42.2000 34.8000 44.8000 ;
	    RECT 35.8000 44.7000 36.2000 44.8000 ;
	    RECT 33.4000 41.8000 34.8000 42.2000 ;
	    RECT 34.0000 41.1000 34.8000 41.8000 ;
	    RECT 36.6000 41.1000 37.0000 44.8000 ;
	    RECT 37.4000 41.1000 37.8000 49.9000 ;
	    RECT 40.3000 49.2000 40.7000 49.9000 ;
	    RECT 39.8000 48.8000 40.7000 49.2000 ;
	    RECT 38.2000 47.8000 38.6000 48.6000 ;
	    RECT 40.3000 48.2000 40.7000 48.8000 ;
	    RECT 39.8000 47.9000 40.7000 48.2000 ;
	    RECT 39.8000 41.1000 40.2000 47.9000 ;
	    RECT 40.6000 45.1000 41.0000 45.2000 ;
	    RECT 42.2000 45.1000 42.6000 49.9000 ;
	    RECT 40.6000 44.8000 42.6000 45.1000 ;
	    RECT 40.6000 44.4000 41.0000 44.8000 ;
	    RECT 42.2000 41.1000 42.6000 44.8000 ;
	    RECT 43.0000 47.7000 43.4000 49.9000 ;
	    RECT 45.1000 49.2000 45.7000 49.9000 ;
	    RECT 45.1000 48.9000 45.8000 49.2000 ;
	    RECT 47.4000 48.9000 47.8000 49.9000 ;
	    RECT 49.6000 49.2000 50.0000 49.9000 ;
	    RECT 49.6000 48.9000 50.6000 49.2000 ;
	    RECT 45.4000 48.5000 45.8000 48.9000 ;
	    RECT 47.5000 48.6000 47.8000 48.9000 ;
	    RECT 47.5000 48.3000 48.9000 48.6000 ;
	    RECT 48.5000 48.2000 48.9000 48.3000 ;
	    RECT 49.4000 48.2000 49.8000 48.6000 ;
	    RECT 50.2000 48.5000 50.6000 48.9000 ;
	    RECT 44.5000 47.7000 44.9000 47.8000 ;
	    RECT 43.0000 47.4000 44.9000 47.7000 ;
	    RECT 43.0000 45.7000 43.4000 47.4000 ;
	    RECT 46.5000 47.1000 46.9000 47.2000 ;
	    RECT 49.4000 47.1000 49.7000 48.2000 ;
	    RECT 51.8000 47.5000 52.2000 49.9000 ;
	    RECT 52.6000 47.9000 53.0000 49.9000 ;
	    RECT 54.2000 48.9000 54.6000 49.9000 ;
	    RECT 51.0000 47.1000 51.8000 47.2000 ;
	    RECT 46.3000 46.8000 51.8000 47.1000 ;
	    RECT 45.4000 46.4000 45.8000 46.5000 ;
	    RECT 43.9000 46.1000 45.8000 46.4000 ;
	    RECT 43.9000 46.0000 44.3000 46.1000 ;
	    RECT 44.7000 45.7000 45.1000 45.8000 ;
	    RECT 43.0000 45.4000 45.1000 45.7000 ;
	    RECT 43.0000 41.1000 43.4000 45.4000 ;
	    RECT 46.3000 45.2000 46.6000 46.8000 ;
	    RECT 49.9000 46.7000 50.3000 46.8000 ;
	    RECT 49.4000 46.2000 49.8000 46.3000 ;
	    RECT 50.7000 46.2000 51.1000 46.3000 ;
	    RECT 48.6000 45.9000 51.1000 46.2000 ;
	    RECT 52.6000 46.2000 52.9000 47.9000 ;
	    RECT 54.2000 47.8000 54.5000 48.9000 ;
	    RECT 55.0000 47.8000 55.4000 48.6000 ;
	    RECT 53.3000 47.5000 54.5000 47.8000 ;
	    RECT 55.8000 47.6000 56.2000 49.9000 ;
	    RECT 57.4000 48.2000 57.8000 49.9000 ;
	    RECT 57.4000 47.8000 57.9000 48.2000 ;
	    RECT 60.6000 47.8000 61.0000 48.6000 ;
	    RECT 48.6000 45.8000 49.0000 45.9000 ;
	    RECT 52.6000 45.8000 53.0000 46.2000 ;
	    RECT 53.3000 46.0000 53.6000 47.5000 ;
	    RECT 55.8000 47.3000 57.1000 47.6000 ;
	    RECT 54.1000 46.8000 54.6000 47.2000 ;
	    RECT 54.0000 46.4000 54.4000 46.8000 ;
	    RECT 55.9000 46.2000 56.3000 46.6000 ;
	    RECT 49.4000 45.5000 52.2000 45.6000 ;
	    RECT 49.3000 45.4000 52.2000 45.5000 ;
	    RECT 45.4000 44.9000 46.6000 45.2000 ;
	    RECT 47.3000 45.3000 52.2000 45.4000 ;
	    RECT 47.3000 45.1000 49.7000 45.3000 ;
	    RECT 45.4000 44.4000 45.7000 44.9000 ;
	    RECT 45.0000 44.0000 45.7000 44.4000 ;
	    RECT 46.5000 44.5000 46.9000 44.6000 ;
	    RECT 47.3000 44.5000 47.6000 45.1000 ;
	    RECT 46.5000 44.2000 47.6000 44.5000 ;
	    RECT 47.9000 44.5000 50.6000 44.8000 ;
	    RECT 47.9000 44.4000 48.3000 44.5000 ;
	    RECT 50.2000 44.4000 50.6000 44.5000 ;
	    RECT 47.1000 43.7000 47.5000 43.8000 ;
	    RECT 48.5000 43.7000 48.9000 43.8000 ;
	    RECT 45.4000 43.1000 45.8000 43.5000 ;
	    RECT 47.1000 43.4000 48.9000 43.7000 ;
	    RECT 47.5000 43.1000 47.8000 43.4000 ;
	    RECT 50.2000 43.1000 50.6000 43.5000 ;
	    RECT 45.1000 41.1000 45.7000 43.1000 ;
	    RECT 47.4000 41.1000 47.8000 43.1000 ;
	    RECT 49.6000 42.8000 50.6000 43.1000 ;
	    RECT 49.6000 41.1000 50.0000 42.8000 ;
	    RECT 51.8000 41.1000 52.2000 45.3000 ;
	    RECT 52.6000 45.1000 52.9000 45.8000 ;
	    RECT 53.3000 45.7000 53.7000 46.0000 ;
	    RECT 55.8000 45.8000 56.3000 46.2000 ;
	    RECT 56.8000 46.5000 57.1000 47.3000 ;
	    RECT 57.6000 47.2000 57.9000 47.8000 ;
	    RECT 57.4000 46.8000 57.9000 47.2000 ;
	    RECT 56.8000 46.1000 57.3000 46.5000 ;
	    RECT 53.3000 45.6000 55.4000 45.7000 ;
	    RECT 53.4000 45.4000 55.4000 45.6000 ;
	    RECT 52.6000 44.8000 53.3000 45.1000 ;
	    RECT 52.9000 41.1000 53.3000 44.8000 ;
	    RECT 55.0000 41.1000 55.4000 45.4000 ;
	    RECT 56.8000 45.1000 57.1000 46.1000 ;
	    RECT 57.6000 45.1000 57.9000 46.8000 ;
	    RECT 55.8000 44.8000 57.1000 45.1000 ;
	    RECT 55.8000 41.1000 56.2000 44.8000 ;
	    RECT 57.4000 44.6000 57.9000 45.1000 ;
	    RECT 61.4000 47.1000 61.8000 49.9000 ;
	    RECT 64.6000 48.9000 65.0000 49.9000 ;
	    RECT 66.2000 49.2000 66.6000 49.9000 ;
	    RECT 64.4000 48.8000 65.0000 48.9000 ;
	    RECT 66.1000 48.8000 66.6000 49.2000 ;
	    RECT 69.4000 48.8000 69.8000 49.9000 ;
	    RECT 64.4000 48.5000 66.4000 48.8000 ;
	    RECT 62.2000 47.1000 62.6000 47.2000 ;
	    RECT 61.4000 46.8000 62.6000 47.1000 ;
	    RECT 57.4000 41.1000 57.8000 44.6000 ;
	    RECT 61.4000 41.1000 61.8000 46.8000 ;
	    RECT 64.4000 45.2000 64.7000 48.5000 ;
	    RECT 66.5000 48.1000 67.4000 48.2000 ;
	    RECT 68.6000 48.1000 69.0000 48.6000 ;
	    RECT 66.5000 47.8000 69.0000 48.1000 ;
	    RECT 69.5000 47.2000 69.8000 48.8000 ;
	    RECT 71.0000 48.1000 71.4000 49.9000 ;
	    RECT 65.8000 46.8000 66.6000 47.2000 ;
	    RECT 69.4000 46.8000 69.8000 47.2000 ;
	    RECT 70.2000 47.8000 71.4000 48.1000 ;
	    RECT 71.8000 47.8000 72.2000 48.6000 ;
	    RECT 72.6000 47.8000 73.0000 48.6000 ;
	    RECT 73.4000 48.1000 73.8000 49.9000 ;
	    RECT 75.0000 48.9000 75.4000 49.9000 ;
	    RECT 74.2000 48.1000 74.6000 48.6000 ;
	    RECT 73.4000 47.8000 74.6000 48.1000 ;
	    RECT 70.2000 47.2000 70.5000 47.8000 ;
	    RECT 70.2000 46.8000 70.6000 47.2000 ;
	    RECT 65.0000 45.8000 65.8000 46.2000 ;
	    RECT 63.0000 44.9000 64.7000 45.2000 ;
	    RECT 69.5000 45.1000 69.8000 46.8000 ;
	    RECT 70.2000 45.4000 70.6000 46.2000 ;
	    RECT 63.0000 44.8000 63.4000 44.9000 ;
	    RECT 63.1000 44.5000 63.4000 44.8000 ;
	    RECT 69.4000 44.7000 70.3000 45.1000 ;
	    RECT 63.9000 44.5000 65.7000 44.6000 ;
	    RECT 62.2000 41.5000 62.6000 44.5000 ;
	    RECT 63.0000 41.7000 63.4000 44.5000 ;
	    RECT 63.8000 44.3000 65.7000 44.5000 ;
	    RECT 62.3000 41.4000 62.6000 41.5000 ;
	    RECT 63.8000 41.5000 64.2000 44.3000 ;
	    RECT 65.4000 44.1000 65.7000 44.3000 ;
	    RECT 66.3000 44.4000 68.1000 44.7000 ;
	    RECT 66.3000 44.1000 66.6000 44.4000 ;
	    RECT 63.8000 41.4000 64.1000 41.5000 ;
	    RECT 62.3000 41.1000 64.1000 41.4000 ;
	    RECT 64.6000 41.4000 65.0000 44.0000 ;
	    RECT 65.4000 41.7000 65.8000 44.1000 ;
	    RECT 66.2000 41.4000 66.6000 44.1000 ;
	    RECT 64.6000 41.1000 66.6000 41.4000 ;
	    RECT 67.8000 44.1000 68.1000 44.4000 ;
	    RECT 67.8000 41.1000 68.2000 44.1000 ;
	    RECT 69.9000 41.1000 70.3000 44.7000 ;
	    RECT 71.0000 41.1000 71.4000 47.8000 ;
	    RECT 73.4000 41.1000 73.8000 47.8000 ;
	    RECT 75.1000 47.2000 75.4000 48.9000 ;
	    RECT 76.6000 47.9000 77.0000 49.9000 ;
	    RECT 77.4000 48.0000 77.8000 49.9000 ;
	    RECT 79.0000 48.0000 79.4000 49.9000 ;
	    RECT 77.4000 47.9000 79.4000 48.0000 ;
	    RECT 76.7000 47.2000 77.0000 47.9000 ;
	    RECT 77.5000 47.7000 79.3000 47.9000 ;
	    RECT 79.8000 47.5000 80.2000 49.9000 ;
	    RECT 82.0000 49.2000 82.4000 49.9000 ;
	    RECT 81.4000 48.9000 82.4000 49.2000 ;
	    RECT 84.2000 48.9000 84.6000 49.9000 ;
	    RECT 86.3000 49.2000 86.9000 49.9000 ;
	    RECT 86.2000 48.9000 86.9000 49.2000 ;
	    RECT 81.4000 48.5000 81.8000 48.9000 ;
	    RECT 84.2000 48.6000 84.5000 48.9000 ;
	    RECT 82.2000 48.2000 82.6000 48.6000 ;
	    RECT 83.1000 48.3000 84.5000 48.6000 ;
	    RECT 86.2000 48.5000 86.6000 48.9000 ;
	    RECT 83.1000 48.2000 83.5000 48.3000 ;
	    RECT 78.6000 47.2000 79.0000 47.4000 ;
	    RECT 75.0000 46.8000 75.4000 47.2000 ;
	    RECT 76.6000 46.8000 77.9000 47.2000 ;
	    RECT 78.6000 46.9000 79.4000 47.2000 ;
	    RECT 79.0000 46.8000 79.4000 46.9000 ;
	    RECT 80.2000 47.1000 81.0000 47.2000 ;
	    RECT 82.3000 47.1000 82.6000 48.2000 ;
	    RECT 87.1000 47.7000 87.5000 47.8000 ;
	    RECT 88.6000 47.7000 89.0000 49.9000 ;
	    RECT 89.4000 47.9000 89.8000 49.9000 ;
	    RECT 90.2000 48.0000 90.6000 49.9000 ;
	    RECT 91.8000 48.0000 92.2000 49.9000 ;
	    RECT 90.2000 47.9000 92.2000 48.0000 ;
	    RECT 94.2000 47.9000 94.6000 49.9000 ;
	    RECT 94.9000 48.2000 95.3000 48.6000 ;
	    RECT 87.1000 47.4000 89.0000 47.7000 ;
	    RECT 85.1000 47.1000 85.5000 47.2000 ;
	    RECT 80.2000 46.8000 85.7000 47.1000 ;
	    RECT 74.2000 46.1000 74.6000 46.2000 ;
	    RECT 75.1000 46.1000 75.4000 46.8000 ;
	    RECT 74.2000 45.8000 75.4000 46.1000 ;
	    RECT 75.1000 45.1000 75.4000 45.8000 ;
	    RECT 75.8000 45.4000 76.2000 46.2000 ;
	    RECT 76.6000 45.1000 77.0000 45.2000 ;
	    RECT 77.6000 45.1000 77.9000 46.8000 ;
	    RECT 81.7000 46.7000 82.1000 46.8000 ;
	    RECT 78.2000 45.8000 78.6000 46.6000 ;
	    RECT 80.9000 46.2000 81.3000 46.3000 ;
	    RECT 82.2000 46.2000 82.6000 46.3000 ;
	    RECT 80.9000 45.9000 83.4000 46.2000 ;
	    RECT 83.0000 45.8000 83.4000 45.9000 ;
	    RECT 84.6000 46.1000 85.0000 46.2000 ;
	    RECT 85.4000 46.1000 85.7000 46.8000 ;
	    RECT 86.2000 46.4000 86.6000 46.5000 ;
	    RECT 86.2000 46.1000 88.1000 46.4000 ;
	    RECT 84.6000 45.8000 85.7000 46.1000 ;
	    RECT 87.7000 46.0000 88.1000 46.1000 ;
	    RECT 79.8000 45.5000 82.6000 45.6000 ;
	    RECT 79.8000 45.4000 82.7000 45.5000 ;
	    RECT 79.8000 45.3000 84.7000 45.4000 ;
	    RECT 75.0000 44.7000 75.9000 45.1000 ;
	    RECT 76.6000 44.8000 77.3000 45.1000 ;
	    RECT 77.6000 44.8000 78.1000 45.1000 ;
	    RECT 75.5000 41.1000 75.9000 44.7000 ;
	    RECT 77.0000 44.2000 77.3000 44.8000 ;
	    RECT 76.6000 43.8000 77.4000 44.2000 ;
	    RECT 77.7000 41.1000 78.1000 44.8000 ;
	    RECT 79.8000 41.1000 80.2000 45.3000 ;
	    RECT 82.3000 45.1000 84.7000 45.3000 ;
	    RECT 81.4000 44.5000 84.1000 44.8000 ;
	    RECT 81.4000 44.4000 81.8000 44.5000 ;
	    RECT 83.7000 44.4000 84.1000 44.5000 ;
	    RECT 84.4000 44.5000 84.7000 45.1000 ;
	    RECT 85.4000 45.2000 85.7000 45.8000 ;
	    RECT 86.9000 45.7000 87.3000 45.8000 ;
	    RECT 88.6000 45.7000 89.0000 47.4000 ;
	    RECT 89.5000 47.2000 89.8000 47.9000 ;
	    RECT 90.3000 47.7000 92.1000 47.9000 ;
	    RECT 91.4000 47.2000 91.8000 47.4000 ;
	    RECT 89.4000 46.8000 90.7000 47.2000 ;
	    RECT 91.4000 46.9000 92.2000 47.2000 ;
	    RECT 91.8000 46.8000 92.2000 46.9000 ;
	    RECT 92.6000 47.1000 93.0000 47.2000 ;
	    RECT 93.4000 47.1000 93.8000 47.2000 ;
	    RECT 92.6000 46.8000 93.8000 47.1000 ;
	    RECT 86.9000 45.4000 89.0000 45.7000 ;
	    RECT 85.4000 44.9000 86.6000 45.2000 ;
	    RECT 85.1000 44.5000 85.5000 44.6000 ;
	    RECT 84.4000 44.2000 85.5000 44.5000 ;
	    RECT 86.3000 44.4000 86.6000 44.9000 ;
	    RECT 86.3000 44.0000 87.0000 44.4000 ;
	    RECT 83.1000 43.7000 83.5000 43.8000 ;
	    RECT 84.5000 43.7000 84.9000 43.8000 ;
	    RECT 81.4000 43.1000 81.8000 43.5000 ;
	    RECT 83.1000 43.4000 84.9000 43.7000 ;
	    RECT 84.2000 43.1000 84.5000 43.4000 ;
	    RECT 86.2000 43.1000 86.6000 43.5000 ;
	    RECT 81.4000 42.8000 82.4000 43.1000 ;
	    RECT 82.0000 41.1000 82.4000 42.8000 ;
	    RECT 84.2000 41.1000 84.6000 43.1000 ;
	    RECT 86.3000 41.1000 86.9000 43.1000 ;
	    RECT 88.6000 41.1000 89.0000 45.4000 ;
	    RECT 89.4000 45.1000 89.8000 45.2000 ;
	    RECT 90.4000 45.1000 90.7000 46.8000 ;
	    RECT 91.0000 45.8000 91.4000 46.6000 ;
	    RECT 93.4000 46.4000 93.8000 46.8000 ;
	    RECT 92.6000 46.1000 93.0000 46.2000 ;
	    RECT 94.2000 46.1000 94.5000 47.9000 ;
	    RECT 95.0000 47.8000 95.4000 48.2000 ;
	    RECT 97.4000 47.9000 97.8000 49.9000 ;
	    RECT 98.1000 48.2000 98.5000 48.6000 ;
	    RECT 96.6000 46.4000 97.0000 47.2000 ;
	    RECT 95.0000 46.1000 95.4000 46.2000 ;
	    RECT 92.6000 45.8000 93.4000 46.1000 ;
	    RECT 94.2000 45.8000 95.4000 46.1000 ;
	    RECT 95.8000 46.1000 96.2000 46.2000 ;
	    RECT 97.4000 46.1000 97.7000 47.9000 ;
	    RECT 98.2000 47.8000 98.6000 48.2000 ;
	    RECT 99.0000 47.9000 99.4000 49.9000 ;
	    RECT 99.8000 48.0000 100.2000 49.9000 ;
	    RECT 101.4000 48.0000 101.8000 49.9000 ;
	    RECT 99.8000 47.9000 101.8000 48.0000 ;
	    RECT 102.2000 48.0000 102.6000 49.9000 ;
	    RECT 103.8000 48.0000 104.2000 49.9000 ;
	    RECT 102.2000 47.9000 104.2000 48.0000 ;
	    RECT 104.6000 47.9000 105.0000 49.9000 ;
	    RECT 107.0000 47.9000 107.4000 49.9000 ;
	    RECT 107.7000 48.2000 108.1000 48.6000 ;
	    RECT 99.1000 47.2000 99.4000 47.9000 ;
	    RECT 99.9000 47.7000 101.7000 47.9000 ;
	    RECT 102.3000 47.7000 104.1000 47.9000 ;
	    RECT 101.0000 47.2000 101.4000 47.4000 ;
	    RECT 102.6000 47.2000 103.0000 47.4000 ;
	    RECT 104.6000 47.2000 104.9000 47.9000 ;
	    RECT 98.2000 47.1000 98.6000 47.2000 ;
	    RECT 99.0000 47.1000 100.3000 47.2000 ;
	    RECT 98.2000 46.8000 100.3000 47.1000 ;
	    RECT 101.0000 47.1000 101.8000 47.2000 ;
	    RECT 102.2000 47.1000 103.0000 47.2000 ;
	    RECT 101.0000 46.9000 103.0000 47.1000 ;
	    RECT 103.7000 47.1000 105.0000 47.2000 ;
	    RECT 106.2000 47.1000 106.6000 47.2000 ;
	    RECT 101.4000 46.8000 102.6000 46.9000 ;
	    RECT 103.7000 46.8000 106.6000 47.1000 ;
	    RECT 98.2000 46.1000 98.6000 46.2000 ;
	    RECT 95.8000 45.8000 96.6000 46.1000 ;
	    RECT 97.4000 45.8000 98.6000 46.1000 ;
	    RECT 93.0000 45.6000 93.4000 45.8000 ;
	    RECT 95.0000 45.1000 95.3000 45.8000 ;
	    RECT 96.2000 45.6000 96.6000 45.8000 ;
	    RECT 98.2000 45.1000 98.5000 45.8000 ;
	    RECT 99.0000 45.1000 99.4000 45.2000 ;
	    RECT 100.0000 45.1000 100.3000 46.8000 ;
	    RECT 100.6000 46.1000 101.0000 46.6000 ;
	    RECT 103.0000 46.1000 103.4000 46.6000 ;
	    RECT 100.6000 45.8000 103.4000 46.1000 ;
	    RECT 103.7000 45.1000 104.0000 46.8000 ;
	    RECT 106.2000 46.4000 106.6000 46.8000 ;
	    RECT 105.4000 46.1000 105.8000 46.2000 ;
	    RECT 107.0000 46.1000 107.3000 47.9000 ;
	    RECT 107.8000 47.8000 108.2000 48.2000 ;
	    RECT 110.8000 47.1000 111.2000 49.9000 ;
	    RECT 110.3000 46.9000 111.2000 47.1000 ;
	    RECT 113.4000 47.7000 113.8000 49.9000 ;
	    RECT 115.5000 49.2000 116.1000 49.9000 ;
	    RECT 115.5000 48.9000 116.2000 49.2000 ;
	    RECT 117.8000 48.9000 118.2000 49.9000 ;
	    RECT 120.0000 49.2000 120.4000 49.9000 ;
	    RECT 120.0000 48.9000 121.0000 49.2000 ;
	    RECT 115.8000 48.5000 116.2000 48.9000 ;
	    RECT 117.9000 48.6000 118.2000 48.9000 ;
	    RECT 117.9000 48.3000 119.3000 48.6000 ;
	    RECT 118.9000 48.2000 119.3000 48.3000 ;
	    RECT 119.8000 48.2000 120.2000 48.6000 ;
	    RECT 120.6000 48.5000 121.0000 48.9000 ;
	    RECT 114.9000 47.7000 115.3000 47.8000 ;
	    RECT 113.4000 47.4000 115.3000 47.7000 ;
	    RECT 110.3000 46.8000 111.1000 46.9000 ;
	    RECT 107.8000 46.1000 108.2000 46.2000 ;
	    RECT 105.4000 45.8000 106.2000 46.1000 ;
	    RECT 107.0000 45.8000 108.2000 46.1000 ;
	    RECT 105.8000 45.6000 106.2000 45.8000 ;
	    RECT 104.6000 45.1000 105.0000 45.2000 ;
	    RECT 107.8000 45.1000 108.1000 45.8000 ;
	    RECT 110.3000 45.2000 110.6000 46.8000 ;
	    RECT 111.4000 45.8000 112.2000 46.2000 ;
	    RECT 113.4000 45.7000 113.8000 47.4000 ;
	    RECT 116.9000 47.1000 117.8000 47.2000 ;
	    RECT 119.8000 47.1000 120.1000 48.2000 ;
	    RECT 122.2000 47.5000 122.6000 49.9000 ;
	    RECT 124.3000 48.2000 124.7000 49.9000 ;
	    RECT 123.8000 47.9000 124.7000 48.2000 ;
	    RECT 126.2000 48.9000 126.6000 49.9000 ;
	    RECT 121.4000 47.1000 122.2000 47.2000 ;
	    RECT 116.7000 46.8000 122.2000 47.1000 ;
	    RECT 123.0000 46.8000 123.4000 47.6000 ;
	    RECT 115.8000 46.4000 116.2000 46.5000 ;
	    RECT 114.3000 46.1000 116.2000 46.4000 ;
	    RECT 114.3000 46.0000 114.7000 46.1000 ;
	    RECT 115.1000 45.7000 115.5000 45.8000 ;
	    RECT 109.4000 45.1000 109.8000 45.2000 ;
	    RECT 110.2000 45.1000 110.6000 45.2000 ;
	    RECT 89.4000 44.8000 90.1000 45.1000 ;
	    RECT 90.4000 44.8000 90.9000 45.1000 ;
	    RECT 89.8000 44.2000 90.1000 44.8000 ;
	    RECT 89.8000 43.8000 90.2000 44.2000 ;
	    RECT 90.5000 41.1000 90.9000 44.8000 ;
	    RECT 92.6000 44.8000 94.6000 45.1000 ;
	    RECT 92.6000 41.1000 93.0000 44.8000 ;
	    RECT 94.2000 41.1000 94.6000 44.8000 ;
	    RECT 95.0000 41.1000 95.4000 45.1000 ;
	    RECT 95.8000 44.8000 97.8000 45.1000 ;
	    RECT 95.8000 41.1000 96.2000 44.8000 ;
	    RECT 97.4000 41.1000 97.8000 44.8000 ;
	    RECT 98.2000 41.1000 98.6000 45.1000 ;
	    RECT 99.0000 44.8000 99.7000 45.1000 ;
	    RECT 100.0000 44.8000 100.5000 45.1000 ;
	    RECT 99.4000 44.2000 99.7000 44.8000 ;
	    RECT 99.0000 43.8000 99.8000 44.2000 ;
	    RECT 100.1000 41.1000 100.5000 44.8000 ;
	    RECT 103.5000 44.8000 104.0000 45.1000 ;
	    RECT 104.3000 44.8000 105.0000 45.1000 ;
	    RECT 105.4000 44.8000 107.4000 45.1000 ;
	    RECT 103.5000 41.1000 103.9000 44.8000 ;
	    RECT 104.3000 44.2000 104.6000 44.8000 ;
	    RECT 104.2000 43.8000 105.0000 44.2000 ;
	    RECT 105.4000 41.1000 105.8000 44.8000 ;
	    RECT 107.0000 41.1000 107.4000 44.8000 ;
	    RECT 107.8000 42.1000 108.2000 45.1000 ;
	    RECT 109.4000 44.8000 110.6000 45.1000 ;
	    RECT 110.3000 43.5000 110.6000 44.8000 ;
	    RECT 112.6000 44.8000 113.0000 45.6000 ;
	    RECT 113.4000 45.4000 115.5000 45.7000 ;
	    RECT 111.0000 43.8000 111.4000 44.6000 ;
	    RECT 112.6000 44.1000 112.9000 44.8000 ;
	    RECT 113.4000 44.1000 113.8000 45.4000 ;
	    RECT 116.7000 45.2000 117.0000 46.8000 ;
	    RECT 120.3000 46.7000 120.7000 46.8000 ;
	    RECT 119.8000 46.2000 120.2000 46.3000 ;
	    RECT 121.1000 46.2000 121.5000 46.3000 ;
	    RECT 119.0000 45.9000 121.5000 46.2000 ;
	    RECT 123.8000 46.1000 124.2000 47.9000 ;
	    RECT 126.2000 47.2000 126.5000 48.9000 ;
	    RECT 127.0000 47.8000 127.4000 48.6000 ;
	    RECT 127.9000 48.2000 128.3000 48.6000 ;
	    RECT 127.8000 47.8000 128.2000 48.2000 ;
	    RECT 128.6000 47.9000 129.0000 49.9000 ;
	    RECT 131.0000 47.9000 131.4000 49.9000 ;
	    RECT 133.1000 48.4000 133.5000 49.9000 ;
	    RECT 133.1000 47.9000 133.8000 48.4000 ;
	    RECT 126.2000 46.8000 126.6000 47.2000 ;
	    RECT 127.0000 47.1000 127.3000 47.8000 ;
	    RECT 128.7000 47.1000 129.0000 47.9000 ;
	    RECT 131.1000 47.8000 131.4000 47.9000 ;
	    RECT 131.1000 47.6000 132.0000 47.8000 ;
	    RECT 131.1000 47.5000 133.2000 47.6000 ;
	    RECT 131.7000 47.3000 133.2000 47.5000 ;
	    RECT 132.8000 47.2000 133.2000 47.3000 ;
	    RECT 127.0000 46.8000 129.0000 47.1000 ;
	    RECT 125.4000 46.1000 125.8000 46.2000 ;
	    RECT 119.0000 45.8000 119.4000 45.9000 ;
	    RECT 123.8000 45.8000 125.8000 46.1000 ;
	    RECT 119.8000 45.5000 122.6000 45.6000 ;
	    RECT 119.7000 45.4000 122.6000 45.5000 ;
	    RECT 115.8000 44.9000 117.0000 45.2000 ;
	    RECT 117.7000 45.3000 122.6000 45.4000 ;
	    RECT 117.7000 45.1000 120.1000 45.3000 ;
	    RECT 115.8000 44.4000 116.1000 44.9000 ;
	    RECT 112.6000 43.8000 113.8000 44.1000 ;
	    RECT 115.4000 44.0000 116.1000 44.4000 ;
	    RECT 116.9000 44.5000 117.3000 44.6000 ;
	    RECT 117.7000 44.5000 118.0000 45.1000 ;
	    RECT 116.9000 44.2000 118.0000 44.5000 ;
	    RECT 118.3000 44.5000 121.0000 44.8000 ;
	    RECT 118.3000 44.4000 118.7000 44.5000 ;
	    RECT 120.6000 44.4000 121.0000 44.5000 ;
	    RECT 110.3000 43.2000 112.1000 43.5000 ;
	    RECT 110.3000 43.1000 110.6000 43.2000 ;
	    RECT 109.4000 42.1000 109.8000 42.2000 ;
	    RECT 107.8000 41.8000 109.8000 42.1000 ;
	    RECT 107.8000 41.1000 108.2000 41.8000 ;
	    RECT 110.2000 41.1000 110.6000 43.1000 ;
	    RECT 111.8000 43.1000 112.1000 43.2000 ;
	    RECT 111.8000 41.1000 112.2000 43.1000 ;
	    RECT 113.4000 41.1000 113.8000 43.8000 ;
	    RECT 117.5000 43.7000 117.9000 43.8000 ;
	    RECT 118.9000 43.7000 119.3000 43.8000 ;
	    RECT 115.8000 43.1000 116.2000 43.5000 ;
	    RECT 117.5000 43.4000 119.3000 43.7000 ;
	    RECT 117.9000 43.1000 118.2000 43.4000 ;
	    RECT 120.6000 43.1000 121.0000 43.5000 ;
	    RECT 115.5000 41.1000 116.1000 43.1000 ;
	    RECT 117.8000 41.1000 118.2000 43.1000 ;
	    RECT 120.0000 42.8000 121.0000 43.1000 ;
	    RECT 120.0000 41.1000 120.4000 42.8000 ;
	    RECT 122.2000 41.1000 122.6000 45.3000 ;
	    RECT 123.8000 41.1000 124.2000 45.8000 ;
	    RECT 125.4000 45.4000 125.8000 45.8000 ;
	    RECT 126.2000 46.1000 126.5000 46.8000 ;
	    RECT 127.0000 46.1000 127.4000 46.2000 ;
	    RECT 126.2000 45.8000 127.4000 46.1000 ;
	    RECT 127.8000 46.1000 128.2000 46.2000 ;
	    RECT 128.7000 46.1000 129.0000 46.8000 ;
	    RECT 129.4000 46.4000 129.8000 47.2000 ;
	    RECT 131.0000 46.4000 131.4000 47.2000 ;
	    RECT 132.0000 46.9000 132.4000 47.0000 ;
	    RECT 131.9000 46.6000 132.4000 46.9000 ;
	    RECT 131.9000 46.2000 132.2000 46.6000 ;
	    RECT 130.2000 46.1000 130.6000 46.2000 ;
	    RECT 127.8000 45.8000 129.0000 46.1000 ;
	    RECT 129.8000 45.8000 130.6000 46.1000 ;
	    RECT 131.8000 45.8000 132.2000 46.2000 ;
	    RECT 124.6000 44.4000 125.0000 45.2000 ;
	    RECT 126.2000 45.1000 126.5000 45.8000 ;
	    RECT 127.9000 45.1000 128.2000 45.8000 ;
	    RECT 129.8000 45.6000 130.2000 45.8000 ;
	    RECT 132.8000 45.5000 133.1000 47.2000 ;
	    RECT 133.5000 46.2000 133.8000 47.9000 ;
	    RECT 135.0000 47.6000 135.4000 49.9000 ;
	    RECT 136.6000 47.6000 137.0000 49.9000 ;
	    RECT 138.2000 47.6000 138.6000 49.9000 ;
	    RECT 139.8000 47.6000 140.2000 49.9000 ;
	    RECT 133.4000 45.8000 133.8000 46.2000 ;
	    RECT 131.9000 45.2000 133.1000 45.5000 ;
	    RECT 125.7000 44.7000 126.6000 45.1000 ;
	    RECT 125.7000 41.1000 126.1000 44.7000 ;
	    RECT 127.8000 41.1000 128.2000 45.1000 ;
	    RECT 128.6000 44.8000 130.6000 45.1000 ;
	    RECT 128.6000 41.1000 129.0000 44.8000 ;
	    RECT 130.2000 41.1000 130.6000 44.8000 ;
	    RECT 131.9000 43.1000 132.2000 45.2000 ;
	    RECT 133.5000 45.1000 133.8000 45.8000 ;
	    RECT 134.2000 47.2000 135.4000 47.6000 ;
	    RECT 135.9000 47.2000 137.0000 47.6000 ;
	    RECT 137.5000 47.2000 138.6000 47.6000 ;
	    RECT 139.3000 47.2000 140.2000 47.6000 ;
	    RECT 141.4000 47.5000 141.8000 49.9000 ;
	    RECT 143.6000 49.2000 144.0000 49.9000 ;
	    RECT 143.0000 48.9000 144.0000 49.2000 ;
	    RECT 145.8000 48.9000 146.2000 49.9000 ;
	    RECT 147.9000 49.2000 148.5000 49.9000 ;
	    RECT 147.8000 48.9000 148.5000 49.2000 ;
	    RECT 143.0000 48.5000 143.4000 48.9000 ;
	    RECT 145.8000 48.6000 146.1000 48.9000 ;
	    RECT 143.8000 47.8000 144.2000 48.6000 ;
	    RECT 144.7000 48.3000 146.1000 48.6000 ;
	    RECT 147.8000 48.5000 148.2000 48.9000 ;
	    RECT 144.7000 48.2000 145.1000 48.3000 ;
	    RECT 147.0000 48.1000 147.4000 48.2000 ;
	    RECT 147.0000 47.8000 149.0000 48.1000 ;
	    RECT 134.2000 45.8000 134.6000 47.2000 ;
	    RECT 135.9000 46.9000 136.3000 47.2000 ;
	    RECT 137.5000 46.9000 137.9000 47.2000 ;
	    RECT 139.3000 46.9000 139.7000 47.2000 ;
	    RECT 135.0000 46.5000 136.3000 46.9000 ;
	    RECT 136.7000 46.5000 137.9000 46.9000 ;
	    RECT 138.4000 46.5000 139.7000 46.9000 ;
	    RECT 141.8000 47.1000 142.6000 47.2000 ;
	    RECT 143.9000 47.1000 144.2000 47.8000 ;
	    RECT 148.6000 47.7000 149.1000 47.8000 ;
	    RECT 150.2000 47.7000 150.6000 49.9000 ;
	    RECT 148.6000 47.4000 150.6000 47.7000 ;
	    RECT 151.0000 47.5000 151.4000 49.9000 ;
	    RECT 153.2000 49.2000 153.6000 49.9000 ;
	    RECT 152.6000 48.9000 153.6000 49.2000 ;
	    RECT 155.4000 48.9000 155.8000 49.9000 ;
	    RECT 157.5000 49.2000 158.1000 49.9000 ;
	    RECT 157.4000 48.9000 158.1000 49.2000 ;
	    RECT 152.6000 48.5000 153.0000 48.9000 ;
	    RECT 155.4000 48.6000 155.7000 48.9000 ;
	    RECT 153.4000 48.2000 153.8000 48.6000 ;
	    RECT 154.3000 48.3000 155.7000 48.6000 ;
	    RECT 157.4000 48.5000 157.8000 48.9000 ;
	    RECT 154.3000 48.2000 154.7000 48.3000 ;
	    RECT 146.7000 47.1000 147.1000 47.2000 ;
	    RECT 141.8000 46.8000 147.3000 47.1000 ;
	    RECT 143.3000 46.7000 143.7000 46.8000 ;
	    RECT 135.9000 45.8000 136.3000 46.5000 ;
	    RECT 137.5000 45.8000 137.9000 46.5000 ;
	    RECT 139.3000 45.8000 139.7000 46.5000 ;
	    RECT 142.5000 46.2000 142.9000 46.3000 ;
	    RECT 143.8000 46.2000 144.2000 46.3000 ;
	    RECT 142.5000 45.9000 145.0000 46.2000 ;
	    RECT 144.6000 45.8000 145.0000 45.9000 ;
	    RECT 134.2000 45.4000 135.4000 45.8000 ;
	    RECT 135.9000 45.4000 137.0000 45.8000 ;
	    RECT 137.5000 45.4000 138.6000 45.8000 ;
	    RECT 139.3000 45.4000 140.2000 45.8000 ;
	    RECT 131.8000 41.1000 132.2000 43.1000 ;
	    RECT 133.4000 41.1000 133.8000 45.1000 ;
	    RECT 135.0000 41.1000 135.4000 45.4000 ;
	    RECT 136.6000 41.1000 137.0000 45.4000 ;
	    RECT 138.2000 41.1000 138.6000 45.4000 ;
	    RECT 139.8000 41.1000 140.2000 45.4000 ;
	    RECT 141.4000 45.5000 144.2000 45.6000 ;
	    RECT 141.4000 45.4000 144.3000 45.5000 ;
	    RECT 141.4000 45.3000 146.3000 45.4000 ;
	    RECT 141.4000 41.1000 141.8000 45.3000 ;
	    RECT 143.9000 45.1000 146.3000 45.3000 ;
	    RECT 143.0000 44.5000 145.7000 44.8000 ;
	    RECT 143.0000 44.4000 143.4000 44.5000 ;
	    RECT 145.3000 44.4000 145.7000 44.5000 ;
	    RECT 146.0000 44.5000 146.3000 45.1000 ;
	    RECT 147.0000 45.2000 147.3000 46.8000 ;
	    RECT 147.8000 46.4000 148.2000 46.5000 ;
	    RECT 147.8000 46.1000 149.7000 46.4000 ;
	    RECT 149.3000 46.0000 149.7000 46.1000 ;
	    RECT 148.5000 45.7000 148.9000 45.8000 ;
	    RECT 150.2000 45.7000 150.6000 47.4000 ;
	    RECT 151.4000 47.1000 152.2000 47.2000 ;
	    RECT 153.5000 47.1000 153.8000 48.2000 ;
	    RECT 159.8000 48.1000 160.2000 49.9000 ;
	    RECT 163.0000 48.9000 163.4000 49.9000 ;
	    RECT 162.2000 48.1000 162.6000 48.6000 ;
	    RECT 159.8000 47.8000 162.6000 48.1000 ;
	    RECT 158.3000 47.7000 158.7000 47.8000 ;
	    RECT 159.8000 47.7000 160.2000 47.8000 ;
	    RECT 158.3000 47.4000 160.2000 47.7000 ;
	    RECT 156.3000 47.1000 156.7000 47.2000 ;
	    RECT 151.4000 46.8000 156.9000 47.1000 ;
	    RECT 152.9000 46.7000 153.3000 46.8000 ;
	    RECT 152.1000 46.2000 152.5000 46.3000 ;
	    RECT 152.1000 46.1000 154.6000 46.2000 ;
	    RECT 155.0000 46.1000 155.4000 46.2000 ;
	    RECT 152.1000 45.9000 155.4000 46.1000 ;
	    RECT 154.2000 45.8000 155.4000 45.9000 ;
	    RECT 155.8000 46.1000 156.2000 46.2000 ;
	    RECT 156.6000 46.1000 156.9000 46.8000 ;
	    RECT 157.4000 46.4000 157.8000 46.5000 ;
	    RECT 157.4000 46.1000 159.3000 46.4000 ;
	    RECT 155.8000 45.8000 156.9000 46.1000 ;
	    RECT 158.9000 46.0000 159.3000 46.1000 ;
	    RECT 148.5000 45.4000 150.6000 45.7000 ;
	    RECT 147.0000 44.9000 148.2000 45.2000 ;
	    RECT 146.7000 44.5000 147.1000 44.6000 ;
	    RECT 146.0000 44.2000 147.1000 44.5000 ;
	    RECT 147.9000 44.4000 148.2000 44.9000 ;
	    RECT 147.9000 44.0000 148.6000 44.4000 ;
	    RECT 144.7000 43.7000 145.1000 43.8000 ;
	    RECT 146.1000 43.7000 146.5000 43.8000 ;
	    RECT 143.0000 43.1000 143.4000 43.5000 ;
	    RECT 144.7000 43.4000 146.5000 43.7000 ;
	    RECT 145.8000 43.1000 146.1000 43.4000 ;
	    RECT 147.8000 43.1000 148.2000 43.5000 ;
	    RECT 143.0000 42.8000 144.0000 43.1000 ;
	    RECT 143.6000 41.1000 144.0000 42.8000 ;
	    RECT 145.8000 41.1000 146.2000 43.1000 ;
	    RECT 147.9000 41.1000 148.5000 43.1000 ;
	    RECT 150.2000 41.1000 150.6000 45.4000 ;
	    RECT 151.0000 45.5000 153.8000 45.6000 ;
	    RECT 151.0000 45.4000 153.9000 45.5000 ;
	    RECT 151.0000 45.3000 155.9000 45.4000 ;
	    RECT 151.0000 41.1000 151.4000 45.3000 ;
	    RECT 153.5000 45.1000 155.9000 45.3000 ;
	    RECT 152.6000 44.5000 155.3000 44.8000 ;
	    RECT 152.6000 44.4000 153.0000 44.5000 ;
	    RECT 154.9000 44.4000 155.3000 44.5000 ;
	    RECT 155.6000 44.5000 155.9000 45.1000 ;
	    RECT 156.6000 45.2000 156.9000 45.8000 ;
	    RECT 158.1000 45.7000 158.5000 45.8000 ;
	    RECT 159.8000 45.7000 160.2000 47.4000 ;
	    RECT 163.1000 47.2000 163.4000 48.9000 ;
	    RECT 163.0000 46.8000 163.4000 47.2000 ;
	    RECT 158.1000 45.4000 160.2000 45.7000 ;
	    RECT 156.6000 44.9000 157.8000 45.2000 ;
	    RECT 156.3000 44.5000 156.7000 44.6000 ;
	    RECT 155.6000 44.2000 156.7000 44.5000 ;
	    RECT 157.5000 44.4000 157.8000 44.9000 ;
	    RECT 158.2000 44.8000 158.6000 45.4000 ;
	    RECT 157.5000 44.0000 158.2000 44.4000 ;
	    RECT 154.3000 43.7000 154.7000 43.8000 ;
	    RECT 155.7000 43.7000 156.1000 43.8000 ;
	    RECT 152.6000 43.1000 153.0000 43.5000 ;
	    RECT 154.3000 43.4000 156.1000 43.7000 ;
	    RECT 155.4000 43.1000 155.7000 43.4000 ;
	    RECT 157.4000 43.1000 157.8000 43.5000 ;
	    RECT 152.6000 42.8000 153.6000 43.1000 ;
	    RECT 153.2000 41.1000 153.6000 42.8000 ;
	    RECT 155.4000 41.1000 155.8000 43.1000 ;
	    RECT 157.5000 41.1000 158.1000 43.1000 ;
	    RECT 159.8000 41.1000 160.2000 45.4000 ;
	    RECT 163.1000 45.1000 163.4000 46.8000 ;
	    RECT 163.8000 46.1000 164.2000 46.2000 ;
	    RECT 164.6000 46.1000 165.0000 49.9000 ;
	    RECT 165.4000 47.8000 165.8000 48.6000 ;
	    RECT 163.8000 45.8000 165.0000 46.1000 ;
	    RECT 163.8000 45.4000 164.2000 45.8000 ;
	    RECT 163.0000 44.7000 163.9000 45.1000 ;
	    RECT 163.5000 42.2000 163.9000 44.7000 ;
	    RECT 163.5000 41.8000 164.2000 42.2000 ;
	    RECT 163.5000 41.1000 163.9000 41.8000 ;
	    RECT 164.6000 41.1000 165.0000 45.8000 ;
	    RECT 166.2000 47.7000 166.6000 49.9000 ;
	    RECT 168.3000 49.2000 168.9000 49.9000 ;
	    RECT 168.3000 48.9000 169.0000 49.2000 ;
	    RECT 170.6000 48.9000 171.0000 49.9000 ;
	    RECT 172.8000 49.2000 173.2000 49.9000 ;
	    RECT 172.8000 48.9000 173.8000 49.2000 ;
	    RECT 168.6000 48.5000 169.0000 48.9000 ;
	    RECT 170.7000 48.6000 171.0000 48.9000 ;
	    RECT 170.7000 48.3000 172.1000 48.6000 ;
	    RECT 171.7000 48.2000 172.1000 48.3000 ;
	    RECT 172.6000 48.2000 173.0000 48.6000 ;
	    RECT 173.4000 48.5000 173.8000 48.9000 ;
	    RECT 167.7000 47.7000 168.1000 47.8000 ;
	    RECT 166.2000 47.4000 168.1000 47.7000 ;
	    RECT 166.2000 45.7000 166.6000 47.4000 ;
	    RECT 169.7000 47.1000 170.1000 47.2000 ;
	    RECT 172.6000 47.1000 172.9000 48.2000 ;
	    RECT 175.0000 47.5000 175.4000 49.9000 ;
	    RECT 175.8000 47.8000 176.2000 48.6000 ;
	    RECT 174.2000 47.1000 175.0000 47.2000 ;
	    RECT 169.5000 46.8000 175.0000 47.1000 ;
	    RECT 168.6000 46.4000 169.0000 46.5000 ;
	    RECT 167.1000 46.1000 169.0000 46.4000 ;
	    RECT 169.5000 46.2000 169.8000 46.8000 ;
	    RECT 173.1000 46.7000 173.5000 46.8000 ;
	    RECT 172.6000 46.2000 173.0000 46.3000 ;
	    RECT 173.9000 46.2000 174.3000 46.3000 ;
	    RECT 167.1000 46.0000 167.5000 46.1000 ;
	    RECT 169.4000 45.8000 169.8000 46.2000 ;
	    RECT 171.8000 45.9000 174.3000 46.2000 ;
	    RECT 171.8000 45.8000 172.2000 45.9000 ;
	    RECT 167.9000 45.7000 168.3000 45.8000 ;
	    RECT 166.2000 45.4000 168.3000 45.7000 ;
	    RECT 166.2000 41.1000 166.6000 45.4000 ;
	    RECT 169.5000 45.2000 169.8000 45.8000 ;
	    RECT 172.6000 45.5000 175.4000 45.6000 ;
	    RECT 172.5000 45.4000 175.4000 45.5000 ;
	    RECT 168.6000 44.9000 169.8000 45.2000 ;
	    RECT 170.5000 45.3000 175.4000 45.4000 ;
	    RECT 170.5000 45.1000 172.9000 45.3000 ;
	    RECT 168.6000 44.4000 168.9000 44.9000 ;
	    RECT 168.2000 44.0000 168.9000 44.4000 ;
	    RECT 169.7000 44.5000 170.1000 44.6000 ;
	    RECT 170.5000 44.5000 170.8000 45.1000 ;
	    RECT 169.7000 44.2000 170.8000 44.5000 ;
	    RECT 171.1000 44.5000 173.8000 44.8000 ;
	    RECT 171.1000 44.4000 171.5000 44.5000 ;
	    RECT 173.4000 44.4000 173.8000 44.5000 ;
	    RECT 170.3000 43.7000 170.7000 43.8000 ;
	    RECT 171.7000 43.7000 172.1000 43.8000 ;
	    RECT 168.6000 43.1000 169.0000 43.5000 ;
	    RECT 170.3000 43.4000 172.1000 43.7000 ;
	    RECT 170.7000 43.1000 171.0000 43.4000 ;
	    RECT 173.4000 43.1000 173.8000 43.5000 ;
	    RECT 168.3000 41.1000 168.9000 43.1000 ;
	    RECT 170.6000 41.1000 171.0000 43.1000 ;
	    RECT 172.8000 42.8000 173.8000 43.1000 ;
	    RECT 172.8000 41.1000 173.2000 42.8000 ;
	    RECT 175.0000 41.1000 175.4000 45.3000 ;
	    RECT 176.6000 41.1000 177.0000 49.9000 ;
	    RECT 177.4000 47.7000 177.8000 49.9000 ;
	    RECT 179.5000 49.2000 180.1000 49.9000 ;
	    RECT 179.5000 48.9000 180.2000 49.2000 ;
	    RECT 181.8000 48.9000 182.2000 49.9000 ;
	    RECT 184.0000 49.2000 184.4000 49.9000 ;
	    RECT 184.0000 48.9000 185.0000 49.2000 ;
	    RECT 179.8000 48.5000 180.2000 48.9000 ;
	    RECT 181.9000 48.6000 182.2000 48.9000 ;
	    RECT 181.9000 48.3000 183.3000 48.6000 ;
	    RECT 182.9000 48.2000 183.3000 48.3000 ;
	    RECT 183.8000 48.2000 184.2000 48.6000 ;
	    RECT 184.6000 48.5000 185.0000 48.9000 ;
	    RECT 178.9000 47.7000 179.3000 47.8000 ;
	    RECT 177.4000 47.4000 179.3000 47.7000 ;
	    RECT 177.4000 45.7000 177.8000 47.4000 ;
	    RECT 180.9000 47.1000 181.3000 47.2000 ;
	    RECT 183.0000 47.1000 183.4000 47.2000 ;
	    RECT 183.8000 47.1000 184.1000 48.2000 ;
	    RECT 186.2000 47.5000 186.6000 49.9000 ;
	    RECT 187.0000 47.9000 187.4000 49.9000 ;
	    RECT 189.1000 48.4000 189.5000 49.9000 ;
	    RECT 189.1000 47.9000 189.8000 48.4000 ;
	    RECT 187.1000 47.8000 187.4000 47.9000 ;
	    RECT 187.1000 47.6000 188.0000 47.8000 ;
	    RECT 187.1000 47.5000 189.2000 47.6000 ;
	    RECT 187.7000 47.3000 189.2000 47.5000 ;
	    RECT 188.8000 47.2000 189.2000 47.3000 ;
	    RECT 185.4000 47.1000 186.2000 47.2000 ;
	    RECT 180.7000 46.8000 186.2000 47.1000 ;
	    RECT 179.8000 46.4000 180.2000 46.5000 ;
	    RECT 178.3000 46.1000 180.2000 46.4000 ;
	    RECT 178.3000 46.0000 178.7000 46.1000 ;
	    RECT 179.1000 45.7000 179.5000 45.8000 ;
	    RECT 177.4000 45.4000 179.5000 45.7000 ;
	    RECT 177.4000 41.1000 177.8000 45.4000 ;
	    RECT 180.7000 45.2000 181.0000 46.8000 ;
	    RECT 184.3000 46.7000 184.7000 46.8000 ;
	    RECT 187.0000 46.4000 187.4000 47.2000 ;
	    RECT 188.0000 46.9000 188.4000 47.0000 ;
	    RECT 187.9000 46.6000 188.4000 46.9000 ;
	    RECT 185.1000 46.2000 185.5000 46.3000 ;
	    RECT 187.9000 46.2000 188.2000 46.6000 ;
	    RECT 181.4000 46.1000 181.8000 46.2000 ;
	    RECT 183.0000 46.1000 185.5000 46.2000 ;
	    RECT 181.4000 45.9000 185.5000 46.1000 ;
	    RECT 181.4000 45.8000 183.4000 45.9000 ;
	    RECT 187.8000 45.8000 188.2000 46.2000 ;
	    RECT 183.8000 45.5000 186.6000 45.6000 ;
	    RECT 188.8000 45.5000 189.1000 47.2000 ;
	    RECT 189.5000 46.2000 189.8000 47.9000 ;
	    RECT 190.2000 47.5000 190.6000 49.9000 ;
	    RECT 192.4000 49.2000 192.8000 49.9000 ;
	    RECT 191.8000 48.9000 192.8000 49.2000 ;
	    RECT 194.6000 48.9000 195.0000 49.9000 ;
	    RECT 196.7000 49.2000 197.3000 49.9000 ;
	    RECT 196.6000 48.9000 197.3000 49.2000 ;
	    RECT 191.8000 48.5000 192.2000 48.9000 ;
	    RECT 194.6000 48.6000 194.9000 48.9000 ;
	    RECT 192.6000 48.2000 193.0000 48.6000 ;
	    RECT 193.5000 48.3000 194.9000 48.6000 ;
	    RECT 196.6000 48.5000 197.0000 48.9000 ;
	    RECT 193.5000 48.2000 193.9000 48.3000 ;
	    RECT 190.6000 47.1000 191.4000 47.2000 ;
	    RECT 192.7000 47.1000 193.0000 48.2000 ;
	    RECT 197.5000 47.7000 197.9000 47.8000 ;
	    RECT 199.0000 47.7000 199.4000 49.9000 ;
	    RECT 200.1000 49.2000 200.5000 49.9000 ;
	    RECT 199.8000 48.8000 200.5000 49.2000 ;
	    RECT 200.1000 48.4000 200.5000 48.8000 ;
	    RECT 197.5000 47.4000 199.4000 47.7000 ;
	    RECT 195.5000 47.1000 195.9000 47.2000 ;
	    RECT 190.6000 46.8000 196.1000 47.1000 ;
	    RECT 192.1000 46.7000 192.5000 46.8000 ;
	    RECT 189.4000 45.8000 189.8000 46.2000 ;
	    RECT 191.3000 46.2000 191.7000 46.3000 ;
	    RECT 192.6000 46.2000 193.0000 46.3000 ;
	    RECT 195.8000 46.2000 196.1000 46.8000 ;
	    RECT 196.6000 46.4000 197.0000 46.5000 ;
	    RECT 191.3000 45.9000 193.8000 46.2000 ;
	    RECT 193.4000 45.8000 193.8000 45.9000 ;
	    RECT 195.8000 45.8000 196.2000 46.2000 ;
	    RECT 196.6000 46.1000 198.5000 46.4000 ;
	    RECT 198.1000 46.0000 198.5000 46.1000 ;
	    RECT 183.7000 45.4000 186.6000 45.5000 ;
	    RECT 179.8000 44.9000 181.0000 45.2000 ;
	    RECT 181.7000 45.3000 186.6000 45.4000 ;
	    RECT 181.7000 45.1000 184.1000 45.3000 ;
	    RECT 179.8000 44.4000 180.1000 44.9000 ;
	    RECT 179.4000 44.0000 180.1000 44.4000 ;
	    RECT 180.9000 44.5000 181.3000 44.6000 ;
	    RECT 181.7000 44.5000 182.0000 45.1000 ;
	    RECT 180.9000 44.2000 182.0000 44.5000 ;
	    RECT 182.3000 44.5000 185.0000 44.8000 ;
	    RECT 182.3000 44.4000 182.7000 44.5000 ;
	    RECT 184.6000 44.4000 185.0000 44.5000 ;
	    RECT 181.5000 43.7000 181.9000 43.8000 ;
	    RECT 182.9000 43.7000 183.3000 43.8000 ;
	    RECT 179.8000 43.1000 180.2000 43.5000 ;
	    RECT 181.5000 43.4000 183.3000 43.7000 ;
	    RECT 181.9000 43.1000 182.2000 43.4000 ;
	    RECT 184.6000 43.1000 185.0000 43.5000 ;
	    RECT 179.5000 41.1000 180.1000 43.1000 ;
	    RECT 181.8000 41.1000 182.2000 43.1000 ;
	    RECT 184.0000 42.8000 185.0000 43.1000 ;
	    RECT 184.0000 41.1000 184.4000 42.8000 ;
	    RECT 186.2000 41.1000 186.6000 45.3000 ;
	    RECT 187.9000 45.2000 189.1000 45.5000 ;
	    RECT 187.9000 43.1000 188.2000 45.2000 ;
	    RECT 189.5000 45.1000 189.8000 45.8000 ;
	    RECT 187.8000 41.1000 188.2000 43.1000 ;
	    RECT 189.4000 41.1000 189.8000 45.1000 ;
	    RECT 190.2000 45.5000 193.0000 45.6000 ;
	    RECT 190.2000 45.4000 193.1000 45.5000 ;
	    RECT 190.2000 45.3000 195.1000 45.4000 ;
	    RECT 190.2000 41.1000 190.6000 45.3000 ;
	    RECT 192.7000 45.1000 195.1000 45.3000 ;
	    RECT 191.8000 44.5000 194.5000 44.8000 ;
	    RECT 191.8000 44.4000 192.2000 44.5000 ;
	    RECT 194.1000 44.4000 194.5000 44.5000 ;
	    RECT 194.8000 44.5000 195.1000 45.1000 ;
	    RECT 195.8000 45.2000 196.1000 45.8000 ;
	    RECT 197.3000 45.7000 197.7000 45.8000 ;
	    RECT 199.0000 45.7000 199.4000 47.4000 ;
	    RECT 197.3000 45.4000 199.4000 45.7000 ;
	    RECT 195.8000 44.9000 197.0000 45.2000 ;
	    RECT 195.5000 44.5000 195.9000 44.6000 ;
	    RECT 194.8000 44.2000 195.9000 44.5000 ;
	    RECT 196.7000 44.4000 197.0000 44.9000 ;
	    RECT 196.7000 44.0000 197.4000 44.4000 ;
	    RECT 193.5000 43.7000 193.9000 43.8000 ;
	    RECT 194.9000 43.7000 195.3000 43.8000 ;
	    RECT 191.8000 43.1000 192.2000 43.5000 ;
	    RECT 193.5000 43.4000 195.3000 43.7000 ;
	    RECT 194.6000 43.1000 194.9000 43.4000 ;
	    RECT 196.6000 43.1000 197.0000 43.5000 ;
	    RECT 191.8000 42.8000 192.8000 43.1000 ;
	    RECT 192.4000 41.1000 192.8000 42.8000 ;
	    RECT 194.6000 41.1000 195.0000 43.1000 ;
	    RECT 196.7000 41.1000 197.3000 43.1000 ;
	    RECT 199.0000 41.1000 199.4000 45.4000 ;
	    RECT 199.8000 47.9000 200.5000 48.4000 ;
	    RECT 202.2000 47.9000 202.6000 49.9000 ;
	    RECT 203.0000 48.0000 203.4000 49.9000 ;
	    RECT 204.6000 48.0000 205.0000 49.9000 ;
	    RECT 203.0000 47.9000 205.0000 48.0000 ;
	    RECT 205.4000 47.9000 205.8000 49.9000 ;
	    RECT 199.8000 46.2000 200.1000 47.9000 ;
	    RECT 202.2000 47.8000 202.5000 47.9000 ;
	    RECT 201.6000 47.6000 202.5000 47.8000 ;
	    RECT 203.1000 47.7000 204.9000 47.9000 ;
	    RECT 200.4000 47.5000 202.5000 47.6000 ;
	    RECT 200.4000 47.3000 201.9000 47.5000 ;
	    RECT 200.4000 47.2000 200.8000 47.3000 ;
	    RECT 203.4000 47.2000 203.8000 47.4000 ;
	    RECT 205.4000 47.2000 205.7000 47.9000 ;
	    RECT 206.2000 47.6000 206.6000 49.9000 ;
	    RECT 206.2000 47.3000 207.3000 47.6000 ;
	    RECT 199.8000 45.8000 200.2000 46.2000 ;
	    RECT 199.8000 45.1000 200.1000 45.8000 ;
	    RECT 200.5000 45.5000 200.8000 47.2000 ;
	    RECT 202.2000 47.1000 202.6000 47.2000 ;
	    RECT 203.0000 47.1000 203.8000 47.2000 ;
	    RECT 201.2000 46.9000 201.6000 47.0000 ;
	    RECT 202.2000 46.9000 203.8000 47.1000 ;
	    RECT 201.2000 46.6000 201.7000 46.9000 ;
	    RECT 201.4000 46.2000 201.7000 46.6000 ;
	    RECT 202.2000 46.8000 203.4000 46.9000 ;
	    RECT 204.5000 46.8000 205.8000 47.2000 ;
	    RECT 201.4000 45.8000 201.8000 46.2000 ;
	    RECT 202.2000 45.8000 202.6000 46.8000 ;
	    RECT 203.8000 45.8000 204.2000 46.6000 ;
	    RECT 200.5000 45.2000 201.7000 45.5000 ;
	    RECT 199.8000 41.1000 200.2000 45.1000 ;
	    RECT 201.4000 43.1000 201.7000 45.2000 ;
	    RECT 204.5000 45.1000 204.8000 46.8000 ;
	    RECT 206.2000 46.1000 206.6000 46.6000 ;
	    RECT 205.4000 45.8000 206.6000 46.1000 ;
	    RECT 207.0000 45.8000 207.3000 47.3000 ;
	    RECT 207.8000 47.1000 208.2000 49.9000 ;
	    RECT 210.2000 47.5000 210.6000 49.9000 ;
	    RECT 212.4000 49.2000 212.8000 49.9000 ;
	    RECT 211.8000 48.9000 212.8000 49.2000 ;
	    RECT 214.6000 48.9000 215.0000 49.9000 ;
	    RECT 216.7000 49.2000 217.3000 49.9000 ;
	    RECT 216.6000 48.9000 217.3000 49.2000 ;
	    RECT 211.8000 48.5000 212.2000 48.9000 ;
	    RECT 214.6000 48.6000 214.9000 48.9000 ;
	    RECT 212.6000 48.2000 213.0000 48.6000 ;
	    RECT 213.5000 48.3000 214.9000 48.6000 ;
	    RECT 216.6000 48.5000 217.0000 48.9000 ;
	    RECT 213.5000 48.2000 213.9000 48.3000 ;
	    RECT 209.4000 47.1000 209.8000 47.2000 ;
	    RECT 207.8000 46.8000 209.8000 47.1000 ;
	    RECT 210.6000 47.1000 211.4000 47.2000 ;
	    RECT 212.7000 47.1000 213.0000 48.2000 ;
	    RECT 217.5000 47.7000 217.9000 47.8000 ;
	    RECT 219.0000 47.7000 219.4000 49.9000 ;
	    RECT 217.5000 47.4000 219.4000 47.7000 ;
	    RECT 219.8000 47.5000 220.2000 49.9000 ;
	    RECT 222.0000 49.2000 222.4000 49.9000 ;
	    RECT 221.4000 48.9000 222.4000 49.2000 ;
	    RECT 224.2000 48.9000 224.6000 49.9000 ;
	    RECT 226.3000 49.2000 226.9000 49.9000 ;
	    RECT 226.2000 48.9000 226.9000 49.2000 ;
	    RECT 221.4000 48.5000 221.8000 48.9000 ;
	    RECT 224.2000 48.6000 224.5000 48.9000 ;
	    RECT 222.2000 47.8000 222.6000 48.6000 ;
	    RECT 223.1000 48.3000 224.5000 48.6000 ;
	    RECT 226.2000 48.5000 226.6000 48.9000 ;
	    RECT 223.1000 48.2000 223.5000 48.3000 ;
	    RECT 215.5000 47.1000 215.9000 47.2000 ;
	    RECT 210.6000 46.8000 216.1000 47.1000 ;
	    RECT 207.8000 46.2000 208.2000 46.8000 ;
	    RECT 212.1000 46.7000 212.5000 46.8000 ;
	    RECT 205.4000 45.2000 205.7000 45.8000 ;
	    RECT 207.0000 45.4000 207.6000 45.8000 ;
	    RECT 205.4000 45.1000 205.8000 45.2000 ;
	    RECT 207.0000 45.1000 207.3000 45.4000 ;
	    RECT 207.9000 45.1000 208.2000 46.2000 ;
	    RECT 211.3000 46.2000 211.7000 46.3000 ;
	    RECT 212.6000 46.2000 213.0000 46.3000 ;
	    RECT 215.8000 46.2000 216.1000 46.8000 ;
	    RECT 216.6000 46.4000 217.0000 46.5000 ;
	    RECT 211.3000 45.9000 213.8000 46.2000 ;
	    RECT 213.4000 45.8000 213.8000 45.9000 ;
	    RECT 215.8000 45.8000 216.2000 46.2000 ;
	    RECT 216.6000 46.1000 218.5000 46.4000 ;
	    RECT 218.1000 46.0000 218.5000 46.1000 ;
	    RECT 204.3000 44.8000 204.8000 45.1000 ;
	    RECT 205.1000 44.8000 205.8000 45.1000 ;
	    RECT 206.2000 44.8000 207.3000 45.1000 ;
	    RECT 201.4000 41.1000 201.8000 43.1000 ;
	    RECT 204.3000 41.1000 204.7000 44.8000 ;
	    RECT 205.1000 44.2000 205.4000 44.8000 ;
	    RECT 205.0000 43.8000 205.4000 44.2000 ;
	    RECT 206.2000 41.1000 206.6000 44.8000 ;
	    RECT 207.8000 41.1000 208.2000 45.1000 ;
	    RECT 210.2000 45.5000 213.0000 45.6000 ;
	    RECT 210.2000 45.4000 213.1000 45.5000 ;
	    RECT 210.2000 45.3000 215.1000 45.4000 ;
	    RECT 210.2000 41.1000 210.6000 45.3000 ;
	    RECT 212.7000 45.1000 215.1000 45.3000 ;
	    RECT 211.8000 44.5000 214.5000 44.8000 ;
	    RECT 211.8000 44.4000 212.2000 44.5000 ;
	    RECT 214.1000 44.4000 214.5000 44.5000 ;
	    RECT 214.8000 44.5000 215.1000 45.1000 ;
	    RECT 215.8000 45.2000 216.1000 45.8000 ;
	    RECT 217.3000 45.7000 217.7000 45.8000 ;
	    RECT 219.0000 45.7000 219.4000 47.4000 ;
	    RECT 220.2000 47.1000 221.0000 47.2000 ;
	    RECT 222.3000 47.1000 222.6000 47.8000 ;
	    RECT 227.1000 47.7000 227.5000 47.8000 ;
	    RECT 228.6000 47.7000 229.0000 49.9000 ;
	    RECT 227.1000 47.4000 229.0000 47.7000 ;
	    RECT 225.1000 47.1000 225.5000 47.2000 ;
	    RECT 220.2000 46.8000 225.7000 47.1000 ;
	    RECT 221.7000 46.7000 222.1000 46.8000 ;
	    RECT 220.9000 46.2000 221.3000 46.3000 ;
	    RECT 222.2000 46.2000 222.6000 46.3000 ;
	    RECT 225.4000 46.2000 225.7000 46.8000 ;
	    RECT 226.2000 46.4000 226.6000 46.5000 ;
	    RECT 220.9000 45.9000 223.4000 46.2000 ;
	    RECT 223.0000 45.8000 223.4000 45.9000 ;
	    RECT 225.4000 45.8000 225.8000 46.2000 ;
	    RECT 226.2000 46.1000 228.1000 46.4000 ;
	    RECT 227.7000 46.0000 228.1000 46.1000 ;
	    RECT 217.3000 45.4000 219.4000 45.7000 ;
	    RECT 215.8000 44.9000 217.0000 45.2000 ;
	    RECT 215.5000 44.5000 215.9000 44.6000 ;
	    RECT 214.8000 44.2000 215.9000 44.5000 ;
	    RECT 216.7000 44.4000 217.0000 44.9000 ;
	    RECT 216.7000 44.0000 217.4000 44.4000 ;
	    RECT 213.5000 43.7000 213.9000 43.8000 ;
	    RECT 214.9000 43.7000 215.3000 43.8000 ;
	    RECT 211.8000 43.1000 212.2000 43.5000 ;
	    RECT 213.5000 43.4000 215.3000 43.7000 ;
	    RECT 214.6000 43.1000 214.9000 43.4000 ;
	    RECT 216.6000 43.1000 217.0000 43.5000 ;
	    RECT 211.8000 42.8000 212.8000 43.1000 ;
	    RECT 212.4000 41.1000 212.8000 42.8000 ;
	    RECT 214.6000 41.1000 215.0000 43.1000 ;
	    RECT 216.7000 41.1000 217.3000 43.1000 ;
	    RECT 219.0000 41.1000 219.4000 45.4000 ;
	    RECT 219.8000 45.5000 222.6000 45.6000 ;
	    RECT 219.8000 45.4000 222.7000 45.5000 ;
	    RECT 219.8000 45.3000 224.7000 45.4000 ;
	    RECT 219.8000 41.1000 220.2000 45.3000 ;
	    RECT 222.3000 45.1000 224.7000 45.3000 ;
	    RECT 221.4000 44.5000 224.1000 44.8000 ;
	    RECT 221.4000 44.4000 221.8000 44.5000 ;
	    RECT 223.7000 44.4000 224.1000 44.5000 ;
	    RECT 224.4000 44.5000 224.7000 45.1000 ;
	    RECT 225.4000 45.2000 225.7000 45.8000 ;
	    RECT 226.9000 45.7000 227.3000 45.8000 ;
	    RECT 228.6000 45.7000 229.0000 47.4000 ;
	    RECT 226.9000 45.4000 229.0000 45.7000 ;
	    RECT 225.4000 44.9000 226.6000 45.2000 ;
	    RECT 225.1000 44.5000 225.5000 44.6000 ;
	    RECT 224.4000 44.2000 225.5000 44.5000 ;
	    RECT 226.3000 44.4000 226.6000 44.9000 ;
	    RECT 226.3000 44.0000 227.0000 44.4000 ;
	    RECT 223.1000 43.7000 223.5000 43.8000 ;
	    RECT 224.5000 43.7000 224.9000 43.8000 ;
	    RECT 221.4000 43.1000 221.8000 43.5000 ;
	    RECT 223.1000 43.4000 224.9000 43.7000 ;
	    RECT 224.2000 43.1000 224.5000 43.4000 ;
	    RECT 226.2000 43.1000 226.6000 43.5000 ;
	    RECT 221.4000 42.8000 222.4000 43.1000 ;
	    RECT 222.0000 41.1000 222.4000 42.8000 ;
	    RECT 224.2000 41.1000 224.6000 43.1000 ;
	    RECT 226.3000 41.1000 226.9000 43.1000 ;
	    RECT 228.6000 41.1000 229.0000 45.4000 ;
	    RECT 229.4000 47.7000 229.8000 49.9000 ;
	    RECT 231.5000 49.2000 232.1000 49.9000 ;
	    RECT 231.5000 48.9000 232.2000 49.2000 ;
	    RECT 233.8000 48.9000 234.2000 49.9000 ;
	    RECT 236.0000 49.2000 236.4000 49.9000 ;
	    RECT 236.0000 48.9000 237.0000 49.2000 ;
	    RECT 231.8000 48.5000 232.2000 48.9000 ;
	    RECT 233.9000 48.6000 234.2000 48.9000 ;
	    RECT 233.9000 48.3000 235.3000 48.6000 ;
	    RECT 234.9000 48.2000 235.3000 48.3000 ;
	    RECT 235.8000 48.2000 236.2000 48.6000 ;
	    RECT 236.6000 48.5000 237.0000 48.9000 ;
	    RECT 230.9000 47.7000 231.3000 47.8000 ;
	    RECT 229.4000 47.4000 231.3000 47.7000 ;
	    RECT 229.4000 45.7000 229.8000 47.4000 ;
	    RECT 232.9000 47.1000 233.3000 47.2000 ;
	    RECT 235.8000 47.1000 236.1000 48.2000 ;
	    RECT 238.2000 47.5000 238.6000 49.9000 ;
	    RECT 239.0000 47.7000 239.4000 49.9000 ;
	    RECT 241.1000 49.2000 241.7000 49.9000 ;
	    RECT 241.1000 48.9000 241.8000 49.2000 ;
	    RECT 243.4000 48.9000 243.8000 49.9000 ;
	    RECT 245.6000 49.2000 246.0000 49.9000 ;
	    RECT 245.6000 48.9000 246.6000 49.2000 ;
	    RECT 241.4000 48.5000 241.8000 48.9000 ;
	    RECT 243.5000 48.6000 243.8000 48.9000 ;
	    RECT 243.5000 48.3000 244.9000 48.6000 ;
	    RECT 244.5000 48.2000 244.9000 48.3000 ;
	    RECT 245.4000 48.2000 245.8000 48.6000 ;
	    RECT 246.2000 48.5000 246.6000 48.9000 ;
	    RECT 240.5000 47.7000 240.9000 47.8000 ;
	    RECT 239.0000 47.4000 240.9000 47.7000 ;
	    RECT 237.4000 47.1000 238.2000 47.2000 ;
	    RECT 232.7000 46.8000 238.2000 47.1000 ;
	    RECT 231.8000 46.4000 232.2000 46.5000 ;
	    RECT 230.3000 46.1000 232.2000 46.4000 ;
	    RECT 232.7000 46.2000 233.0000 46.8000 ;
	    RECT 236.3000 46.7000 236.7000 46.8000 ;
	    RECT 235.8000 46.2000 236.2000 46.3000 ;
	    RECT 237.1000 46.2000 237.5000 46.3000 ;
	    RECT 230.3000 46.0000 230.7000 46.1000 ;
	    RECT 232.6000 45.8000 233.0000 46.2000 ;
	    RECT 235.0000 45.9000 237.5000 46.2000 ;
	    RECT 235.0000 45.8000 235.4000 45.9000 ;
	    RECT 231.1000 45.7000 231.5000 45.8000 ;
	    RECT 229.4000 45.4000 231.5000 45.7000 ;
	    RECT 229.4000 41.1000 229.8000 45.4000 ;
	    RECT 232.7000 45.2000 233.0000 45.8000 ;
	    RECT 239.0000 45.7000 239.4000 47.4000 ;
	    RECT 242.5000 47.1000 242.9000 47.2000 ;
	    RECT 245.4000 47.1000 245.7000 48.2000 ;
	    RECT 247.8000 47.5000 248.2000 49.9000 ;
	    RECT 248.6000 48.0000 249.0000 49.9000 ;
	    RECT 250.2000 48.0000 250.6000 49.9000 ;
	    RECT 248.6000 47.9000 250.6000 48.0000 ;
	    RECT 251.0000 47.9000 251.4000 49.9000 ;
	    RECT 251.8000 47.9000 252.2000 49.9000 ;
	    RECT 252.6000 48.0000 253.0000 49.9000 ;
	    RECT 254.2000 48.0000 254.6000 49.9000 ;
	    RECT 252.6000 47.9000 254.6000 48.0000 ;
	    RECT 256.6000 47.9000 257.0000 49.9000 ;
	    RECT 257.3000 48.2000 257.7000 48.6000 ;
	    RECT 248.7000 47.7000 250.5000 47.9000 ;
	    RECT 249.0000 47.2000 249.4000 47.4000 ;
	    RECT 251.0000 47.2000 251.3000 47.9000 ;
	    RECT 251.9000 47.2000 252.2000 47.9000 ;
	    RECT 252.7000 47.7000 254.5000 47.9000 ;
	    RECT 253.8000 47.2000 254.2000 47.4000 ;
	    RECT 247.0000 47.1000 247.8000 47.2000 ;
	    RECT 242.3000 46.8000 247.8000 47.1000 ;
	    RECT 248.6000 46.9000 249.4000 47.2000 ;
	    RECT 248.6000 46.8000 249.0000 46.9000 ;
	    RECT 250.1000 46.8000 251.4000 47.2000 ;
	    RECT 251.8000 46.8000 253.1000 47.2000 ;
	    RECT 253.8000 46.9000 254.6000 47.2000 ;
	    RECT 254.2000 46.8000 254.6000 46.9000 ;
	    RECT 241.4000 46.4000 241.8000 46.5000 ;
	    RECT 239.9000 46.1000 241.8000 46.4000 ;
	    RECT 242.3000 46.2000 242.6000 46.8000 ;
	    RECT 245.9000 46.7000 246.3000 46.8000 ;
	    RECT 245.4000 46.2000 245.8000 46.3000 ;
	    RECT 246.7000 46.2000 247.1000 46.3000 ;
	    RECT 239.9000 46.0000 240.3000 46.1000 ;
	    RECT 242.2000 45.8000 242.6000 46.2000 ;
	    RECT 244.6000 45.9000 247.1000 46.2000 ;
	    RECT 244.6000 45.8000 245.0000 45.9000 ;
	    RECT 240.7000 45.7000 241.1000 45.8000 ;
	    RECT 235.8000 45.5000 238.6000 45.6000 ;
	    RECT 235.7000 45.4000 238.6000 45.5000 ;
	    RECT 231.8000 44.9000 233.0000 45.2000 ;
	    RECT 233.7000 45.3000 238.6000 45.4000 ;
	    RECT 233.7000 45.1000 236.1000 45.3000 ;
	    RECT 231.8000 44.4000 232.1000 44.9000 ;
	    RECT 231.4000 44.0000 232.1000 44.4000 ;
	    RECT 232.9000 44.5000 233.3000 44.6000 ;
	    RECT 233.7000 44.5000 234.0000 45.1000 ;
	    RECT 232.9000 44.2000 234.0000 44.5000 ;
	    RECT 234.3000 44.5000 237.0000 44.8000 ;
	    RECT 234.3000 44.4000 234.7000 44.5000 ;
	    RECT 236.6000 44.4000 237.0000 44.5000 ;
	    RECT 233.5000 43.7000 233.9000 43.8000 ;
	    RECT 234.9000 43.7000 235.3000 43.8000 ;
	    RECT 231.8000 43.1000 232.2000 43.5000 ;
	    RECT 233.5000 43.4000 235.3000 43.7000 ;
	    RECT 233.9000 43.1000 234.2000 43.4000 ;
	    RECT 236.6000 43.1000 237.0000 43.5000 ;
	    RECT 231.5000 41.1000 232.1000 43.1000 ;
	    RECT 233.8000 41.1000 234.2000 43.1000 ;
	    RECT 236.0000 42.8000 237.0000 43.1000 ;
	    RECT 236.0000 41.1000 236.4000 42.8000 ;
	    RECT 238.2000 41.1000 238.6000 45.3000 ;
	    RECT 239.0000 45.4000 241.1000 45.7000 ;
	    RECT 239.0000 41.1000 239.4000 45.4000 ;
	    RECT 242.3000 45.2000 242.6000 45.8000 ;
	    RECT 245.4000 45.5000 248.2000 45.6000 ;
	    RECT 245.3000 45.4000 248.2000 45.5000 ;
	    RECT 241.4000 44.9000 242.6000 45.2000 ;
	    RECT 243.3000 45.3000 248.2000 45.4000 ;
	    RECT 243.3000 45.1000 245.7000 45.3000 ;
	    RECT 241.4000 44.4000 241.7000 44.9000 ;
	    RECT 241.0000 44.0000 241.7000 44.4000 ;
	    RECT 242.5000 44.5000 242.9000 44.6000 ;
	    RECT 243.3000 44.5000 243.6000 45.1000 ;
	    RECT 242.5000 44.2000 243.6000 44.5000 ;
	    RECT 243.9000 44.5000 246.6000 44.8000 ;
	    RECT 243.9000 44.4000 244.3000 44.5000 ;
	    RECT 246.2000 44.4000 246.6000 44.5000 ;
	    RECT 243.1000 43.7000 243.5000 43.8000 ;
	    RECT 244.5000 43.7000 244.9000 43.8000 ;
	    RECT 241.4000 43.1000 241.8000 43.5000 ;
	    RECT 243.1000 43.4000 244.9000 43.7000 ;
	    RECT 243.5000 43.1000 243.8000 43.4000 ;
	    RECT 246.2000 43.1000 246.6000 43.5000 ;
	    RECT 241.1000 41.1000 241.7000 43.1000 ;
	    RECT 243.4000 41.1000 243.8000 43.1000 ;
	    RECT 245.6000 42.8000 246.6000 43.1000 ;
	    RECT 245.6000 41.1000 246.0000 42.8000 ;
	    RECT 247.8000 41.1000 248.2000 45.3000 ;
	    RECT 250.1000 45.1000 250.4000 46.8000 ;
	    RECT 249.9000 44.8000 250.4000 45.1000 ;
	    RECT 251.8000 45.1000 252.2000 45.2000 ;
	    RECT 252.8000 45.1000 253.1000 46.8000 ;
	    RECT 253.4000 45.8000 253.8000 46.6000 ;
	    RECT 255.8000 46.4000 256.2000 47.2000 ;
	    RECT 255.0000 46.1000 255.4000 46.2000 ;
	    RECT 256.6000 46.1000 256.9000 47.9000 ;
	    RECT 257.4000 47.8000 257.8000 48.2000 ;
	    RECT 258.2000 47.7000 258.6000 49.9000 ;
	    RECT 260.3000 49.2000 260.9000 49.9000 ;
	    RECT 260.3000 48.9000 261.0000 49.2000 ;
	    RECT 262.6000 48.9000 263.0000 49.9000 ;
	    RECT 264.8000 49.2000 265.2000 49.9000 ;
	    RECT 264.8000 48.9000 265.8000 49.2000 ;
	    RECT 260.6000 48.5000 261.0000 48.9000 ;
	    RECT 262.7000 48.6000 263.0000 48.9000 ;
	    RECT 262.7000 48.3000 264.1000 48.6000 ;
	    RECT 263.7000 48.2000 264.1000 48.3000 ;
	    RECT 264.6000 48.2000 265.0000 48.6000 ;
	    RECT 265.4000 48.5000 265.8000 48.9000 ;
	    RECT 259.7000 47.7000 260.1000 47.8000 ;
	    RECT 258.2000 47.4000 260.1000 47.7000 ;
	    RECT 257.4000 46.1000 257.8000 46.2000 ;
	    RECT 255.0000 45.8000 255.8000 46.1000 ;
	    RECT 256.6000 45.8000 257.8000 46.1000 ;
	    RECT 255.4000 45.6000 255.8000 45.8000 ;
	    RECT 257.4000 45.1000 257.7000 45.8000 ;
	    RECT 258.2000 45.7000 258.6000 47.4000 ;
	    RECT 261.7000 47.1000 262.1000 47.2000 ;
	    RECT 264.6000 47.1000 264.9000 48.2000 ;
	    RECT 267.0000 47.5000 267.4000 49.9000 ;
	    RECT 268.1000 49.2000 268.5000 49.9000 ;
	    RECT 268.1000 48.8000 269.0000 49.2000 ;
	    RECT 268.1000 48.2000 268.5000 48.8000 ;
	    RECT 268.1000 47.9000 269.0000 48.2000 ;
	    RECT 266.2000 47.1000 267.0000 47.2000 ;
	    RECT 261.5000 46.8000 267.0000 47.1000 ;
	    RECT 260.6000 46.4000 261.0000 46.5000 ;
	    RECT 259.1000 46.1000 261.0000 46.4000 ;
	    RECT 261.5000 46.2000 261.8000 46.8000 ;
	    RECT 265.1000 46.7000 265.5000 46.8000 ;
	    RECT 264.6000 46.2000 265.0000 46.3000 ;
	    RECT 265.9000 46.2000 266.3000 46.3000 ;
	    RECT 259.1000 46.0000 259.5000 46.1000 ;
	    RECT 261.4000 45.8000 261.8000 46.2000 ;
	    RECT 263.8000 45.9000 266.3000 46.2000 ;
	    RECT 263.8000 45.8000 264.2000 45.9000 ;
	    RECT 259.9000 45.7000 260.3000 45.8000 ;
	    RECT 258.2000 45.4000 260.3000 45.7000 ;
	    RECT 251.8000 44.8000 252.5000 45.1000 ;
	    RECT 252.8000 44.8000 253.3000 45.1000 ;
	    RECT 249.9000 41.1000 250.3000 44.8000 ;
	    RECT 252.2000 44.2000 252.5000 44.8000 ;
	    RECT 252.2000 43.8000 252.6000 44.2000 ;
	    RECT 252.9000 41.1000 253.3000 44.8000 ;
	    RECT 255.0000 44.8000 257.0000 45.1000 ;
	    RECT 255.0000 41.1000 255.4000 44.8000 ;
	    RECT 256.6000 41.1000 257.0000 44.8000 ;
	    RECT 257.4000 41.1000 257.8000 45.1000 ;
	    RECT 258.2000 41.1000 258.6000 45.4000 ;
	    RECT 261.5000 45.2000 261.8000 45.8000 ;
	    RECT 264.6000 45.5000 267.4000 45.6000 ;
	    RECT 264.5000 45.4000 267.4000 45.5000 ;
	    RECT 260.6000 44.9000 261.8000 45.2000 ;
	    RECT 262.5000 45.3000 267.4000 45.4000 ;
	    RECT 262.5000 45.1000 264.9000 45.3000 ;
	    RECT 260.6000 44.4000 260.9000 44.9000 ;
	    RECT 260.2000 44.0000 260.9000 44.4000 ;
	    RECT 261.7000 44.5000 262.1000 44.6000 ;
	    RECT 262.5000 44.5000 262.8000 45.1000 ;
	    RECT 261.7000 44.2000 262.8000 44.5000 ;
	    RECT 263.1000 44.5000 265.8000 44.8000 ;
	    RECT 263.1000 44.4000 263.5000 44.5000 ;
	    RECT 265.4000 44.4000 265.8000 44.5000 ;
	    RECT 262.3000 43.7000 262.7000 43.8000 ;
	    RECT 263.7000 43.7000 264.1000 43.8000 ;
	    RECT 260.6000 43.1000 261.0000 43.5000 ;
	    RECT 262.3000 43.4000 264.1000 43.7000 ;
	    RECT 262.7000 43.1000 263.0000 43.4000 ;
	    RECT 265.4000 43.1000 265.8000 43.5000 ;
	    RECT 260.3000 41.1000 260.9000 43.1000 ;
	    RECT 262.6000 41.1000 263.0000 43.1000 ;
	    RECT 264.8000 42.8000 265.8000 43.1000 ;
	    RECT 264.8000 41.1000 265.2000 42.8000 ;
	    RECT 267.0000 41.1000 267.4000 45.3000 ;
	    RECT 267.8000 44.4000 268.2000 45.2000 ;
	    RECT 268.6000 41.1000 269.0000 47.9000 ;
	    RECT 0.6000 36.2000 1.0000 39.9000 ;
	    RECT 2.8000 37.2000 3.6000 39.9000 ;
	    RECT 2.8000 36.8000 4.2000 37.2000 ;
	    RECT 1.3000 36.2000 1.7000 36.3000 ;
	    RECT 0.6000 35.9000 1.7000 36.2000 ;
	    RECT 2.8000 36.2000 3.6000 36.8000 ;
	    RECT 4.6000 36.2000 5.0000 36.3000 ;
	    RECT 5.4000 36.2000 5.8000 39.9000 ;
	    RECT 2.8000 35.9000 3.8000 36.2000 ;
	    RECT 4.6000 35.9000 5.8000 36.2000 ;
	    RECT 6.2000 36.2000 6.6000 39.9000 ;
	    RECT 7.1000 36.2000 7.5000 36.3000 ;
	    RECT 6.2000 35.9000 7.5000 36.2000 ;
	    RECT 8.4000 35.9000 9.2000 39.9000 ;
	    RECT 10.2000 36.2000 10.6000 36.3000 ;
	    RECT 11.0000 36.2000 11.4000 39.9000 ;
	    RECT 10.2000 35.9000 11.4000 36.2000 ;
	    RECT 1.4000 35.6000 1.7000 35.9000 ;
	    RECT 1.4000 35.3000 3.1000 35.6000 ;
	    RECT 2.7000 35.2000 3.1000 35.3000 ;
	    RECT 3.5000 35.2000 3.8000 35.9000 ;
	    RECT 7.7000 35.2000 8.1000 35.3000 ;
	    RECT 8.7000 35.2000 9.0000 35.9000 ;
	    RECT 1.6000 34.9000 2.0000 35.0000 ;
	    RECT 3.5000 34.9000 4.2000 35.2000 ;
	    RECT 1.6000 34.6000 2.9000 34.9000 ;
	    RECT 2.6000 34.3000 2.9000 34.6000 ;
	    RECT 3.3000 34.8000 4.2000 34.9000 ;
	    RECT 7.3000 34.9000 8.1000 35.2000 ;
	    RECT 7.3000 34.8000 7.7000 34.9000 ;
	    RECT 8.6000 34.8000 9.0000 35.2000 ;
	    RECT 11.8000 35.1000 12.2000 35.2000 ;
	    RECT 12.6000 35.1000 13.0000 39.9000 ;
	    RECT 11.8000 34.8000 13.0000 35.1000 ;
	    RECT 3.3000 34.6000 3.8000 34.8000 ;
	    RECT 2.6000 33.9000 3.0000 34.3000 ;
	    RECT 1.3000 33.4000 1.7000 33.5000 ;
	    RECT 0.6000 33.1000 1.7000 33.4000 ;
	    RECT 0.6000 31.1000 1.0000 33.1000 ;
	    RECT 3.3000 32.9000 3.6000 34.6000 ;
	    RECT 8.7000 34.2000 9.0000 34.8000 ;
	    RECT 8.7000 33.9000 9.2000 34.2000 ;
	    RECT 4.6000 33.4000 5.0000 33.5000 ;
	    RECT 7.1000 33.4000 7.5000 33.5000 ;
	    RECT 4.6000 33.1000 5.8000 33.4000 ;
	    RECT 2.8000 31.1000 3.6000 32.9000 ;
	    RECT 5.4000 31.1000 5.8000 33.1000 ;
	    RECT 6.2000 33.1000 7.5000 33.4000 ;
	    RECT 7.8000 33.2000 8.6000 33.6000 ;
	    RECT 6.2000 31.1000 6.6000 33.1000 ;
	    RECT 8.9000 32.9000 9.2000 33.9000 ;
	    RECT 9.6000 33.8000 10.0000 34.2000 ;
	    RECT 9.6000 33.6000 9.9000 33.8000 ;
	    RECT 9.5000 33.2000 9.9000 33.6000 ;
	    RECT 10.2000 33.4000 10.6000 33.5000 ;
	    RECT 10.2000 33.1000 11.4000 33.4000 ;
	    RECT 8.4000 32.2000 9.2000 32.9000 ;
	    RECT 8.4000 31.8000 9.8000 32.2000 ;
	    RECT 8.4000 31.1000 9.2000 31.8000 ;
	    RECT 11.0000 31.1000 11.4000 33.1000 ;
	    RECT 12.6000 31.1000 13.0000 34.8000 ;
	    RECT 14.2000 34.1000 14.6000 39.9000 ;
	    RECT 15.0000 35.8000 15.4000 36.6000 ;
	    RECT 16.1000 36.3000 16.5000 39.9000 ;
	    RECT 19.3000 39.2000 19.7000 39.9000 ;
	    RECT 19.3000 38.8000 20.2000 39.2000 ;
	    RECT 18.6000 36.8000 19.0000 37.2000 ;
	    RECT 16.1000 35.9000 17.0000 36.3000 ;
	    RECT 18.6000 36.2000 18.9000 36.8000 ;
	    RECT 19.3000 36.2000 19.7000 38.8000 ;
	    RECT 22.7000 36.3000 23.1000 39.9000 ;
	    RECT 18.2000 35.9000 18.9000 36.2000 ;
	    RECT 19.2000 35.9000 19.7000 36.2000 ;
	    RECT 22.2000 35.9000 23.1000 36.3000 ;
	    RECT 15.0000 35.1000 15.4000 35.2000 ;
	    RECT 15.8000 35.1000 16.2000 35.6000 ;
	    RECT 15.0000 34.8000 16.2000 35.1000 ;
	    RECT 16.6000 34.2000 16.9000 35.9000 ;
	    RECT 18.2000 35.8000 18.6000 35.9000 ;
	    RECT 19.2000 34.2000 19.5000 35.9000 ;
	    RECT 19.8000 34.4000 20.2000 35.2000 ;
	    RECT 22.3000 34.2000 22.6000 35.9000 ;
	    RECT 15.0000 34.1000 15.4000 34.2000 ;
	    RECT 14.2000 33.8000 15.4000 34.1000 ;
	    RECT 15.8000 34.1000 16.2000 34.2000 ;
	    RECT 16.6000 34.1000 17.0000 34.2000 ;
	    RECT 15.8000 33.8000 17.0000 34.1000 ;
	    RECT 18.2000 33.8000 19.5000 34.2000 ;
	    RECT 20.6000 34.1000 21.0000 34.2000 ;
	    RECT 20.2000 33.8000 21.0000 34.1000 ;
	    RECT 22.2000 34.1000 22.6000 34.2000 ;
	    RECT 23.8000 34.8000 24.2000 35.2000 ;
	    RECT 24.6000 35.1000 25.0000 39.9000 ;
	    RECT 26.7000 36.2000 27.1000 39.9000 ;
	    RECT 27.4000 36.8000 27.8000 37.2000 ;
	    RECT 27.5000 36.2000 27.8000 36.8000 ;
	    RECT 29.9000 36.3000 30.3000 39.9000 ;
	    RECT 26.7000 35.9000 27.2000 36.2000 ;
	    RECT 27.5000 35.9000 28.2000 36.2000 ;
	    RECT 29.4000 35.9000 30.3000 36.3000 ;
	    RECT 31.3000 39.2000 31.7000 39.9000 ;
	    RECT 31.3000 38.8000 32.2000 39.2000 ;
	    RECT 31.3000 36.3000 31.7000 38.8000 ;
	    RECT 31.3000 35.9000 32.2000 36.3000 ;
	    RECT 26.2000 35.1000 26.6000 35.2000 ;
	    RECT 24.6000 34.8000 26.6000 35.1000 ;
	    RECT 23.8000 34.1000 24.1000 34.8000 ;
	    RECT 22.2000 33.8000 24.1000 34.1000 ;
	    RECT 14.2000 33.1000 14.6000 33.8000 ;
	    RECT 14.2000 32.8000 15.1000 33.1000 ;
	    RECT 14.7000 31.1000 15.1000 32.8000 ;
	    RECT 16.6000 32.1000 16.9000 33.8000 ;
	    RECT 18.3000 33.1000 18.6000 33.8000 ;
	    RECT 20.2000 33.6000 20.6000 33.8000 ;
	    RECT 19.1000 33.1000 20.9000 33.3000 ;
	    RECT 16.6000 31.1000 17.0000 32.1000 ;
	    RECT 18.2000 31.1000 18.6000 33.1000 ;
	    RECT 19.0000 33.0000 21.0000 33.1000 ;
	    RECT 19.0000 31.1000 19.4000 33.0000 ;
	    RECT 20.6000 31.1000 21.0000 33.0000 ;
	    RECT 22.3000 32.2000 22.6000 33.8000 ;
	    RECT 23.8000 32.4000 24.2000 33.2000 ;
	    RECT 22.2000 31.1000 22.6000 32.2000 ;
	    RECT 24.6000 31.1000 25.0000 34.8000 ;
	    RECT 26.2000 34.4000 26.6000 34.8000 ;
	    RECT 26.9000 35.1000 27.2000 35.9000 ;
	    RECT 27.8000 35.8000 28.2000 35.9000 ;
	    RECT 27.8000 35.1000 28.2000 35.2000 ;
	    RECT 26.9000 34.8000 28.2000 35.1000 ;
	    RECT 26.9000 34.2000 27.2000 34.8000 ;
	    RECT 29.5000 34.2000 29.8000 35.9000 ;
	    RECT 30.2000 34.8000 30.6000 35.6000 ;
	    RECT 31.0000 34.8000 31.4000 35.6000 ;
	    RECT 25.4000 34.1000 25.8000 34.2000 ;
	    RECT 25.4000 33.8000 26.2000 34.1000 ;
	    RECT 26.9000 33.8000 28.2000 34.2000 ;
	    RECT 29.4000 33.8000 29.8000 34.2000 ;
	    RECT 25.8000 33.6000 26.2000 33.8000 ;
	    RECT 25.5000 33.1000 27.3000 33.3000 ;
	    RECT 27.8000 33.1000 28.1000 33.8000 ;
	    RECT 25.4000 33.0000 27.4000 33.1000 ;
	    RECT 25.4000 31.1000 25.8000 33.0000 ;
	    RECT 27.0000 31.1000 27.4000 33.0000 ;
	    RECT 27.8000 31.1000 28.2000 33.1000 ;
	    RECT 29.5000 32.2000 29.8000 33.8000 ;
	    RECT 29.4000 31.1000 29.8000 32.2000 ;
	    RECT 31.8000 34.2000 32.1000 35.9000 ;
	    RECT 33.4000 35.8000 33.8000 36.6000 ;
	    RECT 31.8000 33.8000 32.2000 34.2000 ;
	    RECT 31.8000 32.1000 32.1000 33.8000 ;
	    RECT 32.6000 33.1000 33.0000 33.2000 ;
	    RECT 34.2000 33.1000 34.6000 39.9000 ;
	    RECT 35.8000 36.2000 36.2000 39.9000 ;
	    RECT 36.6000 36.2000 37.0000 36.3000 ;
	    RECT 38.0000 36.2000 38.8000 39.9000 ;
	    RECT 35.8000 35.9000 37.0000 36.2000 ;
	    RECT 37.8000 35.9000 38.8000 36.2000 ;
	    RECT 39.9000 36.2000 40.3000 36.3000 ;
	    RECT 40.6000 36.2000 41.0000 39.9000 ;
	    RECT 39.9000 35.9000 41.0000 36.2000 ;
	    RECT 37.8000 35.2000 38.1000 35.9000 ;
	    RECT 39.9000 35.6000 40.2000 35.9000 ;
	    RECT 38.5000 35.3000 40.2000 35.6000 ;
	    RECT 38.5000 35.2000 38.9000 35.3000 ;
	    RECT 37.4000 35.1000 38.1000 35.2000 ;
	    RECT 35.0000 34.9000 38.1000 35.1000 ;
	    RECT 39.6000 34.9000 40.0000 35.0000 ;
	    RECT 35.0000 34.8000 38.3000 34.9000 ;
	    RECT 35.0000 34.2000 35.3000 34.8000 ;
	    RECT 37.8000 34.6000 38.3000 34.8000 ;
	    RECT 35.0000 33.4000 35.4000 34.2000 ;
	    RECT 36.6000 33.4000 37.0000 33.5000 ;
	    RECT 32.6000 32.8000 34.6000 33.1000 ;
	    RECT 35.8000 33.1000 37.0000 33.4000 ;
	    RECT 32.6000 32.4000 33.0000 32.8000 ;
	    RECT 31.8000 31.1000 32.2000 32.1000 ;
	    RECT 33.7000 31.1000 34.1000 32.8000 ;
	    RECT 35.8000 31.1000 36.2000 33.1000 ;
	    RECT 38.0000 32.9000 38.3000 34.6000 ;
	    RECT 38.7000 34.6000 40.0000 34.9000 ;
	    RECT 38.7000 34.3000 39.0000 34.6000 ;
	    RECT 38.6000 33.9000 39.0000 34.3000 ;
	    RECT 39.9000 33.4000 40.3000 33.5000 ;
	    RECT 39.9000 33.1000 41.0000 33.4000 ;
	    RECT 38.0000 31.1000 38.8000 32.9000 ;
	    RECT 40.6000 31.1000 41.0000 33.1000 ;
	    RECT 41.4000 32.4000 41.8000 33.2000 ;
	    RECT 42.2000 33.1000 42.6000 39.9000 ;
	    RECT 44.3000 36.3000 44.7000 39.9000 ;
	    RECT 43.8000 35.9000 44.7000 36.3000 ;
	    RECT 43.9000 34.2000 44.2000 35.9000 ;
	    RECT 44.6000 34.8000 45.0000 35.6000 ;
	    RECT 43.8000 33.8000 44.2000 34.2000 ;
	    RECT 43.0000 33.1000 43.4000 33.2000 ;
	    RECT 42.2000 32.8000 43.4000 33.1000 ;
	    RECT 42.2000 31.1000 42.6000 32.8000 ;
	    RECT 43.0000 32.4000 43.4000 32.8000 ;
	    RECT 43.9000 32.2000 44.2000 33.8000 ;
	    RECT 45.4000 33.4000 45.8000 34.2000 ;
	    RECT 43.8000 31.1000 44.2000 32.2000 ;
	    RECT 46.2000 31.1000 46.6000 39.9000 ;
	    RECT 47.8000 36.4000 48.2000 39.9000 ;
	    RECT 47.7000 35.9000 48.2000 36.4000 ;
	    RECT 49.4000 36.2000 49.8000 39.9000 ;
	    RECT 48.5000 35.9000 49.8000 36.2000 ;
	    RECT 47.7000 34.2000 48.0000 35.9000 ;
	    RECT 48.5000 34.9000 48.8000 35.9000 ;
	    RECT 50.2000 35.6000 50.6000 39.9000 ;
	    RECT 52.3000 37.9000 52.9000 39.9000 ;
	    RECT 54.6000 37.9000 55.0000 39.9000 ;
	    RECT 56.8000 38.2000 57.2000 39.9000 ;
	    RECT 56.8000 37.9000 57.8000 38.2000 ;
	    RECT 52.6000 37.5000 53.0000 37.9000 ;
	    RECT 54.7000 37.6000 55.0000 37.9000 ;
	    RECT 54.3000 37.3000 56.1000 37.6000 ;
	    RECT 57.4000 37.5000 57.8000 37.9000 ;
	    RECT 54.3000 37.2000 54.7000 37.3000 ;
	    RECT 55.7000 37.2000 56.1000 37.3000 ;
	    RECT 52.2000 36.6000 52.9000 37.0000 ;
	    RECT 52.6000 36.1000 52.9000 36.6000 ;
	    RECT 53.7000 36.5000 54.8000 36.8000 ;
	    RECT 53.7000 36.4000 54.1000 36.5000 ;
	    RECT 52.6000 35.8000 53.8000 36.1000 ;
	    RECT 50.2000 35.3000 52.3000 35.6000 ;
	    RECT 48.3000 34.5000 48.8000 34.9000 ;
	    RECT 47.0000 34.1000 47.4000 34.2000 ;
	    RECT 47.7000 34.1000 48.2000 34.2000 ;
	    RECT 47.0000 33.8000 48.2000 34.1000 ;
	    RECT 47.7000 33.1000 48.0000 33.8000 ;
	    RECT 48.5000 33.7000 48.8000 34.5000 ;
	    RECT 49.3000 34.8000 49.8000 35.2000 ;
	    RECT 49.3000 34.4000 49.7000 34.8000 ;
	    RECT 48.5000 33.4000 49.8000 33.7000 ;
	    RECT 47.7000 32.8000 48.2000 33.1000 ;
	    RECT 47.8000 31.1000 48.2000 32.8000 ;
	    RECT 49.4000 31.1000 49.8000 33.4000 ;
	    RECT 50.2000 33.6000 50.6000 35.3000 ;
	    RECT 51.9000 35.2000 52.3000 35.3000 ;
	    RECT 53.5000 35.2000 53.8000 35.8000 ;
	    RECT 54.5000 35.9000 54.8000 36.5000 ;
	    RECT 55.1000 36.5000 55.5000 36.6000 ;
	    RECT 57.4000 36.5000 57.8000 36.6000 ;
	    RECT 55.1000 36.2000 57.8000 36.5000 ;
	    RECT 54.5000 35.7000 56.9000 35.9000 ;
	    RECT 59.0000 35.7000 59.4000 39.9000 ;
	    RECT 61.4000 37.9000 61.8000 39.9000 ;
	    RECT 61.5000 37.8000 61.8000 37.9000 ;
	    RECT 63.0000 37.9000 63.4000 39.9000 ;
	    RECT 63.0000 37.8000 63.3000 37.9000 ;
	    RECT 61.5000 37.5000 63.3000 37.8000 ;
	    RECT 61.5000 36.2000 61.8000 37.5000 ;
	    RECT 62.2000 36.4000 62.6000 37.2000 ;
	    RECT 61.4000 35.8000 61.8000 36.2000 ;
	    RECT 54.5000 35.6000 59.4000 35.7000 ;
	    RECT 56.5000 35.5000 59.4000 35.6000 ;
	    RECT 56.6000 35.4000 59.4000 35.5000 ;
	    RECT 51.1000 34.9000 51.5000 35.0000 ;
	    RECT 51.1000 34.6000 53.0000 34.9000 ;
	    RECT 53.4000 34.8000 53.8000 35.2000 ;
	    RECT 55.8000 35.1000 56.2000 35.2000 ;
	    RECT 55.8000 34.8000 58.3000 35.1000 ;
	    RECT 52.6000 34.5000 53.0000 34.6000 ;
	    RECT 53.5000 34.2000 53.8000 34.8000 ;
	    RECT 56.6000 34.7000 57.0000 34.8000 ;
	    RECT 57.9000 34.7000 58.3000 34.8000 ;
	    RECT 57.1000 34.2000 57.5000 34.3000 ;
	    RECT 61.5000 34.2000 61.8000 35.8000 ;
	    RECT 62.6000 34.8000 63.4000 35.2000 ;
	    RECT 63.8000 35.1000 64.2000 36.2000 ;
	    RECT 63.8000 34.8000 64.9000 35.1000 ;
	    RECT 64.6000 34.2000 64.9000 34.8000 ;
	    RECT 53.5000 33.9000 59.0000 34.2000 ;
	    RECT 61.5000 34.1000 62.3000 34.2000 ;
	    RECT 61.5000 33.9000 62.4000 34.1000 ;
	    RECT 53.7000 33.8000 54.1000 33.9000 ;
	    RECT 50.2000 33.3000 52.1000 33.6000 ;
	    RECT 50.2000 31.1000 50.6000 33.3000 ;
	    RECT 51.7000 33.2000 52.1000 33.3000 ;
	    RECT 56.6000 32.8000 56.9000 33.9000 ;
	    RECT 58.2000 33.8000 59.0000 33.9000 ;
	    RECT 55.7000 32.7000 56.1000 32.8000 ;
	    RECT 52.6000 32.1000 53.0000 32.5000 ;
	    RECT 54.7000 32.4000 56.1000 32.7000 ;
	    RECT 56.6000 32.4000 57.0000 32.8000 ;
	    RECT 54.7000 32.1000 55.0000 32.4000 ;
	    RECT 57.4000 32.1000 57.8000 32.5000 ;
	    RECT 52.3000 31.8000 53.0000 32.1000 ;
	    RECT 52.3000 31.1000 52.9000 31.8000 ;
	    RECT 54.6000 31.1000 55.0000 32.1000 ;
	    RECT 56.8000 31.8000 57.8000 32.1000 ;
	    RECT 56.8000 31.1000 57.2000 31.8000 ;
	    RECT 59.0000 31.1000 59.4000 33.5000 ;
	    RECT 62.0000 31.1000 62.4000 33.9000 ;
	    RECT 64.6000 33.4000 65.0000 34.2000 ;
	    RECT 65.4000 33.1000 65.8000 39.9000 ;
	    RECT 66.2000 35.8000 66.6000 36.6000 ;
	    RECT 67.8000 34.1000 68.2000 39.9000 ;
	    RECT 69.9000 39.2000 70.3000 39.9000 ;
	    RECT 69.4000 38.8000 70.3000 39.2000 ;
	    RECT 69.9000 36.2000 70.3000 38.8000 ;
	    RECT 70.6000 36.8000 71.0000 37.2000 ;
	    RECT 70.7000 36.2000 71.0000 36.8000 ;
	    RECT 69.9000 35.9000 70.4000 36.2000 ;
	    RECT 70.7000 35.9000 71.4000 36.2000 ;
	    RECT 69.4000 34.4000 69.8000 35.2000 ;
	    RECT 70.1000 34.2000 70.4000 35.9000 ;
	    RECT 71.0000 35.8000 71.4000 35.9000 ;
	    RECT 71.8000 35.6000 72.2000 39.9000 ;
	    RECT 73.9000 37.9000 74.5000 39.9000 ;
	    RECT 76.2000 37.9000 76.6000 39.9000 ;
	    RECT 78.4000 38.2000 78.8000 39.9000 ;
	    RECT 78.4000 37.9000 79.4000 38.2000 ;
	    RECT 74.2000 37.5000 74.6000 37.9000 ;
	    RECT 76.3000 37.6000 76.6000 37.9000 ;
	    RECT 75.9000 37.3000 77.7000 37.6000 ;
	    RECT 79.0000 37.5000 79.4000 37.9000 ;
	    RECT 75.9000 37.2000 76.3000 37.3000 ;
	    RECT 77.3000 37.2000 77.7000 37.3000 ;
	    RECT 73.8000 36.6000 74.5000 37.0000 ;
	    RECT 74.2000 36.1000 74.5000 36.6000 ;
	    RECT 75.3000 36.5000 76.4000 36.8000 ;
	    RECT 75.3000 36.4000 75.7000 36.5000 ;
	    RECT 74.2000 35.8000 75.4000 36.1000 ;
	    RECT 71.8000 35.3000 73.9000 35.6000 ;
	    RECT 68.6000 34.1000 69.0000 34.2000 ;
	    RECT 67.8000 33.8000 69.4000 34.1000 ;
	    RECT 70.1000 33.8000 71.4000 34.2000 ;
	    RECT 67.0000 33.1000 67.4000 33.2000 ;
	    RECT 65.4000 32.8000 67.4000 33.1000 ;
	    RECT 65.9000 31.1000 66.3000 32.8000 ;
	    RECT 67.0000 32.4000 67.4000 32.8000 ;
	    RECT 67.8000 31.1000 68.2000 33.8000 ;
	    RECT 69.0000 33.6000 69.4000 33.8000 ;
	    RECT 68.7000 33.1000 70.5000 33.3000 ;
	    RECT 71.0000 33.1000 71.3000 33.8000 ;
	    RECT 71.8000 33.6000 72.2000 35.3000 ;
	    RECT 73.5000 35.2000 73.9000 35.3000 ;
	    RECT 72.7000 34.9000 73.1000 35.0000 ;
	    RECT 72.7000 34.6000 74.6000 34.9000 ;
	    RECT 74.2000 34.5000 74.6000 34.6000 ;
	    RECT 75.1000 34.2000 75.4000 35.8000 ;
	    RECT 76.1000 35.9000 76.4000 36.5000 ;
	    RECT 76.7000 36.5000 77.1000 36.6000 ;
	    RECT 79.0000 36.5000 79.4000 36.6000 ;
	    RECT 76.7000 36.2000 79.4000 36.5000 ;
	    RECT 76.1000 35.7000 78.5000 35.9000 ;
	    RECT 80.6000 35.7000 81.0000 39.9000 ;
	    RECT 82.2000 37.9000 82.6000 39.9000 ;
	    RECT 82.3000 37.8000 82.6000 37.9000 ;
	    RECT 83.8000 37.9000 84.2000 39.9000 ;
	    RECT 85.4000 37.9000 85.8000 39.9000 ;
	    RECT 83.8000 37.8000 84.1000 37.9000 ;
	    RECT 82.3000 37.5000 84.1000 37.8000 ;
	    RECT 85.5000 37.8000 85.8000 37.9000 ;
	    RECT 87.0000 37.9000 87.4000 39.9000 ;
	    RECT 87.9000 39.6000 89.7000 39.9000 ;
	    RECT 87.9000 39.5000 88.2000 39.6000 ;
	    RECT 87.0000 37.8000 87.3000 37.9000 ;
	    RECT 85.5000 37.5000 87.3000 37.8000 ;
	    RECT 83.0000 36.4000 83.4000 37.2000 ;
	    RECT 83.8000 36.2000 84.1000 37.5000 ;
	    RECT 86.2000 36.4000 86.6000 37.2000 ;
	    RECT 87.0000 36.2000 87.3000 37.5000 ;
	    RECT 87.8000 36.5000 88.2000 39.5000 ;
	    RECT 89.4000 39.5000 89.7000 39.6000 ;
	    RECT 90.2000 39.6000 92.2000 39.9000 ;
	    RECT 88.6000 36.5000 89.0000 39.3000 ;
	    RECT 89.4000 36.7000 89.8000 39.5000 ;
	    RECT 90.2000 37.0000 90.6000 39.6000 ;
	    RECT 91.0000 36.9000 91.4000 39.3000 ;
	    RECT 91.8000 36.9000 92.2000 39.6000 ;
	    RECT 91.0000 36.7000 91.3000 36.9000 ;
	    RECT 89.4000 36.5000 91.3000 36.7000 ;
	    RECT 88.7000 36.2000 89.0000 36.5000 ;
	    RECT 89.5000 36.4000 91.3000 36.5000 ;
	    RECT 91.9000 36.6000 92.2000 36.9000 ;
	    RECT 93.4000 36.9000 93.8000 39.9000 ;
	    RECT 93.4000 36.6000 93.7000 36.9000 ;
	    RECT 91.9000 36.3000 93.7000 36.6000 ;
	    RECT 76.1000 35.6000 81.0000 35.7000 ;
	    RECT 78.1000 35.5000 81.0000 35.6000 ;
	    RECT 78.2000 35.4000 81.0000 35.5000 ;
	    RECT 77.4000 35.1000 77.8000 35.2000 ;
	    RECT 77.4000 34.8000 79.9000 35.1000 ;
	    RECT 81.4000 34.8000 81.8000 36.2000 ;
	    RECT 83.8000 35.8000 84.2000 36.2000 ;
	    RECT 82.2000 34.8000 83.0000 35.2000 ;
	    RECT 78.2000 34.7000 78.6000 34.8000 ;
	    RECT 79.5000 34.7000 79.9000 34.8000 ;
	    RECT 78.7000 34.2000 79.1000 34.3000 ;
	    RECT 83.8000 34.2000 84.1000 35.8000 ;
	    RECT 84.6000 34.8000 85.0000 36.2000 ;
	    RECT 87.0000 35.8000 87.4000 36.2000 ;
	    RECT 88.6000 36.1000 89.0000 36.2000 ;
	    RECT 94.2000 36.1000 94.6000 39.9000 ;
	    RECT 96.2000 36.8000 96.6000 37.2000 ;
	    RECT 96.2000 36.2000 96.5000 36.8000 ;
	    RECT 96.9000 36.2000 97.3000 39.9000 ;
	    RECT 95.8000 36.1000 96.5000 36.2000 ;
	    RECT 88.6000 35.8000 90.3000 36.1000 ;
	    RECT 85.4000 34.8000 86.2000 35.2000 ;
	    RECT 87.0000 34.2000 87.3000 35.8000 ;
	    RECT 75.1000 33.9000 80.6000 34.2000 ;
	    RECT 83.3000 34.1000 84.1000 34.2000 ;
	    RECT 86.5000 34.1000 87.3000 34.2000 ;
	    RECT 75.3000 33.8000 75.7000 33.9000 ;
	    RECT 71.8000 33.3000 73.7000 33.6000 ;
	    RECT 68.6000 33.0000 70.6000 33.1000 ;
	    RECT 68.6000 31.1000 69.0000 33.0000 ;
	    RECT 70.2000 31.1000 70.6000 33.0000 ;
	    RECT 71.0000 31.1000 71.4000 33.1000 ;
	    RECT 71.8000 31.1000 72.2000 33.3000 ;
	    RECT 73.3000 33.2000 73.7000 33.3000 ;
	    RECT 78.2000 33.2000 78.5000 33.9000 ;
	    RECT 79.8000 33.8000 80.6000 33.9000 ;
	    RECT 83.2000 33.9000 84.1000 34.1000 ;
	    RECT 86.4000 33.9000 87.3000 34.1000 ;
	    RECT 77.3000 32.7000 77.7000 32.8000 ;
	    RECT 74.2000 32.1000 74.6000 32.5000 ;
	    RECT 76.3000 32.4000 77.7000 32.7000 ;
	    RECT 78.2000 32.4000 78.6000 33.2000 ;
	    RECT 76.3000 32.1000 76.6000 32.4000 ;
	    RECT 79.0000 32.1000 79.4000 32.5000 ;
	    RECT 73.9000 31.8000 74.6000 32.1000 ;
	    RECT 73.9000 31.1000 74.5000 31.8000 ;
	    RECT 76.2000 31.1000 76.6000 32.1000 ;
	    RECT 78.4000 31.8000 79.4000 32.1000 ;
	    RECT 78.4000 31.1000 78.8000 31.8000 ;
	    RECT 80.6000 31.1000 81.0000 33.5000 ;
	    RECT 83.2000 31.1000 83.6000 33.9000 ;
	    RECT 86.4000 31.1000 86.8000 33.9000 ;
	    RECT 90.0000 32.5000 90.3000 35.8000 ;
	    RECT 94.2000 35.9000 96.5000 36.1000 ;
	    RECT 96.8000 35.9000 97.3000 36.2000 ;
	    RECT 100.3000 36.2000 100.7000 39.9000 ;
	    RECT 101.0000 36.8000 101.4000 37.2000 ;
	    RECT 101.1000 36.2000 101.4000 36.8000 ;
	    RECT 103.5000 36.2000 103.9000 39.9000 ;
	    RECT 104.2000 36.8000 104.6000 37.2000 ;
	    RECT 104.3000 36.2000 104.6000 36.8000 ;
	    RECT 100.3000 35.9000 100.8000 36.2000 ;
	    RECT 101.1000 35.9000 101.8000 36.2000 ;
	    RECT 103.5000 35.9000 104.0000 36.2000 ;
	    RECT 104.3000 36.1000 105.0000 36.2000 ;
	    RECT 106.2000 36.1000 106.6000 36.2000 ;
	    RECT 104.3000 35.9000 106.6000 36.1000 ;
	    RECT 94.2000 35.8000 96.2000 35.9000 ;
	    RECT 90.6000 34.8000 91.4000 35.2000 ;
	    RECT 91.4000 34.1000 92.2000 34.2000 ;
	    RECT 94.2000 34.1000 94.6000 35.8000 ;
	    RECT 96.8000 34.2000 97.1000 35.9000 ;
	    RECT 97.4000 34.4000 97.8000 35.2000 ;
	    RECT 99.8000 34.4000 100.2000 35.2000 ;
	    RECT 100.5000 34.2000 100.8000 35.9000 ;
	    RECT 101.4000 35.8000 101.8000 35.9000 ;
	    RECT 103.0000 34.4000 103.4000 35.2000 ;
	    RECT 103.7000 34.2000 104.0000 35.9000 ;
	    RECT 104.6000 35.8000 106.6000 35.9000 ;
	    RECT 107.0000 35.7000 107.4000 39.9000 ;
	    RECT 109.2000 38.2000 109.6000 39.9000 ;
	    RECT 108.6000 37.9000 109.6000 38.2000 ;
	    RECT 111.4000 37.9000 111.8000 39.9000 ;
	    RECT 113.5000 37.9000 114.1000 39.9000 ;
	    RECT 108.6000 37.5000 109.0000 37.9000 ;
	    RECT 111.4000 37.6000 111.7000 37.9000 ;
	    RECT 110.3000 37.3000 112.1000 37.6000 ;
	    RECT 113.4000 37.5000 113.8000 37.9000 ;
	    RECT 110.3000 37.2000 110.7000 37.3000 ;
	    RECT 111.7000 37.2000 112.1000 37.3000 ;
	    RECT 108.6000 36.5000 109.0000 36.6000 ;
	    RECT 110.9000 36.5000 111.3000 36.6000 ;
	    RECT 108.6000 36.2000 111.3000 36.5000 ;
	    RECT 111.6000 36.5000 112.7000 36.8000 ;
	    RECT 111.6000 35.9000 111.9000 36.5000 ;
	    RECT 112.3000 36.4000 112.7000 36.5000 ;
	    RECT 113.5000 36.6000 114.2000 37.0000 ;
	    RECT 113.5000 36.1000 113.8000 36.6000 ;
	    RECT 109.5000 35.7000 111.9000 35.9000 ;
	    RECT 107.0000 35.6000 111.9000 35.7000 ;
	    RECT 112.6000 35.8000 113.8000 36.1000 ;
	    RECT 107.0000 35.5000 109.9000 35.6000 ;
	    RECT 107.0000 35.4000 109.8000 35.5000 ;
	    RECT 112.6000 35.2000 112.9000 35.8000 ;
	    RECT 115.8000 35.6000 116.2000 39.9000 ;
	    RECT 117.9000 36.2000 118.3000 39.9000 ;
	    RECT 119.8000 39.6000 121.8000 39.9000 ;
	    RECT 118.6000 36.8000 119.0000 37.2000 ;
	    RECT 118.7000 36.2000 119.0000 36.8000 ;
	    RECT 117.9000 35.9000 118.4000 36.2000 ;
	    RECT 118.7000 35.9000 119.4000 36.2000 ;
	    RECT 119.8000 35.9000 120.2000 39.6000 ;
	    RECT 120.6000 35.9000 121.0000 39.3000 ;
	    RECT 121.4000 36.2000 121.8000 39.6000 ;
	    RECT 123.0000 36.2000 123.4000 39.9000 ;
	    RECT 124.6000 37.9000 125.0000 39.9000 ;
	    RECT 124.7000 37.8000 125.0000 37.9000 ;
	    RECT 126.2000 37.9000 126.6000 39.9000 ;
	    RECT 126.2000 37.8000 126.5000 37.9000 ;
	    RECT 124.7000 37.5000 126.5000 37.8000 ;
	    RECT 123.8000 37.1000 124.2000 37.2000 ;
	    RECT 125.4000 37.1000 125.8000 37.2000 ;
	    RECT 123.8000 36.8000 125.8000 37.1000 ;
	    RECT 125.4000 36.4000 125.8000 36.8000 ;
	    RECT 126.2000 36.2000 126.5000 37.5000 ;
	    RECT 121.4000 35.9000 123.4000 36.2000 ;
	    RECT 114.1000 35.3000 116.2000 35.6000 ;
	    RECT 114.1000 35.2000 114.5000 35.3000 ;
	    RECT 110.2000 35.1000 110.6000 35.2000 ;
	    RECT 108.1000 34.8000 110.6000 35.1000 ;
	    RECT 112.6000 34.8000 113.0000 35.2000 ;
	    RECT 114.9000 34.9000 115.3000 35.0000 ;
	    RECT 108.1000 34.7000 108.5000 34.8000 ;
	    RECT 109.4000 34.7000 109.8000 34.8000 ;
	    RECT 108.9000 34.2000 109.3000 34.3000 ;
	    RECT 112.6000 34.2000 112.9000 34.8000 ;
	    RECT 113.4000 34.6000 115.3000 34.9000 ;
	    RECT 113.4000 34.5000 113.8000 34.6000 ;
	    RECT 91.4000 33.8000 94.6000 34.1000 ;
	    RECT 95.8000 33.8000 97.1000 34.2000 ;
	    RECT 98.2000 34.1000 98.6000 34.2000 ;
	    RECT 97.8000 33.8000 98.6000 34.1000 ;
	    RECT 99.0000 34.1000 99.4000 34.2000 ;
	    RECT 99.0000 33.8000 99.8000 34.1000 ;
	    RECT 100.5000 33.8000 101.8000 34.2000 ;
	    RECT 102.2000 34.1000 102.6000 34.2000 ;
	    RECT 102.2000 33.8000 103.0000 34.1000 ;
	    RECT 103.7000 33.8000 105.0000 34.2000 ;
	    RECT 107.4000 33.9000 112.9000 34.2000 ;
	    RECT 107.4000 33.8000 108.2000 33.9000 ;
	    RECT 92.1000 32.8000 93.0000 33.2000 ;
	    RECT 90.0000 32.2000 92.0000 32.5000 ;
	    RECT 90.0000 32.1000 90.6000 32.2000 ;
	    RECT 90.2000 31.1000 90.6000 32.1000 ;
	    RECT 91.7000 31.8000 92.2000 32.2000 ;
	    RECT 91.8000 31.1000 92.2000 31.8000 ;
	    RECT 94.2000 31.1000 94.6000 33.8000 ;
	    RECT 95.0000 32.4000 95.4000 33.2000 ;
	    RECT 95.9000 33.1000 96.2000 33.8000 ;
	    RECT 97.8000 33.6000 98.2000 33.8000 ;
	    RECT 99.4000 33.6000 99.8000 33.8000 ;
	    RECT 96.7000 33.1000 98.5000 33.3000 ;
	    RECT 99.1000 33.1000 100.9000 33.3000 ;
	    RECT 101.4000 33.1000 101.7000 33.8000 ;
	    RECT 102.6000 33.6000 103.0000 33.8000 ;
	    RECT 102.3000 33.1000 104.1000 33.3000 ;
	    RECT 104.6000 33.1000 104.9000 33.8000 ;
	    RECT 95.8000 31.1000 96.2000 33.1000 ;
	    RECT 96.6000 33.0000 98.6000 33.1000 ;
	    RECT 96.6000 31.1000 97.0000 33.0000 ;
	    RECT 98.2000 31.1000 98.6000 33.0000 ;
	    RECT 99.0000 33.0000 101.0000 33.1000 ;
	    RECT 99.0000 31.1000 99.4000 33.0000 ;
	    RECT 100.6000 31.1000 101.0000 33.0000 ;
	    RECT 101.4000 31.1000 101.8000 33.1000 ;
	    RECT 102.2000 33.0000 104.2000 33.1000 ;
	    RECT 102.2000 31.1000 102.6000 33.0000 ;
	    RECT 103.8000 31.1000 104.2000 33.0000 ;
	    RECT 104.6000 32.1000 105.0000 33.1000 ;
	    RECT 106.2000 32.1000 106.6000 32.2000 ;
	    RECT 104.6000 31.8000 106.6000 32.1000 ;
	    RECT 104.6000 31.1000 105.0000 31.8000 ;
	    RECT 107.0000 31.1000 107.4000 33.5000 ;
	    RECT 109.5000 32.8000 109.8000 33.9000 ;
	    RECT 112.3000 33.8000 112.7000 33.9000 ;
	    RECT 115.8000 33.6000 116.2000 35.3000 ;
	    RECT 117.4000 34.4000 117.8000 35.2000 ;
	    RECT 118.1000 34.2000 118.4000 35.9000 ;
	    RECT 119.0000 35.8000 119.4000 35.9000 ;
	    RECT 120.7000 35.6000 121.0000 35.9000 ;
	    RECT 119.8000 34.8000 120.2000 35.6000 ;
	    RECT 120.7000 35.3000 121.7000 35.6000 ;
	    RECT 123.8000 35.4000 124.2000 36.2000 ;
	    RECT 126.2000 35.8000 126.6000 36.2000 ;
	    RECT 121.4000 35.2000 121.7000 35.3000 ;
	    RECT 122.6000 35.2000 123.0000 35.4000 ;
	    RECT 121.4000 34.8000 121.8000 35.2000 ;
	    RECT 122.6000 34.9000 123.4000 35.2000 ;
	    RECT 123.0000 34.8000 123.4000 34.9000 ;
	    RECT 124.6000 34.8000 125.4000 35.2000 ;
	    RECT 120.7000 34.4000 121.1000 34.8000 ;
	    RECT 120.7000 34.2000 121.0000 34.4000 ;
	    RECT 116.6000 34.1000 117.0000 34.2000 ;
	    RECT 118.1000 34.1000 119.4000 34.2000 ;
	    RECT 119.8000 34.1000 120.2000 34.2000 ;
	    RECT 116.6000 33.8000 117.4000 34.1000 ;
	    RECT 118.1000 33.8000 120.2000 34.1000 ;
	    RECT 120.6000 33.8000 121.0000 34.2000 ;
	    RECT 117.0000 33.6000 117.4000 33.8000 ;
	    RECT 114.3000 33.3000 116.2000 33.6000 ;
	    RECT 114.3000 33.2000 114.7000 33.3000 ;
	    RECT 108.6000 32.1000 109.0000 32.5000 ;
	    RECT 109.4000 32.4000 109.8000 32.8000 ;
	    RECT 110.3000 32.7000 110.7000 32.8000 ;
	    RECT 110.3000 32.4000 111.7000 32.7000 ;
	    RECT 111.4000 32.1000 111.7000 32.4000 ;
	    RECT 113.4000 32.1000 113.8000 32.5000 ;
	    RECT 108.6000 31.8000 109.6000 32.1000 ;
	    RECT 109.2000 31.1000 109.6000 31.8000 ;
	    RECT 111.4000 31.1000 111.8000 32.1000 ;
	    RECT 113.4000 31.8000 114.1000 32.1000 ;
	    RECT 113.5000 31.1000 114.1000 31.8000 ;
	    RECT 115.8000 31.1000 116.2000 33.3000 ;
	    RECT 116.7000 33.1000 118.5000 33.3000 ;
	    RECT 119.0000 33.1000 119.3000 33.8000 ;
	    RECT 121.4000 33.1000 121.7000 34.8000 ;
	    RECT 122.2000 33.8000 122.6000 34.6000 ;
	    RECT 126.2000 34.2000 126.5000 35.8000 ;
	    RECT 127.0000 35.7000 127.4000 39.9000 ;
	    RECT 129.2000 38.2000 129.6000 39.9000 ;
	    RECT 128.6000 37.9000 129.6000 38.2000 ;
	    RECT 131.4000 37.9000 131.8000 39.9000 ;
	    RECT 133.5000 37.9000 134.1000 39.9000 ;
	    RECT 128.6000 37.5000 129.0000 37.9000 ;
	    RECT 131.4000 37.6000 131.7000 37.9000 ;
	    RECT 130.3000 37.3000 132.1000 37.6000 ;
	    RECT 133.4000 37.5000 133.8000 37.9000 ;
	    RECT 130.3000 37.2000 130.7000 37.3000 ;
	    RECT 131.7000 37.2000 132.1000 37.3000 ;
	    RECT 128.6000 36.5000 129.0000 36.6000 ;
	    RECT 130.9000 36.5000 131.3000 36.6000 ;
	    RECT 128.6000 36.2000 131.3000 36.5000 ;
	    RECT 131.6000 36.5000 132.7000 36.8000 ;
	    RECT 131.6000 35.9000 131.9000 36.5000 ;
	    RECT 132.3000 36.4000 132.7000 36.5000 ;
	    RECT 133.5000 36.6000 134.2000 37.0000 ;
	    RECT 133.5000 36.1000 133.8000 36.6000 ;
	    RECT 129.5000 35.7000 131.9000 35.9000 ;
	    RECT 127.0000 35.6000 131.9000 35.7000 ;
	    RECT 132.6000 35.8000 133.8000 36.1000 ;
	    RECT 127.0000 35.5000 129.9000 35.6000 ;
	    RECT 127.0000 35.4000 129.8000 35.5000 ;
	    RECT 132.6000 35.2000 132.9000 35.8000 ;
	    RECT 135.8000 35.6000 136.2000 39.9000 ;
	    RECT 137.4000 37.9000 137.8000 39.9000 ;
	    RECT 134.1000 35.3000 136.2000 35.6000 ;
	    RECT 137.5000 35.8000 137.8000 37.9000 ;
	    RECT 139.0000 35.9000 139.4000 39.9000 ;
	    RECT 140.1000 36.2000 140.5000 39.9000 ;
	    RECT 137.5000 35.5000 138.7000 35.8000 ;
	    RECT 134.1000 35.2000 134.5000 35.3000 ;
	    RECT 130.2000 35.1000 130.6000 35.2000 ;
	    RECT 128.1000 34.8000 130.6000 35.1000 ;
	    RECT 132.6000 34.8000 133.0000 35.2000 ;
	    RECT 134.9000 34.9000 135.3000 35.0000 ;
	    RECT 128.1000 34.7000 128.5000 34.8000 ;
	    RECT 129.4000 34.7000 129.8000 34.8000 ;
	    RECT 128.9000 34.2000 129.3000 34.3000 ;
	    RECT 132.6000 34.2000 132.9000 34.8000 ;
	    RECT 133.4000 34.6000 135.3000 34.9000 ;
	    RECT 133.4000 34.5000 133.8000 34.6000 ;
	    RECT 125.7000 34.1000 126.5000 34.2000 ;
	    RECT 125.6000 33.9000 126.5000 34.1000 ;
	    RECT 127.4000 33.9000 132.9000 34.2000 ;
	    RECT 116.6000 33.0000 118.6000 33.1000 ;
	    RECT 116.6000 31.1000 117.0000 33.0000 ;
	    RECT 118.2000 31.1000 118.6000 33.0000 ;
	    RECT 119.0000 31.1000 119.4000 33.1000 ;
	    RECT 121.1000 31.1000 121.9000 33.1000 ;
	    RECT 125.6000 31.1000 126.0000 33.9000 ;
	    RECT 127.4000 33.8000 128.2000 33.9000 ;
	    RECT 127.0000 31.1000 127.4000 33.5000 ;
	    RECT 129.5000 32.8000 129.8000 33.9000 ;
	    RECT 132.3000 33.8000 132.7000 33.9000 ;
	    RECT 135.8000 33.6000 136.2000 35.3000 ;
	    RECT 137.4000 34.8000 137.8000 35.2000 ;
	    RECT 136.6000 33.8000 137.0000 34.6000 ;
	    RECT 137.5000 34.4000 137.8000 34.8000 ;
	    RECT 137.5000 34.1000 138.0000 34.4000 ;
	    RECT 137.6000 34.0000 138.0000 34.1000 ;
	    RECT 138.4000 33.8000 138.7000 35.5000 ;
	    RECT 139.1000 35.2000 139.4000 35.9000 ;
	    RECT 139.0000 34.8000 139.4000 35.2000 ;
	    RECT 138.4000 33.7000 138.8000 33.8000 ;
	    RECT 134.3000 33.3000 136.2000 33.6000 ;
	    RECT 137.3000 33.5000 138.8000 33.7000 ;
	    RECT 134.3000 33.2000 134.7000 33.3000 ;
	    RECT 128.6000 32.1000 129.0000 32.5000 ;
	    RECT 129.4000 32.4000 129.8000 32.8000 ;
	    RECT 130.3000 32.7000 130.7000 32.8000 ;
	    RECT 130.3000 32.4000 131.7000 32.7000 ;
	    RECT 131.4000 32.1000 131.7000 32.4000 ;
	    RECT 133.4000 32.1000 133.8000 32.5000 ;
	    RECT 128.6000 31.8000 129.6000 32.1000 ;
	    RECT 129.2000 31.1000 129.6000 31.8000 ;
	    RECT 131.4000 31.1000 131.8000 32.1000 ;
	    RECT 133.4000 31.8000 134.1000 32.1000 ;
	    RECT 133.5000 31.1000 134.1000 31.8000 ;
	    RECT 135.8000 31.1000 136.2000 33.3000 ;
	    RECT 136.7000 33.4000 138.8000 33.5000 ;
	    RECT 136.7000 33.2000 137.6000 33.4000 ;
	    RECT 136.7000 33.1000 137.0000 33.2000 ;
	    RECT 139.1000 33.1000 139.4000 34.8000 ;
	    RECT 136.6000 31.1000 137.0000 33.1000 ;
	    RECT 138.7000 32.6000 139.4000 33.1000 ;
	    RECT 139.8000 35.9000 140.5000 36.2000 ;
	    RECT 139.8000 35.2000 140.1000 35.9000 ;
	    RECT 142.2000 35.6000 142.6000 39.9000 ;
	    RECT 140.6000 35.4000 142.6000 35.6000 ;
	    RECT 143.0000 35.7000 143.4000 39.9000 ;
	    RECT 145.2000 38.2000 145.6000 39.9000 ;
	    RECT 144.6000 37.9000 145.6000 38.2000 ;
	    RECT 147.4000 37.9000 147.8000 39.9000 ;
	    RECT 149.5000 37.9000 150.1000 39.9000 ;
	    RECT 144.6000 37.5000 145.0000 37.9000 ;
	    RECT 147.4000 37.6000 147.7000 37.9000 ;
	    RECT 146.3000 37.3000 148.1000 37.6000 ;
	    RECT 149.4000 37.5000 149.8000 37.9000 ;
	    RECT 146.3000 37.2000 146.7000 37.3000 ;
	    RECT 147.7000 37.2000 148.1000 37.3000 ;
	    RECT 144.6000 36.5000 145.0000 36.6000 ;
	    RECT 146.9000 36.5000 147.3000 36.6000 ;
	    RECT 144.6000 36.2000 147.3000 36.5000 ;
	    RECT 147.6000 36.5000 148.7000 36.8000 ;
	    RECT 147.6000 35.9000 147.9000 36.5000 ;
	    RECT 148.3000 36.4000 148.7000 36.5000 ;
	    RECT 149.5000 36.6000 150.2000 37.0000 ;
	    RECT 149.5000 36.1000 149.8000 36.6000 ;
	    RECT 145.5000 35.7000 147.9000 35.9000 ;
	    RECT 143.0000 35.6000 147.9000 35.7000 ;
	    RECT 148.6000 35.8000 149.8000 36.1000 ;
	    RECT 143.0000 35.5000 145.9000 35.6000 ;
	    RECT 143.0000 35.4000 145.8000 35.5000 ;
	    RECT 140.5000 35.3000 142.6000 35.4000 ;
	    RECT 139.8000 34.8000 140.2000 35.2000 ;
	    RECT 140.5000 35.0000 140.9000 35.3000 ;
	    RECT 146.2000 35.1000 146.6000 35.2000 ;
	    RECT 139.8000 33.1000 140.1000 34.8000 ;
	    RECT 140.5000 33.5000 140.8000 35.0000 ;
	    RECT 144.1000 34.8000 146.6000 35.1000 ;
	    RECT 144.1000 34.7000 144.5000 34.8000 ;
	    RECT 145.4000 34.7000 145.8000 34.8000 ;
	    RECT 141.2000 34.2000 141.6000 34.6000 ;
	    RECT 144.9000 34.2000 145.3000 34.3000 ;
	    RECT 148.6000 34.2000 148.9000 35.8000 ;
	    RECT 151.8000 35.6000 152.2000 39.9000 ;
	    RECT 150.1000 35.3000 152.2000 35.6000 ;
	    RECT 150.1000 35.2000 150.5000 35.3000 ;
	    RECT 150.9000 34.9000 151.3000 35.0000 ;
	    RECT 149.4000 34.6000 151.3000 34.9000 ;
	    RECT 149.4000 34.5000 149.8000 34.6000 ;
	    RECT 141.3000 33.8000 141.8000 34.2000 ;
	    RECT 143.4000 33.9000 148.9000 34.2000 ;
	    RECT 143.4000 33.8000 144.2000 33.9000 ;
	    RECT 140.5000 33.2000 141.7000 33.5000 ;
	    RECT 138.7000 31.1000 139.1000 32.6000 ;
	    RECT 139.8000 31.1000 140.2000 33.1000 ;
	    RECT 141.4000 32.1000 141.7000 33.2000 ;
	    RECT 142.2000 32.4000 142.6000 33.2000 ;
	    RECT 141.4000 31.1000 141.8000 32.1000 ;
	    RECT 143.0000 31.1000 143.4000 33.5000 ;
	    RECT 145.5000 33.2000 145.8000 33.9000 ;
	    RECT 148.3000 33.8000 148.7000 33.9000 ;
	    RECT 151.8000 33.6000 152.2000 35.3000 ;
	    RECT 150.3000 33.3000 152.2000 33.6000 ;
	    RECT 152.6000 33.4000 153.0000 34.2000 ;
	    RECT 153.4000 34.1000 153.8000 39.9000 ;
	    RECT 154.2000 35.8000 154.6000 36.6000 ;
	    RECT 155.0000 34.1000 155.4000 34.2000 ;
	    RECT 153.4000 33.8000 155.4000 34.1000 ;
	    RECT 150.3000 33.2000 150.7000 33.3000 ;
	    RECT 144.6000 32.1000 145.0000 32.5000 ;
	    RECT 145.4000 32.4000 145.8000 33.2000 ;
	    RECT 146.3000 32.7000 146.7000 32.8000 ;
	    RECT 146.3000 32.4000 147.7000 32.7000 ;
	    RECT 147.4000 32.1000 147.7000 32.4000 ;
	    RECT 149.4000 32.1000 149.8000 32.5000 ;
	    RECT 144.6000 31.8000 145.6000 32.1000 ;
	    RECT 145.2000 31.1000 145.6000 31.8000 ;
	    RECT 147.4000 31.1000 147.8000 32.1000 ;
	    RECT 149.4000 31.8000 150.1000 32.1000 ;
	    RECT 149.5000 31.1000 150.1000 31.8000 ;
	    RECT 151.8000 31.1000 152.2000 33.3000 ;
	    RECT 153.4000 33.1000 153.8000 33.8000 ;
	    RECT 155.0000 33.4000 155.4000 33.8000 ;
	    RECT 155.8000 33.1000 156.2000 39.9000 ;
	    RECT 156.6000 35.8000 157.0000 36.6000 ;
	    RECT 153.4000 32.8000 154.3000 33.1000 ;
	    RECT 155.8000 32.8000 156.7000 33.1000 ;
	    RECT 153.9000 31.1000 154.3000 32.8000 ;
	    RECT 156.3000 32.2000 156.7000 32.8000 ;
	    RECT 155.8000 31.8000 156.7000 32.2000 ;
	    RECT 156.3000 31.1000 156.7000 31.8000 ;
	    RECT 157.4000 31.1000 157.8000 39.9000 ;
	    RECT 160.6000 35.6000 161.0000 39.9000 ;
	    RECT 162.7000 37.9000 163.3000 39.9000 ;
	    RECT 165.0000 37.9000 165.4000 39.9000 ;
	    RECT 167.2000 38.2000 167.6000 39.9000 ;
	    RECT 167.2000 37.9000 168.2000 38.2000 ;
	    RECT 163.0000 37.5000 163.4000 37.9000 ;
	    RECT 165.1000 37.6000 165.4000 37.9000 ;
	    RECT 164.7000 37.3000 166.5000 37.6000 ;
	    RECT 167.8000 37.5000 168.2000 37.9000 ;
	    RECT 164.7000 37.2000 165.1000 37.3000 ;
	    RECT 166.1000 37.2000 166.5000 37.3000 ;
	    RECT 162.6000 36.6000 163.3000 37.0000 ;
	    RECT 163.0000 36.1000 163.3000 36.6000 ;
	    RECT 164.1000 36.5000 165.2000 36.8000 ;
	    RECT 164.1000 36.4000 164.5000 36.5000 ;
	    RECT 163.0000 35.8000 164.2000 36.1000 ;
	    RECT 160.6000 35.3000 162.7000 35.6000 ;
	    RECT 160.6000 33.6000 161.0000 35.3000 ;
	    RECT 162.3000 35.2000 162.7000 35.3000 ;
	    RECT 163.9000 35.2000 164.2000 35.8000 ;
	    RECT 164.9000 35.9000 165.2000 36.5000 ;
	    RECT 165.5000 36.5000 165.9000 36.6000 ;
	    RECT 167.8000 36.5000 168.2000 36.6000 ;
	    RECT 165.5000 36.2000 168.2000 36.5000 ;
	    RECT 164.9000 35.7000 167.3000 35.9000 ;
	    RECT 169.4000 35.7000 169.8000 39.9000 ;
	    RECT 164.9000 35.6000 169.8000 35.7000 ;
	    RECT 166.9000 35.5000 169.8000 35.6000 ;
	    RECT 167.0000 35.4000 169.8000 35.5000 ;
	    RECT 161.5000 34.9000 161.9000 35.0000 ;
	    RECT 161.5000 34.6000 163.4000 34.9000 ;
	    RECT 163.8000 34.8000 164.2000 35.2000 ;
	    RECT 166.2000 35.1000 166.6000 35.2000 ;
	    RECT 166.2000 34.8000 168.7000 35.1000 ;
	    RECT 163.0000 34.5000 163.4000 34.6000 ;
	    RECT 163.9000 34.2000 164.2000 34.8000 ;
	    RECT 167.0000 34.7000 167.4000 34.8000 ;
	    RECT 168.3000 34.7000 168.7000 34.8000 ;
	    RECT 167.5000 34.2000 167.9000 34.3000 ;
	    RECT 163.9000 33.9000 169.4000 34.2000 ;
	    RECT 164.1000 33.8000 164.5000 33.9000 ;
	    RECT 160.6000 33.3000 162.5000 33.6000 ;
	    RECT 158.2000 32.4000 158.6000 33.2000 ;
	    RECT 160.6000 31.1000 161.0000 33.3000 ;
	    RECT 162.1000 33.2000 162.5000 33.3000 ;
	    RECT 167.0000 32.8000 167.3000 33.9000 ;
	    RECT 168.6000 33.8000 169.4000 33.9000 ;
	    RECT 166.1000 32.7000 166.5000 32.8000 ;
	    RECT 163.0000 32.1000 163.4000 32.5000 ;
	    RECT 165.1000 32.4000 166.5000 32.7000 ;
	    RECT 167.0000 32.4000 167.4000 32.8000 ;
	    RECT 165.1000 32.1000 165.4000 32.4000 ;
	    RECT 167.8000 32.1000 168.2000 32.5000 ;
	    RECT 162.7000 31.8000 163.4000 32.1000 ;
	    RECT 162.7000 31.1000 163.3000 31.8000 ;
	    RECT 165.0000 31.1000 165.4000 32.1000 ;
	    RECT 167.2000 31.8000 168.2000 32.1000 ;
	    RECT 167.2000 31.1000 167.6000 31.8000 ;
	    RECT 169.4000 31.1000 169.8000 33.5000 ;
	    RECT 170.2000 32.4000 170.6000 33.2000 ;
	    RECT 171.0000 33.1000 171.4000 39.9000 ;
	    RECT 173.1000 36.3000 173.5000 39.9000 ;
	    RECT 172.6000 35.9000 173.5000 36.3000 ;
	    RECT 172.7000 35.1000 173.0000 35.9000 ;
	    RECT 171.8000 34.8000 173.0000 35.1000 ;
	    RECT 173.4000 34.8000 173.8000 35.6000 ;
	    RECT 171.8000 34.2000 172.1000 34.8000 ;
	    RECT 172.7000 34.2000 173.0000 34.8000 ;
	    RECT 171.8000 33.8000 172.2000 34.2000 ;
	    RECT 172.6000 33.8000 173.0000 34.2000 ;
	    RECT 171.8000 33.1000 172.2000 33.2000 ;
	    RECT 171.0000 32.8000 172.2000 33.1000 ;
	    RECT 171.0000 31.1000 171.4000 32.8000 ;
	    RECT 171.8000 32.4000 172.2000 32.8000 ;
	    RECT 172.7000 32.1000 173.0000 33.8000 ;
	    RECT 172.6000 31.1000 173.0000 32.1000 ;
	    RECT 174.2000 31.1000 174.6000 39.9000 ;
	    RECT 175.8000 36.2000 176.2000 39.9000 ;
	    RECT 177.4000 36.4000 177.8000 39.9000 ;
	    RECT 175.8000 35.9000 177.1000 36.2000 ;
	    RECT 177.4000 35.9000 177.9000 36.4000 ;
	    RECT 175.8000 34.8000 176.3000 35.2000 ;
	    RECT 175.9000 34.4000 176.3000 34.8000 ;
	    RECT 176.8000 34.9000 177.1000 35.9000 ;
	    RECT 176.8000 34.5000 177.3000 34.9000 ;
	    RECT 176.8000 33.7000 177.1000 34.5000 ;
	    RECT 177.6000 34.2000 177.9000 35.9000 ;
	    RECT 179.0000 35.7000 179.4000 39.9000 ;
	    RECT 181.2000 38.2000 181.6000 39.9000 ;
	    RECT 180.6000 37.9000 181.6000 38.2000 ;
	    RECT 183.4000 37.9000 183.8000 39.9000 ;
	    RECT 185.5000 37.9000 186.1000 39.9000 ;
	    RECT 180.6000 37.5000 181.0000 37.9000 ;
	    RECT 183.4000 37.6000 183.7000 37.9000 ;
	    RECT 182.3000 37.3000 184.1000 37.6000 ;
	    RECT 185.4000 37.5000 185.8000 37.9000 ;
	    RECT 182.3000 37.2000 182.7000 37.3000 ;
	    RECT 183.7000 37.2000 184.1000 37.3000 ;
	    RECT 180.6000 36.5000 181.0000 36.6000 ;
	    RECT 182.9000 36.5000 183.3000 36.6000 ;
	    RECT 180.6000 36.2000 183.3000 36.5000 ;
	    RECT 183.6000 36.5000 184.7000 36.8000 ;
	    RECT 183.6000 35.9000 183.9000 36.5000 ;
	    RECT 184.3000 36.4000 184.7000 36.5000 ;
	    RECT 185.5000 36.6000 186.2000 37.0000 ;
	    RECT 185.5000 36.1000 185.8000 36.6000 ;
	    RECT 181.5000 35.7000 183.9000 35.9000 ;
	    RECT 179.0000 35.6000 183.9000 35.7000 ;
	    RECT 184.6000 35.8000 185.8000 36.1000 ;
	    RECT 179.0000 35.5000 181.9000 35.6000 ;
	    RECT 179.0000 35.4000 181.8000 35.5000 ;
	    RECT 182.2000 35.1000 182.6000 35.2000 ;
	    RECT 180.1000 34.8000 182.6000 35.1000 ;
	    RECT 180.1000 34.7000 180.5000 34.8000 ;
	    RECT 181.4000 34.7000 181.8000 34.8000 ;
	    RECT 180.9000 34.2000 181.3000 34.3000 ;
	    RECT 184.6000 34.2000 184.9000 35.8000 ;
	    RECT 187.8000 35.6000 188.2000 39.9000 ;
	    RECT 188.6000 36.2000 189.0000 39.9000 ;
	    RECT 190.2000 36.2000 190.6000 39.9000 ;
	    RECT 188.6000 35.9000 190.6000 36.2000 ;
	    RECT 191.0000 35.9000 191.4000 39.9000 ;
	    RECT 193.1000 36.2000 193.5000 39.9000 ;
	    RECT 193.8000 36.8000 194.2000 37.2000 ;
	    RECT 193.9000 36.2000 194.2000 36.8000 ;
	    RECT 193.1000 35.9000 193.6000 36.2000 ;
	    RECT 193.9000 35.9000 194.6000 36.2000 ;
	    RECT 186.1000 35.3000 188.2000 35.6000 ;
	    RECT 186.1000 35.2000 186.5000 35.3000 ;
	    RECT 186.9000 34.9000 187.3000 35.0000 ;
	    RECT 185.4000 34.6000 187.3000 34.9000 ;
	    RECT 185.4000 34.5000 185.8000 34.6000 ;
	    RECT 177.4000 33.8000 177.9000 34.2000 ;
	    RECT 179.4000 33.9000 184.9000 34.2000 ;
	    RECT 179.4000 33.8000 180.2000 33.9000 ;
	    RECT 175.8000 33.4000 177.1000 33.7000 ;
	    RECT 175.0000 32.4000 175.4000 33.2000 ;
	    RECT 175.8000 31.1000 176.2000 33.4000 ;
	    RECT 177.6000 33.1000 177.9000 33.8000 ;
	    RECT 177.4000 32.8000 177.9000 33.1000 ;
	    RECT 177.4000 31.1000 177.8000 32.8000 ;
	    RECT 179.0000 31.1000 179.4000 33.5000 ;
	    RECT 181.5000 32.8000 181.8000 33.9000 ;
	    RECT 184.3000 33.8000 184.7000 33.9000 ;
	    RECT 187.8000 33.6000 188.2000 35.3000 ;
	    RECT 189.0000 35.2000 189.4000 35.4000 ;
	    RECT 191.0000 35.2000 191.3000 35.9000 ;
	    RECT 188.6000 34.9000 189.4000 35.2000 ;
	    RECT 190.2000 34.9000 191.4000 35.2000 ;
	    RECT 188.6000 34.8000 189.0000 34.9000 ;
	    RECT 189.4000 33.8000 189.8000 34.6000 ;
	    RECT 186.3000 33.3000 188.2000 33.6000 ;
	    RECT 186.3000 33.2000 186.7000 33.3000 ;
	    RECT 180.6000 32.1000 181.0000 32.5000 ;
	    RECT 181.4000 32.4000 181.8000 32.8000 ;
	    RECT 182.3000 32.7000 182.7000 32.8000 ;
	    RECT 182.3000 32.4000 183.7000 32.7000 ;
	    RECT 183.4000 32.1000 183.7000 32.4000 ;
	    RECT 185.4000 32.1000 185.8000 32.5000 ;
	    RECT 180.6000 31.8000 181.6000 32.1000 ;
	    RECT 181.2000 31.1000 181.6000 31.8000 ;
	    RECT 183.4000 31.1000 183.8000 32.1000 ;
	    RECT 185.4000 31.8000 186.1000 32.1000 ;
	    RECT 185.5000 31.1000 186.1000 31.8000 ;
	    RECT 187.8000 31.1000 188.2000 33.3000 ;
	    RECT 190.2000 33.1000 190.5000 34.9000 ;
	    RECT 191.0000 34.8000 191.4000 34.9000 ;
	    RECT 191.8000 35.1000 192.2000 35.2000 ;
	    RECT 192.6000 35.1000 193.0000 35.2000 ;
	    RECT 191.8000 34.8000 193.0000 35.1000 ;
	    RECT 192.6000 34.4000 193.0000 34.8000 ;
	    RECT 193.3000 34.2000 193.6000 35.9000 ;
	    RECT 194.2000 35.8000 194.6000 35.9000 ;
	    RECT 195.0000 35.7000 195.4000 39.9000 ;
	    RECT 197.2000 38.2000 197.6000 39.9000 ;
	    RECT 196.6000 37.9000 197.6000 38.2000 ;
	    RECT 199.4000 37.9000 199.8000 39.9000 ;
	    RECT 201.5000 37.9000 202.1000 39.9000 ;
	    RECT 196.6000 37.5000 197.0000 37.9000 ;
	    RECT 199.4000 37.6000 199.7000 37.9000 ;
	    RECT 198.3000 37.3000 200.1000 37.6000 ;
	    RECT 201.4000 37.5000 201.8000 37.9000 ;
	    RECT 198.3000 37.2000 198.7000 37.3000 ;
	    RECT 199.7000 37.2000 200.1000 37.3000 ;
	    RECT 196.6000 36.5000 197.0000 36.6000 ;
	    RECT 198.9000 36.5000 199.3000 36.6000 ;
	    RECT 196.6000 36.2000 199.3000 36.5000 ;
	    RECT 199.6000 36.5000 200.7000 36.8000 ;
	    RECT 199.6000 35.9000 199.9000 36.5000 ;
	    RECT 200.3000 36.4000 200.7000 36.5000 ;
	    RECT 201.5000 36.6000 202.2000 37.0000 ;
	    RECT 201.5000 36.1000 201.8000 36.6000 ;
	    RECT 197.5000 35.7000 199.9000 35.9000 ;
	    RECT 195.0000 35.6000 199.9000 35.7000 ;
	    RECT 200.6000 35.8000 201.8000 36.1000 ;
	    RECT 195.0000 35.5000 197.9000 35.6000 ;
	    RECT 195.0000 35.4000 197.8000 35.5000 ;
	    RECT 198.2000 35.1000 198.6000 35.2000 ;
	    RECT 196.1000 34.8000 198.6000 35.1000 ;
	    RECT 196.1000 34.7000 196.5000 34.8000 ;
	    RECT 197.4000 34.7000 197.8000 34.8000 ;
	    RECT 196.9000 34.2000 197.3000 34.3000 ;
	    RECT 200.6000 34.2000 200.9000 35.8000 ;
	    RECT 203.8000 35.6000 204.2000 39.9000 ;
	    RECT 205.4000 37.9000 205.8000 39.9000 ;
	    RECT 202.1000 35.3000 204.2000 35.6000 ;
	    RECT 205.5000 35.8000 205.8000 37.9000 ;
	    RECT 207.0000 35.9000 207.4000 39.9000 ;
	    RECT 205.5000 35.5000 206.7000 35.8000 ;
	    RECT 202.1000 35.2000 202.5000 35.3000 ;
	    RECT 202.9000 34.9000 203.3000 35.0000 ;
	    RECT 201.4000 34.6000 203.3000 34.9000 ;
	    RECT 201.4000 34.5000 201.8000 34.6000 ;
	    RECT 191.0000 34.1000 191.4000 34.2000 ;
	    RECT 191.8000 34.1000 192.2000 34.2000 ;
	    RECT 191.0000 33.8000 192.6000 34.1000 ;
	    RECT 193.3000 33.8000 194.6000 34.2000 ;
	    RECT 195.4000 33.9000 200.9000 34.2000 ;
	    RECT 195.4000 33.8000 196.2000 33.9000 ;
	    RECT 192.2000 33.6000 192.6000 33.8000 ;
	    RECT 190.2000 31.1000 190.6000 33.1000 ;
	    RECT 191.0000 32.8000 191.4000 33.2000 ;
	    RECT 191.9000 33.1000 193.7000 33.3000 ;
	    RECT 194.2000 33.1000 194.5000 33.8000 ;
	    RECT 191.8000 33.0000 193.8000 33.1000 ;
	    RECT 190.9000 32.4000 191.3000 32.8000 ;
	    RECT 191.8000 31.1000 192.2000 33.0000 ;
	    RECT 193.4000 31.1000 193.8000 33.0000 ;
	    RECT 194.2000 31.1000 194.6000 33.1000 ;
	    RECT 195.0000 31.1000 195.4000 33.5000 ;
	    RECT 197.5000 32.8000 197.8000 33.9000 ;
	    RECT 200.3000 33.8000 200.9000 33.9000 ;
	    RECT 200.6000 33.2000 200.9000 33.8000 ;
	    RECT 203.8000 33.6000 204.2000 35.3000 ;
	    RECT 205.4000 34.8000 205.8000 35.2000 ;
	    RECT 204.6000 33.8000 205.0000 34.6000 ;
	    RECT 205.5000 34.4000 205.8000 34.8000 ;
	    RECT 205.5000 34.1000 206.0000 34.4000 ;
	    RECT 205.6000 34.0000 206.0000 34.1000 ;
	    RECT 206.4000 33.8000 206.7000 35.5000 ;
	    RECT 207.1000 35.2000 207.4000 35.9000 ;
	    RECT 209.4000 35.7000 209.8000 39.9000 ;
	    RECT 211.6000 38.2000 212.0000 39.9000 ;
	    RECT 211.0000 37.9000 212.0000 38.2000 ;
	    RECT 213.8000 37.9000 214.2000 39.9000 ;
	    RECT 215.9000 37.9000 216.5000 39.9000 ;
	    RECT 211.0000 37.5000 211.4000 37.9000 ;
	    RECT 213.8000 37.6000 214.1000 37.9000 ;
	    RECT 212.7000 37.3000 214.5000 37.6000 ;
	    RECT 215.8000 37.5000 216.2000 37.9000 ;
	    RECT 212.7000 37.2000 213.1000 37.3000 ;
	    RECT 214.1000 37.2000 214.5000 37.3000 ;
	    RECT 211.0000 36.5000 211.4000 36.6000 ;
	    RECT 213.3000 36.5000 213.7000 36.6000 ;
	    RECT 211.0000 36.2000 213.7000 36.5000 ;
	    RECT 214.0000 36.5000 215.1000 36.8000 ;
	    RECT 214.0000 35.9000 214.3000 36.5000 ;
	    RECT 214.7000 36.4000 215.1000 36.5000 ;
	    RECT 215.9000 36.6000 216.6000 37.0000 ;
	    RECT 215.9000 36.1000 216.2000 36.6000 ;
	    RECT 211.9000 35.7000 214.3000 35.9000 ;
	    RECT 209.4000 35.6000 214.3000 35.7000 ;
	    RECT 215.0000 35.8000 216.2000 36.1000 ;
	    RECT 209.4000 35.5000 212.3000 35.6000 ;
	    RECT 209.4000 35.4000 212.2000 35.5000 ;
	    RECT 207.0000 35.1000 207.4000 35.2000 ;
	    RECT 207.8000 35.1000 208.2000 35.2000 ;
	    RECT 212.6000 35.1000 213.0000 35.2000 ;
	    RECT 207.0000 34.8000 208.2000 35.1000 ;
	    RECT 210.5000 34.8000 213.0000 35.1000 ;
	    RECT 206.4000 33.7000 206.8000 33.8000 ;
	    RECT 202.3000 33.3000 204.2000 33.6000 ;
	    RECT 205.3000 33.5000 206.8000 33.7000 ;
	    RECT 202.3000 33.2000 202.7000 33.3000 ;
	    RECT 200.6000 32.8000 201.0000 33.2000 ;
	    RECT 196.6000 32.1000 197.0000 32.5000 ;
	    RECT 197.4000 32.4000 197.8000 32.8000 ;
	    RECT 198.3000 32.7000 198.7000 32.8000 ;
	    RECT 198.3000 32.4000 199.7000 32.7000 ;
	    RECT 199.4000 32.1000 199.7000 32.4000 ;
	    RECT 201.4000 32.1000 201.8000 32.5000 ;
	    RECT 196.6000 31.8000 197.6000 32.1000 ;
	    RECT 197.2000 31.1000 197.6000 31.8000 ;
	    RECT 199.4000 31.1000 199.8000 32.1000 ;
	    RECT 201.4000 31.8000 202.1000 32.1000 ;
	    RECT 201.5000 31.1000 202.1000 31.8000 ;
	    RECT 203.8000 31.1000 204.2000 33.3000 ;
	    RECT 204.7000 33.4000 206.8000 33.5000 ;
	    RECT 204.7000 33.2000 205.6000 33.4000 ;
	    RECT 204.7000 33.1000 205.0000 33.2000 ;
	    RECT 207.1000 33.1000 207.4000 34.8000 ;
	    RECT 210.5000 34.7000 210.9000 34.8000 ;
	    RECT 211.8000 34.7000 212.2000 34.8000 ;
	    RECT 211.3000 34.2000 211.7000 34.3000 ;
	    RECT 215.0000 34.2000 215.3000 35.8000 ;
	    RECT 218.2000 35.6000 218.6000 39.9000 ;
	    RECT 219.8000 37.9000 220.2000 39.9000 ;
	    RECT 216.5000 35.3000 218.6000 35.6000 ;
	    RECT 219.9000 35.8000 220.2000 37.9000 ;
	    RECT 221.4000 35.9000 221.8000 39.9000 ;
	    RECT 219.9000 35.5000 221.1000 35.8000 ;
	    RECT 216.5000 35.2000 216.9000 35.3000 ;
	    RECT 217.3000 34.9000 217.7000 35.0000 ;
	    RECT 215.8000 34.6000 217.7000 34.9000 ;
	    RECT 215.8000 34.5000 216.2000 34.6000 ;
	    RECT 209.8000 33.9000 215.3000 34.2000 ;
	    RECT 209.8000 33.8000 210.6000 33.9000 ;
	    RECT 204.6000 31.1000 205.0000 33.1000 ;
	    RECT 206.7000 32.6000 207.4000 33.1000 ;
	    RECT 206.7000 31.1000 207.1000 32.6000 ;
	    RECT 209.4000 31.1000 209.8000 33.5000 ;
	    RECT 211.9000 32.8000 212.2000 33.9000 ;
	    RECT 214.7000 33.8000 215.1000 33.9000 ;
	    RECT 218.2000 33.6000 218.6000 35.3000 ;
	    RECT 219.8000 34.8000 220.2000 35.2000 ;
	    RECT 219.0000 33.8000 219.4000 34.6000 ;
	    RECT 219.9000 34.4000 220.2000 34.8000 ;
	    RECT 219.9000 34.1000 220.4000 34.4000 ;
	    RECT 220.0000 34.0000 220.4000 34.1000 ;
	    RECT 220.8000 33.8000 221.1000 35.5000 ;
	    RECT 221.5000 35.2000 221.8000 35.9000 ;
	    RECT 222.2000 35.7000 222.6000 39.9000 ;
	    RECT 224.4000 38.2000 224.8000 39.9000 ;
	    RECT 223.8000 37.9000 224.8000 38.2000 ;
	    RECT 226.6000 37.9000 227.0000 39.9000 ;
	    RECT 228.7000 37.9000 229.3000 39.9000 ;
	    RECT 223.8000 37.5000 224.2000 37.9000 ;
	    RECT 226.6000 37.6000 226.9000 37.9000 ;
	    RECT 225.5000 37.3000 227.3000 37.6000 ;
	    RECT 228.6000 37.5000 229.0000 37.9000 ;
	    RECT 225.5000 37.2000 225.9000 37.3000 ;
	    RECT 226.9000 37.2000 227.3000 37.3000 ;
	    RECT 223.8000 36.5000 224.2000 36.6000 ;
	    RECT 226.1000 36.5000 226.5000 36.6000 ;
	    RECT 223.8000 36.2000 226.5000 36.5000 ;
	    RECT 226.8000 36.5000 227.9000 36.8000 ;
	    RECT 226.8000 35.9000 227.1000 36.5000 ;
	    RECT 227.5000 36.4000 227.9000 36.5000 ;
	    RECT 228.7000 36.6000 229.4000 37.0000 ;
	    RECT 228.7000 36.1000 229.0000 36.6000 ;
	    RECT 224.7000 35.7000 227.1000 35.9000 ;
	    RECT 222.2000 35.6000 227.1000 35.7000 ;
	    RECT 227.8000 35.8000 229.0000 36.1000 ;
	    RECT 222.2000 35.5000 225.1000 35.6000 ;
	    RECT 222.2000 35.4000 225.0000 35.5000 ;
	    RECT 221.4000 34.8000 221.8000 35.2000 ;
	    RECT 225.4000 35.1000 225.8000 35.2000 ;
	    RECT 220.8000 33.7000 221.2000 33.8000 ;
	    RECT 216.7000 33.3000 218.6000 33.6000 ;
	    RECT 219.7000 33.5000 221.2000 33.7000 ;
	    RECT 216.7000 33.2000 217.1000 33.3000 ;
	    RECT 211.0000 32.1000 211.4000 32.5000 ;
	    RECT 211.8000 32.4000 212.2000 32.8000 ;
	    RECT 212.7000 32.7000 213.1000 32.8000 ;
	    RECT 212.7000 32.4000 214.1000 32.7000 ;
	    RECT 213.8000 32.1000 214.1000 32.4000 ;
	    RECT 215.8000 32.1000 216.2000 32.5000 ;
	    RECT 211.0000 31.8000 212.0000 32.1000 ;
	    RECT 211.6000 31.1000 212.0000 31.8000 ;
	    RECT 213.8000 31.1000 214.2000 32.1000 ;
	    RECT 215.8000 31.8000 216.5000 32.1000 ;
	    RECT 215.9000 31.1000 216.5000 31.8000 ;
	    RECT 218.2000 31.1000 218.6000 33.3000 ;
	    RECT 219.1000 33.4000 221.2000 33.5000 ;
	    RECT 219.1000 33.2000 220.0000 33.4000 ;
	    RECT 219.1000 33.1000 219.4000 33.2000 ;
	    RECT 221.5000 33.1000 221.8000 34.8000 ;
	    RECT 223.3000 34.8000 225.8000 35.1000 ;
	    RECT 223.3000 34.7000 223.7000 34.8000 ;
	    RECT 224.6000 34.7000 225.0000 34.8000 ;
	    RECT 224.1000 34.2000 224.5000 34.3000 ;
	    RECT 227.8000 34.2000 228.1000 35.8000 ;
	    RECT 231.0000 35.6000 231.4000 39.9000 ;
	    RECT 232.2000 36.8000 232.6000 37.2000 ;
	    RECT 232.2000 36.2000 232.5000 36.8000 ;
	    RECT 232.9000 36.2000 233.3000 39.9000 ;
	    RECT 231.8000 35.9000 232.5000 36.2000 ;
	    RECT 232.8000 35.9000 233.3000 36.2000 ;
	    RECT 235.0000 36.2000 235.4000 39.9000 ;
	    RECT 236.6000 36.2000 237.0000 39.9000 ;
	    RECT 235.0000 35.9000 237.0000 36.2000 ;
	    RECT 237.4000 35.9000 237.8000 39.9000 ;
	    RECT 238.6000 36.8000 239.0000 37.2000 ;
	    RECT 238.6000 36.2000 238.9000 36.8000 ;
	    RECT 239.3000 36.2000 239.7000 39.9000 ;
	    RECT 242.7000 36.3000 243.1000 39.9000 ;
	    RECT 238.2000 35.9000 238.9000 36.2000 ;
	    RECT 239.2000 35.9000 239.7000 36.2000 ;
	    RECT 242.2000 35.9000 243.1000 36.3000 ;
	    RECT 243.8000 35.9000 244.2000 39.9000 ;
	    RECT 244.6000 36.2000 245.0000 39.9000 ;
	    RECT 246.2000 36.2000 246.6000 39.9000 ;
	    RECT 244.6000 35.9000 246.6000 36.2000 ;
	    RECT 231.8000 35.8000 232.2000 35.9000 ;
	    RECT 229.3000 35.3000 231.4000 35.6000 ;
	    RECT 229.3000 35.2000 229.7000 35.3000 ;
	    RECT 230.1000 34.9000 230.5000 35.0000 ;
	    RECT 228.6000 34.6000 230.5000 34.9000 ;
	    RECT 228.6000 34.5000 229.0000 34.6000 ;
	    RECT 222.6000 33.9000 228.1000 34.2000 ;
	    RECT 222.6000 33.8000 223.4000 33.9000 ;
	    RECT 219.0000 31.1000 219.4000 33.1000 ;
	    RECT 221.1000 32.6000 221.8000 33.1000 ;
	    RECT 221.1000 31.1000 221.5000 32.6000 ;
	    RECT 222.2000 31.1000 222.6000 33.5000 ;
	    RECT 224.7000 33.2000 225.0000 33.9000 ;
	    RECT 225.4000 33.8000 225.8000 33.9000 ;
	    RECT 227.5000 33.8000 227.9000 33.9000 ;
	    RECT 231.0000 33.6000 231.4000 35.3000 ;
	    RECT 232.8000 34.2000 233.1000 35.9000 ;
	    RECT 237.4000 35.2000 237.7000 35.9000 ;
	    RECT 238.2000 35.8000 238.6000 35.9000 ;
	    RECT 233.4000 34.4000 233.8000 35.2000 ;
	    RECT 236.6000 34.9000 237.8000 35.2000 ;
	    RECT 231.8000 33.8000 233.1000 34.2000 ;
	    RECT 234.2000 34.1000 234.6000 34.2000 ;
	    RECT 233.8000 33.8000 234.6000 34.1000 ;
	    RECT 235.8000 33.8000 236.2000 34.6000 ;
	    RECT 229.5000 33.3000 231.4000 33.6000 ;
	    RECT 229.5000 33.2000 229.9000 33.3000 ;
	    RECT 223.8000 32.1000 224.2000 32.5000 ;
	    RECT 224.6000 32.4000 225.0000 33.2000 ;
	    RECT 225.5000 32.7000 225.9000 32.8000 ;
	    RECT 225.5000 32.4000 226.9000 32.7000 ;
	    RECT 226.6000 32.1000 226.9000 32.4000 ;
	    RECT 228.6000 32.1000 229.0000 32.5000 ;
	    RECT 223.8000 31.8000 224.8000 32.1000 ;
	    RECT 224.4000 31.1000 224.8000 31.8000 ;
	    RECT 226.6000 31.1000 227.0000 32.1000 ;
	    RECT 228.6000 31.8000 229.3000 32.1000 ;
	    RECT 228.7000 31.1000 229.3000 31.8000 ;
	    RECT 231.0000 31.1000 231.4000 33.3000 ;
	    RECT 231.9000 33.1000 232.2000 33.8000 ;
	    RECT 233.8000 33.6000 234.2000 33.8000 ;
	    RECT 232.7000 33.1000 234.5000 33.3000 ;
	    RECT 236.6000 33.1000 236.9000 34.9000 ;
	    RECT 237.4000 34.8000 237.8000 34.9000 ;
	    RECT 239.2000 34.2000 239.5000 35.9000 ;
	    RECT 239.8000 34.4000 240.2000 35.2000 ;
	    RECT 242.3000 34.2000 242.6000 35.9000 ;
	    RECT 243.0000 34.8000 243.4000 35.6000 ;
	    RECT 243.9000 35.2000 244.2000 35.9000 ;
	    RECT 245.8000 35.2000 246.2000 35.4000 ;
	    RECT 243.8000 34.9000 245.0000 35.2000 ;
	    RECT 245.8000 34.9000 246.6000 35.2000 ;
	    RECT 247.8000 35.1000 248.2000 39.9000 ;
	    RECT 250.7000 36.3000 251.1000 39.9000 ;
	    RECT 250.2000 35.9000 251.1000 36.3000 ;
	    RECT 243.8000 34.8000 244.2000 34.9000 ;
	    RECT 238.2000 33.8000 239.5000 34.2000 ;
	    RECT 240.6000 34.1000 241.0000 34.2000 ;
	    RECT 240.2000 33.8000 241.0000 34.1000 ;
	    RECT 242.2000 33.8000 242.6000 34.2000 ;
	    RECT 237.4000 33.1000 237.8000 33.2000 ;
	    RECT 238.3000 33.1000 238.6000 33.8000 ;
	    RECT 240.2000 33.6000 240.6000 33.8000 ;
	    RECT 239.1000 33.1000 240.9000 33.3000 ;
	    RECT 242.3000 33.2000 242.6000 33.8000 ;
	    RECT 231.8000 31.1000 232.2000 33.1000 ;
	    RECT 232.6000 33.0000 234.6000 33.1000 ;
	    RECT 232.6000 31.1000 233.0000 33.0000 ;
	    RECT 234.2000 31.1000 234.6000 33.0000 ;
	    RECT 236.6000 31.1000 237.0000 33.1000 ;
	    RECT 237.4000 32.8000 238.6000 33.1000 ;
	    RECT 237.3000 32.4000 237.7000 32.8000 ;
	    RECT 238.2000 31.1000 238.6000 32.8000 ;
	    RECT 239.0000 33.0000 241.0000 33.1000 ;
	    RECT 239.0000 31.1000 239.4000 33.0000 ;
	    RECT 240.6000 31.1000 241.0000 33.0000 ;
	    RECT 242.2000 32.8000 242.6000 33.2000 ;
	    RECT 243.8000 32.8000 244.2000 33.2000 ;
	    RECT 244.7000 33.1000 245.0000 34.9000 ;
	    RECT 246.2000 34.8000 246.6000 34.9000 ;
	    RECT 247.0000 34.8000 248.2000 35.1000 ;
	    RECT 245.4000 33.8000 245.8000 34.6000 ;
	    RECT 247.0000 34.2000 247.3000 34.8000 ;
	    RECT 247.0000 33.8000 247.4000 34.2000 ;
	    RECT 242.3000 32.1000 242.6000 32.8000 ;
	    RECT 243.9000 32.4000 244.3000 32.8000 ;
	    RECT 242.2000 31.1000 242.6000 32.1000 ;
	    RECT 244.6000 31.1000 245.0000 33.1000 ;
	    RECT 247.8000 31.1000 248.2000 34.8000 ;
	    RECT 250.3000 34.2000 250.6000 35.9000 ;
	    RECT 250.2000 33.8000 250.6000 34.2000 ;
	    RECT 250.3000 33.1000 250.6000 33.8000 ;
	    RECT 252.6000 34.1000 253.0000 39.9000 ;
	    RECT 254.7000 36.2000 255.1000 39.9000 ;
	    RECT 255.4000 36.8000 255.8000 37.2000 ;
	    RECT 255.5000 36.2000 255.8000 36.8000 ;
	    RECT 254.7000 35.9000 255.2000 36.2000 ;
	    RECT 255.5000 35.9000 256.2000 36.2000 ;
	    RECT 254.2000 34.4000 254.6000 35.2000 ;
	    RECT 254.9000 34.2000 255.2000 35.9000 ;
	    RECT 255.8000 35.8000 256.2000 35.9000 ;
	    RECT 256.6000 35.9000 257.0000 39.9000 ;
	    RECT 258.2000 37.9000 258.6000 39.9000 ;
	    RECT 256.6000 35.2000 256.9000 35.9000 ;
	    RECT 258.2000 35.8000 258.5000 37.9000 ;
	    RECT 261.1000 36.2000 261.5000 39.9000 ;
	    RECT 261.8000 36.8000 262.2000 37.2000 ;
	    RECT 261.9000 36.2000 262.2000 36.8000 ;
	    RECT 261.1000 35.9000 261.6000 36.2000 ;
	    RECT 261.9000 35.9000 262.6000 36.2000 ;
	    RECT 257.3000 35.5000 258.5000 35.8000 ;
	    RECT 256.6000 34.8000 257.0000 35.2000 ;
	    RECT 253.4000 34.1000 253.8000 34.2000 ;
	    RECT 252.6000 33.8000 254.2000 34.1000 ;
	    RECT 254.9000 33.8000 256.2000 34.2000 ;
	    RECT 251.8000 33.1000 252.2000 33.2000 ;
	    RECT 250.2000 32.8000 252.2000 33.1000 ;
	    RECT 250.3000 32.1000 250.6000 32.8000 ;
	    RECT 251.8000 32.4000 252.2000 32.8000 ;
	    RECT 250.2000 31.1000 250.6000 32.1000 ;
	    RECT 252.6000 31.1000 253.0000 33.8000 ;
	    RECT 253.8000 33.6000 254.2000 33.8000 ;
	    RECT 253.5000 33.1000 255.3000 33.3000 ;
	    RECT 255.8000 33.1000 256.1000 33.8000 ;
	    RECT 256.6000 33.1000 256.9000 34.8000 ;
	    RECT 257.3000 33.8000 257.6000 35.5000 ;
	    RECT 261.3000 35.2000 261.6000 35.9000 ;
	    RECT 262.2000 35.8000 262.6000 35.9000 ;
	    RECT 258.2000 34.8000 258.6000 35.2000 ;
	    RECT 258.2000 34.4000 258.5000 34.8000 ;
	    RECT 258.0000 34.1000 258.5000 34.4000 ;
	    RECT 259.0000 34.1000 259.4000 34.6000 ;
	    RECT 260.6000 34.4000 261.0000 35.2000 ;
	    RECT 261.3000 34.8000 261.8000 35.2000 ;
	    RECT 261.3000 34.2000 261.6000 34.8000 ;
	    RECT 259.8000 34.1000 260.2000 34.2000 ;
	    RECT 258.0000 34.0000 258.4000 34.1000 ;
	    RECT 259.0000 33.8000 260.6000 34.1000 ;
	    RECT 261.3000 33.8000 262.6000 34.2000 ;
	    RECT 263.0000 34.1000 263.4000 39.9000 ;
	    RECT 264.6000 35.9000 265.0000 39.9000 ;
	    RECT 265.4000 36.2000 265.8000 39.9000 ;
	    RECT 267.0000 36.2000 267.4000 39.9000 ;
	    RECT 265.4000 35.9000 267.4000 36.2000 ;
	    RECT 264.7000 35.2000 265.0000 35.9000 ;
	    RECT 266.6000 35.2000 267.0000 35.4000 ;
	    RECT 264.6000 34.9000 265.8000 35.2000 ;
	    RECT 266.6000 35.1000 267.4000 35.2000 ;
	    RECT 268.6000 35.1000 269.0000 39.9000 ;
	    RECT 266.6000 34.9000 269.0000 35.1000 ;
	    RECT 264.6000 34.8000 265.0000 34.9000 ;
	    RECT 263.8000 34.1000 264.2000 34.2000 ;
	    RECT 263.0000 33.8000 264.2000 34.1000 ;
	    RECT 257.2000 33.7000 257.6000 33.8000 ;
	    RECT 257.2000 33.5000 258.7000 33.7000 ;
	    RECT 260.2000 33.6000 260.6000 33.8000 ;
	    RECT 257.2000 33.4000 259.3000 33.5000 ;
	    RECT 258.4000 33.2000 259.3000 33.4000 ;
	    RECT 259.0000 33.1000 259.3000 33.2000 ;
	    RECT 259.9000 33.1000 261.7000 33.3000 ;
	    RECT 262.2000 33.1000 262.5000 33.8000 ;
	    RECT 253.4000 33.0000 255.4000 33.1000 ;
	    RECT 253.4000 31.1000 253.8000 33.0000 ;
	    RECT 255.0000 31.1000 255.4000 33.0000 ;
	    RECT 255.8000 31.1000 256.2000 33.1000 ;
	    RECT 256.6000 32.6000 257.3000 33.1000 ;
	    RECT 256.9000 32.2000 257.3000 32.6000 ;
	    RECT 256.6000 31.8000 257.3000 32.2000 ;
	    RECT 256.9000 31.1000 257.3000 31.8000 ;
	    RECT 259.0000 31.1000 259.4000 33.1000 ;
	    RECT 259.8000 33.0000 261.8000 33.1000 ;
	    RECT 259.8000 31.1000 260.2000 33.0000 ;
	    RECT 261.4000 31.1000 261.8000 33.0000 ;
	    RECT 262.2000 31.1000 262.6000 33.1000 ;
	    RECT 263.0000 31.1000 263.4000 33.8000 ;
	    RECT 263.8000 32.4000 264.2000 33.2000 ;
	    RECT 264.6000 32.8000 265.0000 33.2000 ;
	    RECT 265.5000 33.1000 265.8000 34.9000 ;
	    RECT 267.0000 34.8000 269.0000 34.9000 ;
	    RECT 266.2000 33.8000 266.6000 34.6000 ;
	    RECT 264.7000 32.4000 265.1000 32.8000 ;
	    RECT 265.4000 31.1000 265.8000 33.1000 ;
	    RECT 267.8000 32.4000 268.2000 33.2000 ;
	    RECT 268.6000 31.1000 269.0000 34.8000 ;
	    RECT 1.4000 26.1000 1.8000 29.9000 ;
	    RECT 3.0000 28.9000 3.4000 29.9000 ;
	    RECT 3.0000 27.2000 3.3000 28.9000 ;
	    RECT 5.9000 28.2000 6.3000 29.9000 ;
	    RECT 5.4000 27.9000 6.3000 28.2000 ;
	    RECT 8.6000 27.9000 9.0000 29.9000 ;
	    RECT 11.0000 28.9000 11.4000 29.9000 ;
	    RECT 9.3000 28.2000 9.7000 28.6000 ;
	    RECT 9.4000 28.1000 9.8000 28.2000 ;
	    RECT 11.0000 28.1000 11.3000 28.9000 ;
	    RECT 3.0000 27.1000 3.4000 27.2000 ;
	    RECT 3.0000 26.8000 4.1000 27.1000 ;
	    RECT 2.2000 26.1000 2.6000 26.2000 ;
	    RECT 1.4000 25.8000 2.6000 26.1000 ;
	    RECT 1.4000 21.1000 1.8000 25.8000 ;
	    RECT 2.2000 25.4000 2.6000 25.8000 ;
	    RECT 3.0000 25.1000 3.3000 26.8000 ;
	    RECT 3.8000 26.2000 4.1000 26.8000 ;
	    RECT 3.8000 25.8000 4.2000 26.2000 ;
	    RECT 5.4000 26.1000 5.8000 27.9000 ;
	    RECT 7.8000 26.4000 8.2000 27.2000 ;
	    RECT 7.0000 26.1000 7.4000 26.2000 ;
	    RECT 8.6000 26.1000 8.9000 27.9000 ;
	    RECT 9.4000 27.8000 11.3000 28.1000 ;
	    RECT 11.0000 27.2000 11.3000 27.8000 ;
	    RECT 11.0000 26.8000 11.4000 27.2000 ;
	    RECT 11.8000 26.8000 12.2000 27.2000 ;
	    RECT 9.4000 26.1000 9.8000 26.2000 ;
	    RECT 5.4000 25.8000 7.8000 26.1000 ;
	    RECT 8.6000 25.8000 9.8000 26.1000 ;
	    RECT 2.5000 24.7000 3.4000 25.1000 ;
	    RECT 2.5000 21.1000 2.9000 24.7000 ;
	    RECT 5.4000 21.1000 5.8000 25.8000 ;
	    RECT 7.4000 25.6000 7.8000 25.8000 ;
	    RECT 6.2000 24.4000 6.6000 25.2000 ;
	    RECT 9.4000 25.1000 9.7000 25.8000 ;
	    RECT 10.2000 25.4000 10.6000 26.2000 ;
	    RECT 11.0000 25.1000 11.3000 26.8000 ;
	    RECT 11.8000 26.1000 12.1000 26.8000 ;
	    RECT 12.6000 26.1000 13.0000 29.9000 ;
	    RECT 15.5000 28.2000 15.9000 29.9000 ;
	    RECT 16.7000 28.2000 17.1000 28.6000 ;
	    RECT 11.8000 25.8000 13.0000 26.1000 ;
	    RECT 7.0000 24.8000 9.0000 25.1000 ;
	    RECT 7.0000 21.1000 7.4000 24.8000 ;
	    RECT 8.6000 21.1000 9.0000 24.8000 ;
	    RECT 9.4000 21.1000 9.8000 25.1000 ;
	    RECT 10.5000 24.7000 11.4000 25.1000 ;
	    RECT 10.5000 21.1000 10.9000 24.7000 ;
	    RECT 12.6000 21.1000 13.0000 25.8000 ;
	    RECT 15.0000 27.9000 15.9000 28.2000 ;
	    RECT 15.0000 21.1000 15.4000 27.9000 ;
	    RECT 16.6000 27.8000 17.0000 28.2000 ;
	    RECT 17.4000 27.9000 17.8000 29.9000 ;
	    RECT 17.5000 26.2000 17.8000 27.9000 ;
	    RECT 18.2000 26.4000 18.6000 27.2000 ;
	    RECT 16.6000 26.1000 17.0000 26.2000 ;
	    RECT 17.4000 26.1000 17.8000 26.2000 ;
	    RECT 19.0000 26.1000 19.4000 26.2000 ;
	    RECT 19.8000 26.1000 20.2000 29.9000 ;
	    RECT 20.6000 27.8000 21.0000 28.6000 ;
	    RECT 21.7000 28.2000 22.1000 29.9000 ;
	    RECT 21.7000 27.9000 22.6000 28.2000 ;
	    RECT 23.8000 27.9000 24.2000 29.9000 ;
	    RECT 24.6000 28.0000 25.0000 29.9000 ;
	    RECT 26.2000 28.0000 26.6000 29.9000 ;
	    RECT 24.6000 27.9000 26.6000 28.0000 ;
	    RECT 27.8000 28.9000 28.2000 29.9000 ;
	    RECT 16.6000 25.8000 17.8000 26.1000 ;
	    RECT 18.6000 25.8000 20.2000 26.1000 ;
	    RECT 16.7000 25.1000 17.0000 25.8000 ;
	    RECT 18.6000 25.6000 19.0000 25.8000 ;
	    RECT 16.6000 21.1000 17.0000 25.1000 ;
	    RECT 17.4000 24.8000 19.4000 25.1000 ;
	    RECT 17.4000 21.1000 17.8000 24.8000 ;
	    RECT 19.0000 21.1000 19.4000 24.8000 ;
	    RECT 19.8000 21.1000 20.2000 25.8000 ;
	    RECT 20.6000 25.1000 21.0000 25.2000 ;
	    RECT 21.4000 25.1000 21.8000 25.2000 ;
	    RECT 20.6000 24.8000 21.8000 25.1000 ;
	    RECT 21.4000 24.4000 21.8000 24.8000 ;
	    RECT 22.2000 21.1000 22.6000 27.9000 ;
	    RECT 23.0000 27.1000 23.4000 27.6000 ;
	    RECT 23.9000 27.2000 24.2000 27.9000 ;
	    RECT 24.7000 27.7000 26.5000 27.9000 ;
	    RECT 25.8000 27.2000 26.2000 27.4000 ;
	    RECT 27.8000 27.2000 28.1000 28.9000 ;
	    RECT 30.7000 28.2000 31.1000 29.9000 ;
	    RECT 30.2000 27.9000 31.1000 28.2000 ;
	    RECT 23.8000 27.1000 25.1000 27.2000 ;
	    RECT 23.0000 26.8000 25.1000 27.1000 ;
	    RECT 25.8000 27.1000 26.6000 27.2000 ;
	    RECT 27.8000 27.1000 28.2000 27.2000 ;
	    RECT 25.8000 26.9000 28.2000 27.1000 ;
	    RECT 26.2000 26.8000 28.2000 26.9000 ;
	    RECT 23.8000 25.1000 24.2000 25.2000 ;
	    RECT 24.8000 25.1000 25.1000 26.8000 ;
	    RECT 25.4000 25.8000 25.8000 26.6000 ;
	    RECT 27.0000 25.4000 27.4000 26.2000 ;
	    RECT 27.8000 25.1000 28.1000 26.8000 ;
	    RECT 29.4000 25.8000 29.8000 26.2000 ;
	    RECT 29.4000 25.1000 29.7000 25.8000 ;
	    RECT 30.2000 25.1000 30.6000 27.9000 ;
	    RECT 31.0000 26.8000 31.4000 27.2000 ;
	    RECT 31.0000 26.1000 31.3000 26.8000 ;
	    RECT 31.8000 26.1000 32.2000 29.9000 ;
	    RECT 33.4000 27.5000 33.8000 29.9000 ;
	    RECT 35.6000 29.2000 36.0000 29.9000 ;
	    RECT 35.0000 28.9000 36.0000 29.2000 ;
	    RECT 37.8000 28.9000 38.2000 29.9000 ;
	    RECT 39.9000 29.2000 40.5000 29.9000 ;
	    RECT 39.8000 28.9000 40.5000 29.2000 ;
	    RECT 35.0000 28.5000 35.4000 28.9000 ;
	    RECT 37.8000 28.6000 38.1000 28.9000 ;
	    RECT 35.8000 28.2000 36.2000 28.6000 ;
	    RECT 36.7000 28.3000 38.1000 28.6000 ;
	    RECT 39.8000 28.5000 40.2000 28.9000 ;
	    RECT 36.7000 28.2000 37.1000 28.3000 ;
	    RECT 33.8000 27.1000 34.6000 27.2000 ;
	    RECT 35.9000 27.1000 36.2000 28.2000 ;
	    RECT 40.7000 27.7000 41.1000 27.8000 ;
	    RECT 42.2000 27.7000 42.6000 29.9000 ;
	    RECT 40.7000 27.4000 42.6000 27.7000 ;
	    RECT 43.0000 27.5000 43.4000 29.9000 ;
	    RECT 45.2000 29.2000 45.6000 29.9000 ;
	    RECT 44.6000 28.9000 45.6000 29.2000 ;
	    RECT 47.4000 28.9000 47.8000 29.9000 ;
	    RECT 49.5000 29.2000 50.1000 29.9000 ;
	    RECT 49.4000 28.9000 50.1000 29.2000 ;
	    RECT 44.6000 28.5000 45.0000 28.9000 ;
	    RECT 47.4000 28.6000 47.7000 28.9000 ;
	    RECT 45.4000 28.2000 45.8000 28.6000 ;
	    RECT 46.3000 28.3000 47.7000 28.6000 ;
	    RECT 49.4000 28.5000 49.8000 28.9000 ;
	    RECT 46.3000 28.2000 46.7000 28.3000 ;
	    RECT 38.7000 27.1000 39.1000 27.2000 ;
	    RECT 33.8000 26.8000 39.3000 27.1000 ;
	    RECT 35.3000 26.7000 35.7000 26.8000 ;
	    RECT 31.0000 25.8000 32.2000 26.1000 ;
	    RECT 34.5000 26.2000 34.9000 26.3000 ;
	    RECT 39.0000 26.2000 39.3000 26.8000 ;
	    RECT 39.8000 26.4000 40.2000 26.5000 ;
	    RECT 34.5000 25.9000 37.0000 26.2000 ;
	    RECT 36.6000 25.8000 37.0000 25.9000 ;
	    RECT 39.0000 25.8000 39.4000 26.2000 ;
	    RECT 39.8000 26.1000 41.7000 26.4000 ;
	    RECT 41.3000 26.0000 41.7000 26.1000 ;
	    RECT 23.8000 24.8000 24.5000 25.1000 ;
	    RECT 24.8000 24.8000 25.3000 25.1000 ;
	    RECT 24.2000 24.2000 24.5000 24.8000 ;
	    RECT 24.2000 23.8000 24.6000 24.2000 ;
	    RECT 24.9000 21.1000 25.3000 24.8000 ;
	    RECT 27.3000 24.7000 28.2000 25.1000 ;
	    RECT 29.4000 24.8000 30.6000 25.1000 ;
	    RECT 27.3000 21.1000 27.7000 24.7000 ;
	    RECT 30.2000 21.1000 30.6000 24.8000 ;
	    RECT 31.0000 25.1000 31.4000 25.2000 ;
	    RECT 31.8000 25.1000 32.2000 25.8000 ;
	    RECT 31.0000 24.8000 32.2000 25.1000 ;
	    RECT 31.0000 24.4000 31.4000 24.8000 ;
	    RECT 31.8000 21.1000 32.2000 24.8000 ;
	    RECT 33.4000 25.5000 36.2000 25.6000 ;
	    RECT 33.4000 25.4000 36.3000 25.5000 ;
	    RECT 33.4000 25.3000 38.3000 25.4000 ;
	    RECT 33.4000 21.1000 33.8000 25.3000 ;
	    RECT 35.9000 25.1000 38.3000 25.3000 ;
	    RECT 35.0000 24.5000 37.7000 24.8000 ;
	    RECT 35.0000 24.4000 35.4000 24.5000 ;
	    RECT 37.3000 24.4000 37.7000 24.5000 ;
	    RECT 38.0000 24.5000 38.3000 25.1000 ;
	    RECT 39.0000 25.2000 39.3000 25.8000 ;
	    RECT 40.5000 25.7000 40.9000 25.8000 ;
	    RECT 42.2000 25.7000 42.6000 27.4000 ;
	    RECT 43.4000 27.1000 44.2000 27.2000 ;
	    RECT 45.5000 27.1000 45.8000 28.2000 ;
	    RECT 50.3000 27.7000 50.7000 27.8000 ;
	    RECT 51.8000 27.7000 52.2000 29.9000 ;
	    RECT 50.3000 27.4000 52.2000 27.7000 ;
	    RECT 48.3000 27.1000 48.7000 27.2000 ;
	    RECT 43.4000 26.8000 48.9000 27.1000 ;
	    RECT 44.9000 26.7000 45.3000 26.8000 ;
	    RECT 44.1000 26.2000 44.5000 26.3000 ;
	    RECT 45.4000 26.2000 45.8000 26.3000 ;
	    RECT 48.6000 26.2000 48.9000 26.8000 ;
	    RECT 49.4000 26.4000 49.8000 26.5000 ;
	    RECT 44.1000 25.9000 46.6000 26.2000 ;
	    RECT 46.2000 25.8000 46.6000 25.9000 ;
	    RECT 48.6000 25.8000 49.0000 26.2000 ;
	    RECT 49.4000 26.1000 51.3000 26.4000 ;
	    RECT 50.9000 26.0000 51.3000 26.1000 ;
	    RECT 40.5000 25.4000 42.6000 25.7000 ;
	    RECT 39.0000 24.9000 40.2000 25.2000 ;
	    RECT 38.7000 24.5000 39.1000 24.6000 ;
	    RECT 38.0000 24.2000 39.1000 24.5000 ;
	    RECT 39.9000 24.4000 40.2000 24.9000 ;
	    RECT 39.9000 24.0000 40.6000 24.4000 ;
	    RECT 36.7000 23.7000 37.1000 23.8000 ;
	    RECT 38.1000 23.7000 38.5000 23.8000 ;
	    RECT 35.0000 23.1000 35.4000 23.5000 ;
	    RECT 36.7000 23.4000 38.5000 23.7000 ;
	    RECT 37.8000 23.1000 38.1000 23.4000 ;
	    RECT 39.8000 23.1000 40.2000 23.5000 ;
	    RECT 35.0000 22.8000 36.0000 23.1000 ;
	    RECT 35.6000 21.1000 36.0000 22.8000 ;
	    RECT 37.8000 21.1000 38.2000 23.1000 ;
	    RECT 39.9000 21.1000 40.5000 23.1000 ;
	    RECT 42.2000 21.1000 42.6000 25.4000 ;
	    RECT 43.0000 25.5000 45.8000 25.6000 ;
	    RECT 43.0000 25.4000 45.9000 25.5000 ;
	    RECT 43.0000 25.3000 47.9000 25.4000 ;
	    RECT 43.0000 21.1000 43.4000 25.3000 ;
	    RECT 45.5000 25.1000 47.9000 25.3000 ;
	    RECT 44.6000 24.5000 47.3000 24.8000 ;
	    RECT 44.6000 24.4000 45.0000 24.5000 ;
	    RECT 46.9000 24.4000 47.3000 24.5000 ;
	    RECT 47.6000 24.5000 47.9000 25.1000 ;
	    RECT 48.6000 25.2000 48.9000 25.8000 ;
	    RECT 50.1000 25.7000 50.5000 25.8000 ;
	    RECT 51.8000 25.7000 52.2000 27.4000 ;
	    RECT 53.4000 28.9000 53.8000 29.9000 ;
	    RECT 53.4000 27.2000 53.7000 28.9000 ;
	    RECT 54.2000 28.1000 54.6000 28.6000 ;
	    RECT 55.0000 28.1000 55.4000 29.9000 ;
	    RECT 54.2000 27.8000 55.4000 28.1000 ;
	    RECT 55.8000 27.8000 56.2000 28.6000 ;
	    RECT 53.4000 26.8000 53.8000 27.2000 ;
	    RECT 54.2000 26.8000 54.6000 27.2000 ;
	    RECT 50.1000 25.4000 52.2000 25.7000 ;
	    RECT 52.6000 25.4000 53.0000 26.2000 ;
	    RECT 53.4000 26.1000 53.7000 26.8000 ;
	    RECT 54.2000 26.1000 54.5000 26.8000 ;
	    RECT 53.4000 25.8000 54.5000 26.1000 ;
	    RECT 48.6000 24.9000 49.8000 25.2000 ;
	    RECT 48.3000 24.5000 48.7000 24.6000 ;
	    RECT 47.6000 24.2000 48.7000 24.5000 ;
	    RECT 49.5000 24.4000 49.8000 24.9000 ;
	    RECT 49.5000 24.0000 50.2000 24.4000 ;
	    RECT 46.3000 23.7000 46.7000 23.8000 ;
	    RECT 47.7000 23.7000 48.1000 23.8000 ;
	    RECT 44.6000 23.1000 45.0000 23.5000 ;
	    RECT 46.3000 23.4000 48.1000 23.7000 ;
	    RECT 47.4000 23.1000 47.7000 23.4000 ;
	    RECT 49.4000 23.1000 49.8000 23.5000 ;
	    RECT 44.6000 22.8000 45.6000 23.1000 ;
	    RECT 45.2000 21.1000 45.6000 22.8000 ;
	    RECT 47.4000 21.1000 47.8000 23.1000 ;
	    RECT 49.5000 21.1000 50.1000 23.1000 ;
	    RECT 51.8000 21.1000 52.2000 25.4000 ;
	    RECT 53.4000 25.1000 53.7000 25.8000 ;
	    RECT 52.9000 24.7000 53.8000 25.1000 ;
	    RECT 52.9000 21.1000 53.3000 24.7000 ;
	    RECT 55.0000 21.1000 55.4000 27.8000 ;
	    RECT 58.2000 27.5000 58.6000 29.9000 ;
	    RECT 60.4000 29.2000 60.8000 29.9000 ;
	    RECT 59.8000 28.9000 60.8000 29.2000 ;
	    RECT 62.6000 28.9000 63.0000 29.9000 ;
	    RECT 64.7000 29.2000 65.3000 29.9000 ;
	    RECT 64.6000 28.9000 65.3000 29.2000 ;
	    RECT 59.8000 28.5000 60.2000 28.9000 ;
	    RECT 62.6000 28.6000 62.9000 28.9000 ;
	    RECT 60.6000 28.2000 61.0000 28.6000 ;
	    RECT 61.5000 28.3000 62.9000 28.6000 ;
	    RECT 64.6000 28.5000 65.0000 28.9000 ;
	    RECT 61.5000 28.2000 61.9000 28.3000 ;
	    RECT 58.6000 27.1000 59.4000 27.2000 ;
	    RECT 60.7000 27.1000 61.0000 28.2000 ;
	    RECT 65.5000 27.7000 65.9000 27.8000 ;
	    RECT 67.0000 27.7000 67.4000 29.9000 ;
	    RECT 67.8000 28.0000 68.2000 29.9000 ;
	    RECT 69.4000 28.0000 69.8000 29.9000 ;
	    RECT 67.8000 27.9000 69.8000 28.0000 ;
	    RECT 70.2000 27.9000 70.6000 29.9000 ;
	    RECT 71.8000 28.9000 72.2000 29.9000 ;
	    RECT 67.9000 27.7000 69.7000 27.9000 ;
	    RECT 65.5000 27.4000 67.4000 27.7000 ;
	    RECT 63.5000 27.1000 63.9000 27.2000 ;
	    RECT 58.6000 26.8000 64.1000 27.1000 ;
	    RECT 60.1000 26.7000 60.5000 26.8000 ;
	    RECT 59.3000 26.2000 59.7000 26.3000 ;
	    RECT 60.6000 26.2000 61.0000 26.3000 ;
	    RECT 63.8000 26.2000 64.1000 26.8000 ;
	    RECT 64.6000 26.4000 65.0000 26.5000 ;
	    RECT 59.3000 25.9000 61.8000 26.2000 ;
	    RECT 61.4000 25.8000 61.8000 25.9000 ;
	    RECT 63.8000 25.8000 64.2000 26.2000 ;
	    RECT 64.6000 26.1000 66.5000 26.4000 ;
	    RECT 66.1000 26.0000 66.5000 26.1000 ;
	    RECT 58.2000 25.5000 61.0000 25.6000 ;
	    RECT 58.2000 25.4000 61.1000 25.5000 ;
	    RECT 58.2000 25.3000 63.1000 25.4000 ;
	    RECT 58.2000 21.1000 58.6000 25.3000 ;
	    RECT 60.7000 25.1000 63.1000 25.3000 ;
	    RECT 59.8000 24.5000 62.5000 24.8000 ;
	    RECT 59.8000 24.4000 60.2000 24.5000 ;
	    RECT 62.1000 24.4000 62.5000 24.5000 ;
	    RECT 62.8000 24.5000 63.1000 25.1000 ;
	    RECT 63.8000 25.2000 64.1000 25.8000 ;
	    RECT 65.3000 25.7000 65.7000 25.8000 ;
	    RECT 67.0000 25.7000 67.4000 27.4000 ;
	    RECT 68.2000 27.2000 68.6000 27.4000 ;
	    RECT 70.2000 27.2000 70.5000 27.9000 ;
	    RECT 71.8000 27.2000 72.1000 28.9000 ;
	    RECT 72.6000 27.8000 73.0000 28.6000 ;
	    RECT 73.4000 27.5000 73.8000 29.9000 ;
	    RECT 75.6000 29.2000 76.0000 29.9000 ;
	    RECT 75.0000 28.9000 76.0000 29.2000 ;
	    RECT 77.8000 28.9000 78.2000 29.9000 ;
	    RECT 79.9000 29.2000 80.5000 29.9000 ;
	    RECT 79.8000 28.9000 80.5000 29.2000 ;
	    RECT 75.0000 28.5000 75.4000 28.9000 ;
	    RECT 77.8000 28.6000 78.1000 28.9000 ;
	    RECT 75.8000 28.2000 76.2000 28.6000 ;
	    RECT 76.7000 28.3000 78.1000 28.6000 ;
	    RECT 79.8000 28.5000 80.2000 28.9000 ;
	    RECT 76.7000 28.2000 77.1000 28.3000 ;
	    RECT 67.8000 26.9000 68.6000 27.2000 ;
	    RECT 67.8000 26.8000 68.2000 26.9000 ;
	    RECT 69.3000 26.8000 70.6000 27.2000 ;
	    RECT 71.8000 26.8000 72.2000 27.2000 ;
	    RECT 73.8000 27.1000 74.6000 27.2000 ;
	    RECT 75.9000 27.1000 76.2000 28.2000 ;
	    RECT 80.7000 27.7000 81.1000 27.8000 ;
	    RECT 82.2000 27.7000 82.6000 29.9000 ;
	    RECT 80.7000 27.4000 82.6000 27.7000 ;
	    RECT 78.7000 27.1000 79.1000 27.2000 ;
	    RECT 73.8000 26.8000 79.3000 27.1000 ;
	    RECT 68.6000 25.8000 69.0000 26.6000 ;
	    RECT 69.3000 26.1000 69.6000 26.8000 ;
	    RECT 71.0000 26.1000 71.4000 26.2000 ;
	    RECT 69.3000 25.8000 71.4000 26.1000 ;
	    RECT 65.3000 25.4000 67.4000 25.7000 ;
	    RECT 63.8000 24.9000 65.0000 25.2000 ;
	    RECT 63.5000 24.5000 63.9000 24.6000 ;
	    RECT 62.8000 24.2000 63.9000 24.5000 ;
	    RECT 64.7000 24.4000 65.0000 24.9000 ;
	    RECT 64.7000 24.0000 65.4000 24.4000 ;
	    RECT 61.5000 23.7000 61.9000 23.8000 ;
	    RECT 62.9000 23.7000 63.3000 23.8000 ;
	    RECT 59.8000 23.1000 60.2000 23.5000 ;
	    RECT 61.5000 23.4000 63.3000 23.7000 ;
	    RECT 62.6000 23.1000 62.9000 23.4000 ;
	    RECT 64.6000 23.1000 65.0000 23.5000 ;
	    RECT 59.8000 22.8000 60.8000 23.1000 ;
	    RECT 60.4000 21.1000 60.8000 22.8000 ;
	    RECT 62.6000 21.1000 63.0000 23.1000 ;
	    RECT 64.7000 21.1000 65.3000 23.1000 ;
	    RECT 67.0000 21.1000 67.4000 25.4000 ;
	    RECT 69.3000 25.1000 69.6000 25.8000 ;
	    RECT 71.0000 25.4000 71.4000 25.8000 ;
	    RECT 71.8000 25.2000 72.1000 26.8000 ;
	    RECT 75.3000 26.7000 75.7000 26.8000 ;
	    RECT 74.5000 26.2000 74.9000 26.3000 ;
	    RECT 75.8000 26.2000 76.2000 26.3000 ;
	    RECT 74.5000 25.9000 77.0000 26.2000 ;
	    RECT 76.6000 25.8000 77.0000 25.9000 ;
	    RECT 78.2000 26.1000 78.6000 26.2000 ;
	    RECT 79.0000 26.1000 79.3000 26.8000 ;
	    RECT 79.8000 26.4000 80.2000 26.5000 ;
	    RECT 79.8000 26.1000 81.7000 26.4000 ;
	    RECT 78.2000 25.8000 79.3000 26.1000 ;
	    RECT 81.3000 26.0000 81.7000 26.1000 ;
	    RECT 73.4000 25.5000 76.2000 25.6000 ;
	    RECT 73.4000 25.4000 76.3000 25.5000 ;
	    RECT 73.4000 25.3000 78.3000 25.4000 ;
	    RECT 70.2000 25.1000 70.6000 25.2000 ;
	    RECT 71.8000 25.1000 72.2000 25.2000 ;
	    RECT 69.1000 24.8000 69.6000 25.1000 ;
	    RECT 69.9000 24.8000 70.6000 25.1000 ;
	    RECT 69.1000 21.1000 69.5000 24.8000 ;
	    RECT 69.9000 24.2000 70.2000 24.8000 ;
	    RECT 69.8000 23.8000 70.2000 24.2000 ;
	    RECT 71.3000 24.7000 72.2000 25.1000 ;
	    RECT 71.3000 21.1000 71.7000 24.7000 ;
	    RECT 73.4000 21.1000 73.8000 25.3000 ;
	    RECT 75.9000 25.1000 78.3000 25.3000 ;
	    RECT 75.0000 24.5000 77.7000 24.8000 ;
	    RECT 75.0000 24.4000 75.4000 24.5000 ;
	    RECT 77.3000 24.4000 77.7000 24.5000 ;
	    RECT 78.0000 24.5000 78.3000 25.1000 ;
	    RECT 79.0000 25.2000 79.3000 25.8000 ;
	    RECT 80.5000 25.7000 80.9000 25.8000 ;
	    RECT 82.2000 25.7000 82.6000 27.4000 ;
	    RECT 80.5000 25.4000 82.6000 25.7000 ;
	    RECT 79.0000 24.9000 80.2000 25.2000 ;
	    RECT 78.7000 24.5000 79.1000 24.6000 ;
	    RECT 78.0000 24.2000 79.1000 24.5000 ;
	    RECT 79.9000 24.4000 80.2000 24.9000 ;
	    RECT 79.9000 24.0000 80.6000 24.4000 ;
	    RECT 76.7000 23.7000 77.1000 23.8000 ;
	    RECT 78.1000 23.7000 78.5000 23.8000 ;
	    RECT 75.0000 23.1000 75.4000 23.5000 ;
	    RECT 76.7000 23.4000 78.5000 23.7000 ;
	    RECT 77.8000 23.1000 78.1000 23.4000 ;
	    RECT 79.8000 23.1000 80.2000 23.5000 ;
	    RECT 75.0000 22.8000 76.0000 23.1000 ;
	    RECT 75.6000 21.1000 76.0000 22.8000 ;
	    RECT 77.8000 21.1000 78.2000 23.1000 ;
	    RECT 79.9000 21.1000 80.5000 23.1000 ;
	    RECT 82.2000 21.1000 82.6000 25.4000 ;
	    RECT 83.0000 27.7000 83.4000 29.9000 ;
	    RECT 85.1000 29.2000 85.7000 29.9000 ;
	    RECT 85.1000 28.9000 85.8000 29.2000 ;
	    RECT 87.4000 28.9000 87.8000 29.9000 ;
	    RECT 89.6000 29.2000 90.0000 29.9000 ;
	    RECT 89.6000 28.9000 90.6000 29.2000 ;
	    RECT 85.4000 28.5000 85.8000 28.9000 ;
	    RECT 87.5000 28.6000 87.8000 28.9000 ;
	    RECT 87.5000 28.3000 88.9000 28.6000 ;
	    RECT 88.5000 28.2000 88.9000 28.3000 ;
	    RECT 89.4000 28.2000 89.8000 28.6000 ;
	    RECT 90.2000 28.5000 90.6000 28.9000 ;
	    RECT 84.5000 27.7000 84.9000 27.8000 ;
	    RECT 83.0000 27.4000 84.9000 27.7000 ;
	    RECT 83.0000 25.7000 83.4000 27.4000 ;
	    RECT 86.5000 27.1000 86.9000 27.2000 ;
	    RECT 89.4000 27.1000 89.7000 28.2000 ;
	    RECT 91.8000 27.5000 92.2000 29.9000 ;
	    RECT 93.4000 28.9000 93.8000 29.9000 ;
	    RECT 92.6000 27.8000 93.0000 28.6000 ;
	    RECT 93.5000 27.2000 93.8000 28.9000 ;
	    RECT 95.3000 28.2000 95.7000 29.9000 ;
	    RECT 95.3000 27.9000 96.2000 28.2000 ;
	    RECT 91.0000 27.1000 91.8000 27.2000 ;
	    RECT 86.3000 26.8000 91.8000 27.1000 ;
	    RECT 93.4000 26.8000 93.8000 27.2000 ;
	    RECT 85.4000 26.4000 85.8000 26.5000 ;
	    RECT 83.9000 26.1000 85.8000 26.4000 ;
	    RECT 86.3000 26.2000 86.6000 26.8000 ;
	    RECT 89.9000 26.7000 90.3000 26.8000 ;
	    RECT 89.4000 26.2000 89.8000 26.3000 ;
	    RECT 90.7000 26.2000 91.1000 26.3000 ;
	    RECT 83.9000 26.0000 84.3000 26.1000 ;
	    RECT 86.2000 25.8000 86.6000 26.2000 ;
	    RECT 88.6000 25.9000 91.1000 26.2000 ;
	    RECT 88.6000 25.8000 89.0000 25.9000 ;
	    RECT 84.7000 25.7000 85.1000 25.8000 ;
	    RECT 83.0000 25.4000 85.1000 25.7000 ;
	    RECT 83.0000 21.1000 83.4000 25.4000 ;
	    RECT 86.3000 25.2000 86.6000 25.8000 ;
	    RECT 89.4000 25.5000 92.2000 25.6000 ;
	    RECT 89.3000 25.4000 92.2000 25.5000 ;
	    RECT 85.4000 24.9000 86.6000 25.2000 ;
	    RECT 87.3000 25.3000 92.2000 25.4000 ;
	    RECT 87.3000 25.1000 89.7000 25.3000 ;
	    RECT 85.4000 24.4000 85.7000 24.9000 ;
	    RECT 85.0000 24.0000 85.7000 24.4000 ;
	    RECT 86.5000 24.5000 86.9000 24.6000 ;
	    RECT 87.3000 24.5000 87.6000 25.1000 ;
	    RECT 86.5000 24.2000 87.6000 24.5000 ;
	    RECT 87.9000 24.5000 90.6000 24.8000 ;
	    RECT 87.9000 24.4000 88.3000 24.5000 ;
	    RECT 90.2000 24.4000 90.6000 24.5000 ;
	    RECT 87.1000 23.7000 87.5000 23.8000 ;
	    RECT 88.5000 23.7000 88.9000 23.8000 ;
	    RECT 85.4000 23.1000 85.8000 23.5000 ;
	    RECT 87.1000 23.4000 88.9000 23.7000 ;
	    RECT 87.5000 23.1000 87.8000 23.4000 ;
	    RECT 90.2000 23.1000 90.6000 23.5000 ;
	    RECT 85.1000 21.1000 85.7000 23.1000 ;
	    RECT 87.4000 21.1000 87.8000 23.1000 ;
	    RECT 89.6000 22.8000 90.6000 23.1000 ;
	    RECT 89.6000 21.1000 90.0000 22.8000 ;
	    RECT 91.8000 21.1000 92.2000 25.3000 ;
	    RECT 93.5000 25.2000 93.8000 26.8000 ;
	    RECT 94.2000 26.1000 94.6000 26.2000 ;
	    RECT 95.8000 26.1000 96.2000 27.9000 ;
	    RECT 99.0000 27.9000 99.4000 29.9000 ;
	    RECT 101.9000 29.2000 102.3000 29.9000 ;
	    RECT 101.9000 28.8000 102.6000 29.2000 ;
	    RECT 99.7000 28.2000 100.1000 28.6000 ;
	    RECT 101.9000 28.2000 102.3000 28.8000 ;
	    RECT 96.6000 26.8000 97.0000 27.6000 ;
	    RECT 98.2000 26.4000 98.6000 27.2000 ;
	    RECT 94.2000 25.8000 96.2000 26.1000 ;
	    RECT 97.4000 26.1000 97.8000 26.2000 ;
	    RECT 99.0000 26.1000 99.3000 27.9000 ;
	    RECT 99.8000 27.8000 100.2000 28.2000 ;
	    RECT 101.4000 27.9000 102.3000 28.2000 ;
	    RECT 100.6000 26.8000 101.0000 27.6000 ;
	    RECT 99.8000 26.1000 100.2000 26.2000 ;
	    RECT 97.4000 25.8000 98.2000 26.1000 ;
	    RECT 99.0000 25.8000 100.2000 26.1000 ;
	    RECT 94.2000 25.4000 94.6000 25.8000 ;
	    RECT 93.4000 25.1000 93.8000 25.2000 ;
	    RECT 93.4000 24.7000 94.3000 25.1000 ;
	    RECT 93.9000 21.1000 94.3000 24.7000 ;
	    RECT 95.0000 24.4000 95.4000 25.2000 ;
	    RECT 95.8000 21.1000 96.2000 25.8000 ;
	    RECT 97.8000 25.6000 98.2000 25.8000 ;
	    RECT 99.8000 25.1000 100.1000 25.8000 ;
	    RECT 97.4000 24.8000 99.4000 25.1000 ;
	    RECT 97.4000 21.1000 97.8000 24.8000 ;
	    RECT 99.0000 21.1000 99.4000 24.8000 ;
	    RECT 99.8000 21.1000 100.2000 25.1000 ;
	    RECT 101.4000 21.1000 101.8000 27.9000 ;
	    RECT 103.0000 26.1000 103.4000 29.9000 ;
	    RECT 104.6000 28.0000 105.0000 29.9000 ;
	    RECT 106.2000 28.0000 106.6000 29.9000 ;
	    RECT 104.6000 27.9000 106.6000 28.0000 ;
	    RECT 107.0000 28.1000 107.4000 29.9000 ;
	    RECT 108.6000 28.8000 109.0000 29.2000 ;
	    RECT 108.6000 28.1000 108.9000 28.8000 ;
	    RECT 104.7000 27.7000 106.5000 27.9000 ;
	    RECT 107.0000 27.8000 108.9000 28.1000 ;
	    RECT 111.0000 27.9000 111.4000 29.9000 ;
	    RECT 111.7000 28.2000 112.1000 28.6000 ;
	    RECT 103.8000 26.8000 104.2000 27.6000 ;
	    RECT 105.0000 27.2000 105.4000 27.4000 ;
	    RECT 107.0000 27.2000 107.3000 27.8000 ;
	    RECT 104.6000 26.9000 105.4000 27.2000 ;
	    RECT 104.6000 26.8000 105.0000 26.9000 ;
	    RECT 106.1000 26.8000 107.4000 27.2000 ;
	    RECT 104.6000 26.1000 104.9000 26.8000 ;
	    RECT 103.0000 25.8000 104.9000 26.1000 ;
	    RECT 105.4000 25.8000 105.8000 26.6000 ;
	    RECT 102.2000 24.4000 102.6000 25.2000 ;
	    RECT 103.0000 21.1000 103.4000 25.8000 ;
	    RECT 106.1000 25.1000 106.4000 26.8000 ;
	    RECT 110.2000 26.4000 110.6000 27.2000 ;
	    RECT 107.8000 26.1000 108.2000 26.2000 ;
	    RECT 109.4000 26.1000 109.8000 26.2000 ;
	    RECT 111.0000 26.1000 111.3000 27.9000 ;
	    RECT 111.8000 27.8000 112.2000 28.2000 ;
	    RECT 112.6000 27.5000 113.0000 29.9000 ;
	    RECT 114.8000 29.2000 115.2000 29.9000 ;
	    RECT 114.2000 28.9000 115.2000 29.2000 ;
	    RECT 117.0000 28.9000 117.4000 29.9000 ;
	    RECT 119.1000 29.2000 119.7000 29.9000 ;
	    RECT 119.0000 28.9000 119.7000 29.2000 ;
	    RECT 114.2000 28.5000 114.6000 28.9000 ;
	    RECT 117.0000 28.6000 117.3000 28.9000 ;
	    RECT 115.0000 28.2000 115.4000 28.6000 ;
	    RECT 115.9000 28.3000 117.3000 28.6000 ;
	    RECT 119.0000 28.5000 119.4000 28.9000 ;
	    RECT 115.9000 28.2000 116.3000 28.3000 ;
	    RECT 113.0000 27.1000 113.8000 27.2000 ;
	    RECT 115.1000 27.1000 115.4000 28.2000 ;
	    RECT 119.9000 27.7000 120.3000 27.8000 ;
	    RECT 121.4000 27.7000 121.8000 29.9000 ;
	    RECT 122.2000 27.8000 122.6000 28.6000 ;
	    RECT 119.9000 27.4000 121.8000 27.7000 ;
	    RECT 117.9000 27.1000 118.3000 27.2000 ;
	    RECT 113.0000 26.8000 118.5000 27.1000 ;
	    RECT 114.5000 26.7000 114.9000 26.8000 ;
	    RECT 113.7000 26.2000 114.1000 26.3000 ;
	    RECT 115.0000 26.2000 115.4000 26.3000 ;
	    RECT 118.2000 26.2000 118.5000 26.8000 ;
	    RECT 119.0000 26.4000 119.4000 26.5000 ;
	    RECT 111.8000 26.1000 112.2000 26.2000 ;
	    RECT 107.8000 25.8000 110.2000 26.1000 ;
	    RECT 111.0000 25.8000 112.2000 26.1000 ;
	    RECT 113.7000 25.9000 116.2000 26.2000 ;
	    RECT 115.8000 25.8000 116.2000 25.9000 ;
	    RECT 118.2000 25.8000 118.6000 26.2000 ;
	    RECT 119.0000 26.1000 120.9000 26.4000 ;
	    RECT 120.5000 26.0000 120.9000 26.1000 ;
	    RECT 109.8000 25.6000 110.2000 25.8000 ;
	    RECT 111.8000 25.2000 112.1000 25.8000 ;
	    RECT 112.6000 25.5000 115.4000 25.6000 ;
	    RECT 112.6000 25.4000 115.5000 25.5000 ;
	    RECT 112.6000 25.3000 117.5000 25.4000 ;
	    RECT 107.0000 25.1000 107.4000 25.2000 ;
	    RECT 105.9000 24.8000 106.4000 25.1000 ;
	    RECT 106.7000 24.8000 107.4000 25.1000 ;
	    RECT 109.4000 24.8000 111.4000 25.1000 ;
	    RECT 105.9000 21.1000 106.3000 24.8000 ;
	    RECT 106.7000 24.2000 107.0000 24.8000 ;
	    RECT 106.6000 23.8000 107.0000 24.2000 ;
	    RECT 109.4000 21.1000 109.8000 24.8000 ;
	    RECT 111.0000 21.1000 111.4000 24.8000 ;
	    RECT 111.8000 21.1000 112.2000 25.2000 ;
	    RECT 112.6000 21.1000 113.0000 25.3000 ;
	    RECT 115.1000 25.1000 117.5000 25.3000 ;
	    RECT 114.2000 24.5000 116.9000 24.8000 ;
	    RECT 114.2000 24.4000 114.6000 24.5000 ;
	    RECT 116.5000 24.4000 116.9000 24.5000 ;
	    RECT 117.2000 24.5000 117.5000 25.1000 ;
	    RECT 118.2000 25.2000 118.5000 25.8000 ;
	    RECT 119.7000 25.7000 120.1000 25.8000 ;
	    RECT 121.4000 25.7000 121.8000 27.4000 ;
	    RECT 119.7000 25.4000 121.8000 25.7000 ;
	    RECT 118.2000 24.9000 119.4000 25.2000 ;
	    RECT 117.9000 24.5000 118.3000 24.6000 ;
	    RECT 117.2000 24.2000 118.3000 24.5000 ;
	    RECT 119.1000 24.4000 119.4000 24.9000 ;
	    RECT 119.1000 24.0000 119.8000 24.4000 ;
	    RECT 115.9000 23.7000 116.3000 23.8000 ;
	    RECT 117.3000 23.7000 117.7000 23.8000 ;
	    RECT 114.2000 23.1000 114.6000 23.5000 ;
	    RECT 115.9000 23.4000 117.7000 23.7000 ;
	    RECT 117.0000 23.1000 117.3000 23.4000 ;
	    RECT 119.0000 23.1000 119.4000 23.5000 ;
	    RECT 114.2000 22.8000 115.2000 23.1000 ;
	    RECT 114.8000 21.1000 115.2000 22.8000 ;
	    RECT 117.0000 21.1000 117.4000 23.1000 ;
	    RECT 119.1000 21.1000 119.7000 23.1000 ;
	    RECT 121.4000 21.1000 121.8000 25.4000 ;
	    RECT 123.0000 25.1000 123.4000 29.9000 ;
	    RECT 124.1000 29.2000 124.5000 29.9000 ;
	    RECT 123.8000 28.8000 124.5000 29.2000 ;
	    RECT 127.0000 28.9000 127.4000 29.9000 ;
	    RECT 124.1000 28.2000 124.5000 28.8000 ;
	    RECT 124.1000 27.9000 125.0000 28.2000 ;
	    RECT 123.8000 25.1000 124.2000 25.2000 ;
	    RECT 123.0000 24.8000 124.2000 25.1000 ;
	    RECT 123.0000 21.1000 123.4000 24.8000 ;
	    RECT 123.8000 24.4000 124.2000 24.8000 ;
	    RECT 124.6000 21.1000 125.0000 27.9000 ;
	    RECT 126.2000 27.8000 126.6000 28.6000 ;
	    RECT 127.1000 28.1000 127.4000 28.9000 ;
	    RECT 127.8000 28.1000 128.2000 28.2000 ;
	    RECT 127.0000 27.8000 128.2000 28.1000 ;
	    RECT 128.6000 27.9000 129.0000 29.9000 ;
	    RECT 130.2000 28.9000 130.6000 29.9000 ;
	    RECT 125.4000 26.8000 125.8000 27.6000 ;
	    RECT 127.1000 27.2000 127.4000 27.8000 ;
	    RECT 127.0000 26.8000 127.4000 27.2000 ;
	    RECT 126.2000 26.1000 126.6000 26.2000 ;
	    RECT 127.1000 26.1000 127.4000 26.8000 ;
	    RECT 128.6000 26.2000 128.9000 27.9000 ;
	    RECT 130.2000 27.8000 130.5000 28.9000 ;
	    RECT 132.6000 28.8000 133.0000 29.9000 ;
	    RECT 131.0000 27.8000 131.4000 28.6000 ;
	    RECT 131.8000 27.8000 132.2000 28.6000 ;
	    RECT 129.3000 27.5000 130.5000 27.8000 ;
	    RECT 126.2000 25.8000 127.4000 26.1000 ;
	    RECT 127.1000 25.1000 127.4000 25.8000 ;
	    RECT 127.8000 25.4000 128.2000 26.2000 ;
	    RECT 128.6000 25.8000 129.0000 26.2000 ;
	    RECT 129.3000 26.0000 129.6000 27.5000 ;
	    RECT 132.7000 27.2000 133.0000 28.8000 ;
	    RECT 134.5000 28.2000 134.9000 29.9000 ;
	    RECT 134.5000 27.9000 135.4000 28.2000 ;
	    RECT 136.6000 27.9000 137.0000 29.9000 ;
	    RECT 137.4000 28.0000 137.8000 29.9000 ;
	    RECT 139.0000 28.0000 139.4000 29.9000 ;
	    RECT 137.4000 27.9000 139.4000 28.0000 ;
	    RECT 130.1000 27.1000 130.6000 27.2000 ;
	    RECT 131.0000 27.1000 131.4000 27.2000 ;
	    RECT 130.1000 26.8000 131.4000 27.1000 ;
	    RECT 132.6000 26.8000 133.0000 27.2000 ;
	    RECT 130.0000 26.4000 130.4000 26.8000 ;
	    RECT 128.6000 25.1000 128.9000 25.8000 ;
	    RECT 129.3000 25.7000 129.7000 26.0000 ;
	    RECT 129.3000 25.6000 131.4000 25.7000 ;
	    RECT 129.4000 25.4000 131.4000 25.6000 ;
	    RECT 127.0000 24.7000 127.9000 25.1000 ;
	    RECT 128.6000 24.8000 129.3000 25.1000 ;
	    RECT 127.5000 21.1000 127.9000 24.7000 ;
	    RECT 128.9000 21.1000 129.3000 24.8000 ;
	    RECT 131.0000 21.1000 131.4000 25.4000 ;
	    RECT 132.7000 25.1000 133.0000 26.8000 ;
	    RECT 133.4000 26.1000 133.8000 26.2000 ;
	    RECT 134.2000 26.1000 134.6000 26.2000 ;
	    RECT 133.4000 25.8000 134.6000 26.1000 ;
	    RECT 135.0000 26.1000 135.4000 27.9000 ;
	    RECT 135.8000 26.8000 136.2000 27.6000 ;
	    RECT 136.7000 27.2000 137.0000 27.9000 ;
	    RECT 137.5000 27.7000 139.3000 27.9000 ;
	    RECT 138.6000 27.2000 139.0000 27.4000 ;
	    RECT 136.6000 26.8000 137.9000 27.2000 ;
	    RECT 138.6000 26.9000 139.4000 27.2000 ;
	    RECT 139.0000 26.8000 139.4000 26.9000 ;
	    RECT 135.8000 26.1000 136.2000 26.2000 ;
	    RECT 135.0000 25.8000 136.2000 26.1000 ;
	    RECT 133.4000 25.4000 133.8000 25.8000 ;
	    RECT 132.6000 24.7000 133.5000 25.1000 ;
	    RECT 133.1000 24.1000 133.5000 24.7000 ;
	    RECT 134.2000 24.1000 134.6000 25.2000 ;
	    RECT 133.1000 23.8000 134.6000 24.1000 ;
	    RECT 133.1000 21.1000 133.5000 23.8000 ;
	    RECT 135.0000 21.1000 135.4000 25.8000 ;
	    RECT 137.6000 25.2000 137.9000 26.8000 ;
	    RECT 138.2000 26.1000 138.6000 26.6000 ;
	    RECT 139.8000 26.1000 140.2000 29.9000 ;
	    RECT 140.6000 27.8000 141.0000 28.6000 ;
	    RECT 138.2000 25.8000 140.2000 26.1000 ;
	    RECT 136.6000 25.1000 137.0000 25.2000 ;
	    RECT 136.6000 24.8000 137.3000 25.1000 ;
	    RECT 137.6000 24.8000 138.6000 25.2000 ;
	    RECT 137.0000 24.2000 137.3000 24.8000 ;
	    RECT 137.0000 23.8000 137.4000 24.2000 ;
	    RECT 137.7000 21.1000 138.1000 24.8000 ;
	    RECT 139.8000 21.1000 140.2000 25.8000 ;
	    RECT 141.4000 27.7000 141.8000 29.9000 ;
	    RECT 143.5000 29.2000 144.1000 29.9000 ;
	    RECT 143.5000 28.9000 144.2000 29.2000 ;
	    RECT 145.8000 28.9000 146.2000 29.9000 ;
	    RECT 148.0000 29.2000 148.4000 29.9000 ;
	    RECT 148.0000 28.9000 149.0000 29.2000 ;
	    RECT 143.8000 28.5000 144.2000 28.9000 ;
	    RECT 145.9000 28.6000 146.2000 28.9000 ;
	    RECT 145.9000 28.3000 147.3000 28.6000 ;
	    RECT 146.9000 28.2000 147.3000 28.3000 ;
	    RECT 147.8000 28.2000 148.2000 28.6000 ;
	    RECT 148.6000 28.5000 149.0000 28.9000 ;
	    RECT 142.9000 27.7000 143.3000 27.8000 ;
	    RECT 141.4000 27.4000 143.3000 27.7000 ;
	    RECT 141.4000 25.7000 141.8000 27.4000 ;
	    RECT 144.9000 27.1000 145.8000 27.2000 ;
	    RECT 147.8000 27.1000 148.1000 28.2000 ;
	    RECT 150.2000 27.5000 150.6000 29.9000 ;
	    RECT 152.6000 27.9000 153.0000 29.9000 ;
	    RECT 153.3000 28.2000 153.7000 28.6000 ;
	    RECT 149.4000 27.1000 150.2000 27.2000 ;
	    RECT 144.7000 26.8000 150.2000 27.1000 ;
	    RECT 143.8000 26.4000 144.2000 26.5000 ;
	    RECT 142.3000 26.1000 144.2000 26.4000 ;
	    RECT 142.3000 26.0000 142.7000 26.1000 ;
	    RECT 143.1000 25.7000 143.5000 25.8000 ;
	    RECT 141.4000 25.4000 143.5000 25.7000 ;
	    RECT 141.4000 21.1000 141.8000 25.4000 ;
	    RECT 144.7000 25.2000 145.0000 26.8000 ;
	    RECT 148.3000 26.7000 148.7000 26.8000 ;
	    RECT 151.8000 26.4000 152.2000 27.2000 ;
	    RECT 149.1000 26.2000 149.5000 26.3000 ;
	    RECT 147.0000 25.9000 149.5000 26.2000 ;
	    RECT 151.0000 26.1000 151.4000 26.2000 ;
	    RECT 152.6000 26.1000 152.9000 27.9000 ;
	    RECT 153.4000 27.8000 153.8000 28.2000 ;
	    RECT 154.2000 27.5000 154.6000 29.9000 ;
	    RECT 156.4000 29.2000 156.8000 29.9000 ;
	    RECT 155.8000 28.9000 156.8000 29.2000 ;
	    RECT 158.6000 28.9000 159.0000 29.9000 ;
	    RECT 160.7000 29.2000 161.3000 29.9000 ;
	    RECT 160.6000 28.9000 161.3000 29.2000 ;
	    RECT 155.8000 28.5000 156.2000 28.9000 ;
	    RECT 158.6000 28.6000 158.9000 28.9000 ;
	    RECT 156.6000 28.2000 157.0000 28.6000 ;
	    RECT 157.5000 28.3000 158.9000 28.6000 ;
	    RECT 160.6000 28.5000 161.0000 28.9000 ;
	    RECT 157.5000 28.2000 157.9000 28.3000 ;
	    RECT 153.4000 27.1000 153.8000 27.2000 ;
	    RECT 154.6000 27.1000 155.4000 27.2000 ;
	    RECT 156.7000 27.1000 157.0000 28.2000 ;
	    RECT 161.5000 27.7000 161.9000 27.8000 ;
	    RECT 163.0000 27.7000 163.4000 29.9000 ;
	    RECT 165.4000 28.0000 165.8000 29.9000 ;
	    RECT 167.0000 28.0000 167.4000 29.9000 ;
	    RECT 165.4000 27.9000 167.4000 28.0000 ;
	    RECT 167.8000 27.9000 168.2000 29.9000 ;
	    RECT 165.5000 27.7000 167.3000 27.9000 ;
	    RECT 161.5000 27.4000 163.4000 27.7000 ;
	    RECT 159.5000 27.1000 159.9000 27.2000 ;
	    RECT 153.4000 26.8000 160.1000 27.1000 ;
	    RECT 156.1000 26.7000 156.5000 26.8000 ;
	    RECT 155.3000 26.2000 155.7000 26.3000 ;
	    RECT 156.6000 26.2000 157.0000 26.3000 ;
	    RECT 153.4000 26.1000 153.8000 26.2000 ;
	    RECT 147.0000 25.8000 147.4000 25.9000 ;
	    RECT 151.0000 25.8000 151.8000 26.1000 ;
	    RECT 152.6000 25.8000 153.8000 26.1000 ;
	    RECT 155.3000 25.9000 157.8000 26.2000 ;
	    RECT 157.4000 25.8000 157.8000 25.9000 ;
	    RECT 159.0000 26.1000 159.4000 26.2000 ;
	    RECT 159.8000 26.1000 160.1000 26.8000 ;
	    RECT 160.6000 26.4000 161.0000 26.5000 ;
	    RECT 160.6000 26.1000 162.5000 26.4000 ;
	    RECT 159.0000 25.8000 160.1000 26.1000 ;
	    RECT 162.1000 26.0000 162.5000 26.1000 ;
	    RECT 151.4000 25.6000 151.8000 25.8000 ;
	    RECT 147.8000 25.5000 150.6000 25.6000 ;
	    RECT 147.7000 25.4000 150.6000 25.5000 ;
	    RECT 143.8000 24.9000 145.0000 25.2000 ;
	    RECT 145.7000 25.3000 150.6000 25.4000 ;
	    RECT 145.7000 25.1000 148.1000 25.3000 ;
	    RECT 143.8000 24.4000 144.1000 24.9000 ;
	    RECT 143.4000 24.0000 144.1000 24.4000 ;
	    RECT 144.9000 24.5000 145.3000 24.6000 ;
	    RECT 145.7000 24.5000 146.0000 25.1000 ;
	    RECT 144.9000 24.2000 146.0000 24.5000 ;
	    RECT 146.3000 24.5000 149.0000 24.8000 ;
	    RECT 146.3000 24.4000 146.7000 24.5000 ;
	    RECT 148.6000 24.4000 149.0000 24.5000 ;
	    RECT 145.5000 23.7000 145.9000 23.8000 ;
	    RECT 146.9000 23.7000 147.3000 23.8000 ;
	    RECT 143.8000 23.1000 144.2000 23.5000 ;
	    RECT 145.5000 23.4000 147.3000 23.7000 ;
	    RECT 145.9000 23.1000 146.2000 23.4000 ;
	    RECT 148.6000 23.1000 149.0000 23.5000 ;
	    RECT 143.5000 21.1000 144.1000 23.1000 ;
	    RECT 145.8000 21.1000 146.2000 23.1000 ;
	    RECT 148.0000 22.8000 149.0000 23.1000 ;
	    RECT 148.0000 21.1000 148.4000 22.8000 ;
	    RECT 150.2000 21.1000 150.6000 25.3000 ;
	    RECT 153.4000 25.1000 153.7000 25.8000 ;
	    RECT 154.2000 25.5000 157.0000 25.6000 ;
	    RECT 154.2000 25.4000 157.1000 25.5000 ;
	    RECT 154.2000 25.3000 159.1000 25.4000 ;
	    RECT 151.0000 24.8000 153.0000 25.1000 ;
	    RECT 151.0000 21.1000 151.4000 24.8000 ;
	    RECT 152.6000 21.1000 153.0000 24.8000 ;
	    RECT 153.4000 21.1000 153.8000 25.1000 ;
	    RECT 154.2000 21.1000 154.6000 25.3000 ;
	    RECT 156.7000 25.1000 159.1000 25.3000 ;
	    RECT 155.8000 24.5000 158.5000 24.8000 ;
	    RECT 155.8000 24.4000 156.2000 24.5000 ;
	    RECT 158.1000 24.4000 158.5000 24.5000 ;
	    RECT 158.8000 24.5000 159.1000 25.1000 ;
	    RECT 159.8000 25.2000 160.1000 25.8000 ;
	    RECT 161.3000 25.7000 161.7000 25.8000 ;
	    RECT 163.0000 25.7000 163.4000 27.4000 ;
	    RECT 165.8000 27.2000 166.2000 27.4000 ;
	    RECT 167.8000 27.2000 168.1000 27.9000 ;
	    RECT 168.6000 27.5000 169.0000 29.9000 ;
	    RECT 170.8000 29.2000 171.2000 29.9000 ;
	    RECT 170.2000 28.9000 171.2000 29.2000 ;
	    RECT 173.0000 28.9000 173.4000 29.9000 ;
	    RECT 175.1000 29.2000 175.7000 29.9000 ;
	    RECT 175.0000 28.9000 175.7000 29.2000 ;
	    RECT 170.2000 28.5000 170.6000 28.9000 ;
	    RECT 173.0000 28.6000 173.3000 28.9000 ;
	    RECT 171.0000 28.2000 171.4000 28.6000 ;
	    RECT 171.9000 28.3000 173.3000 28.6000 ;
	    RECT 175.0000 28.5000 175.4000 28.9000 ;
	    RECT 171.9000 28.2000 172.3000 28.3000 ;
	    RECT 165.4000 26.9000 166.2000 27.2000 ;
	    RECT 165.4000 26.8000 165.8000 26.9000 ;
	    RECT 166.9000 26.8000 168.2000 27.2000 ;
	    RECT 169.0000 27.1000 169.8000 27.2000 ;
	    RECT 171.1000 27.1000 171.4000 28.2000 ;
	    RECT 175.9000 27.7000 176.3000 27.8000 ;
	    RECT 177.4000 27.7000 177.8000 29.9000 ;
	    RECT 179.0000 28.9000 179.4000 29.9000 ;
	    RECT 178.2000 27.8000 178.6000 28.6000 ;
	    RECT 175.9000 27.4000 177.8000 27.7000 ;
	    RECT 173.9000 27.1000 174.3000 27.2000 ;
	    RECT 169.0000 26.8000 174.5000 27.1000 ;
	    RECT 166.2000 25.8000 166.6000 26.6000 ;
	    RECT 161.3000 25.4000 163.4000 25.7000 ;
	    RECT 159.8000 24.9000 161.0000 25.2000 ;
	    RECT 159.5000 24.5000 159.9000 24.6000 ;
	    RECT 158.8000 24.2000 159.9000 24.5000 ;
	    RECT 160.7000 24.4000 161.0000 24.9000 ;
	    RECT 160.7000 24.0000 161.4000 24.4000 ;
	    RECT 157.5000 23.7000 157.9000 23.8000 ;
	    RECT 158.9000 23.7000 159.3000 23.8000 ;
	    RECT 155.8000 23.1000 156.2000 23.5000 ;
	    RECT 157.5000 23.4000 159.3000 23.7000 ;
	    RECT 158.6000 23.1000 158.9000 23.4000 ;
	    RECT 160.6000 23.1000 161.0000 23.5000 ;
	    RECT 155.8000 22.8000 156.8000 23.1000 ;
	    RECT 156.4000 21.1000 156.8000 22.8000 ;
	    RECT 158.6000 21.1000 159.0000 23.1000 ;
	    RECT 160.7000 21.1000 161.3000 23.1000 ;
	    RECT 163.0000 21.1000 163.4000 25.4000 ;
	    RECT 166.9000 25.1000 167.2000 26.8000 ;
	    RECT 170.5000 26.7000 170.9000 26.8000 ;
	    RECT 169.7000 26.2000 170.1000 26.3000 ;
	    RECT 169.7000 25.9000 172.2000 26.2000 ;
	    RECT 171.8000 25.8000 172.2000 25.9000 ;
	    RECT 168.6000 25.5000 171.4000 25.6000 ;
	    RECT 168.6000 25.4000 171.5000 25.5000 ;
	    RECT 168.6000 25.3000 173.5000 25.4000 ;
	    RECT 167.8000 25.1000 168.2000 25.2000 ;
	    RECT 166.7000 24.8000 167.2000 25.1000 ;
	    RECT 167.5000 24.8000 168.2000 25.1000 ;
	    RECT 166.7000 21.1000 167.1000 24.8000 ;
	    RECT 167.5000 24.2000 167.8000 24.8000 ;
	    RECT 167.4000 23.8000 167.8000 24.2000 ;
	    RECT 168.6000 21.1000 169.0000 25.3000 ;
	    RECT 171.1000 25.1000 173.5000 25.3000 ;
	    RECT 170.2000 24.5000 172.9000 24.8000 ;
	    RECT 170.2000 24.4000 170.6000 24.5000 ;
	    RECT 172.5000 24.4000 172.9000 24.5000 ;
	    RECT 173.2000 24.5000 173.5000 25.1000 ;
	    RECT 174.2000 25.2000 174.5000 26.8000 ;
	    RECT 175.0000 26.4000 175.4000 26.5000 ;
	    RECT 175.0000 26.1000 176.9000 26.4000 ;
	    RECT 176.5000 26.0000 176.9000 26.1000 ;
	    RECT 175.7000 25.7000 176.1000 25.8000 ;
	    RECT 177.4000 25.7000 177.8000 27.4000 ;
	    RECT 179.1000 27.2000 179.4000 28.9000 ;
	    RECT 179.0000 26.8000 179.4000 27.2000 ;
	    RECT 175.7000 25.4000 177.8000 25.7000 ;
	    RECT 174.2000 24.9000 175.4000 25.2000 ;
	    RECT 173.9000 24.5000 174.3000 24.6000 ;
	    RECT 173.2000 24.2000 174.3000 24.5000 ;
	    RECT 175.1000 24.4000 175.4000 24.9000 ;
	    RECT 175.1000 24.0000 175.8000 24.4000 ;
	    RECT 171.9000 23.7000 172.3000 23.8000 ;
	    RECT 173.3000 23.7000 173.7000 23.8000 ;
	    RECT 170.2000 23.1000 170.6000 23.5000 ;
	    RECT 171.9000 23.4000 173.7000 23.7000 ;
	    RECT 173.0000 23.1000 173.3000 23.4000 ;
	    RECT 175.0000 23.1000 175.4000 23.5000 ;
	    RECT 170.2000 22.8000 171.2000 23.1000 ;
	    RECT 170.8000 21.1000 171.2000 22.8000 ;
	    RECT 173.0000 21.1000 173.4000 23.1000 ;
	    RECT 175.1000 21.1000 175.7000 23.1000 ;
	    RECT 177.4000 21.1000 177.8000 25.4000 ;
	    RECT 179.1000 25.1000 179.4000 26.8000 ;
	    RECT 179.8000 26.1000 180.2000 26.2000 ;
	    RECT 180.6000 26.1000 181.0000 29.9000 ;
	    RECT 181.4000 27.8000 181.8000 28.6000 ;
	    RECT 183.0000 27.6000 183.4000 29.9000 ;
	    RECT 184.6000 27.6000 185.0000 29.9000 ;
	    RECT 186.2000 27.6000 186.6000 29.9000 ;
	    RECT 187.8000 27.6000 188.2000 29.9000 ;
	    RECT 183.0000 27.2000 183.9000 27.6000 ;
	    RECT 184.6000 27.2000 185.7000 27.6000 ;
	    RECT 186.2000 27.2000 187.3000 27.6000 ;
	    RECT 187.8000 27.2000 189.0000 27.6000 ;
	    RECT 189.4000 27.5000 189.8000 29.9000 ;
	    RECT 191.6000 29.2000 192.0000 29.9000 ;
	    RECT 191.0000 28.9000 192.0000 29.2000 ;
	    RECT 193.8000 28.9000 194.2000 29.9000 ;
	    RECT 195.9000 29.2000 196.5000 29.9000 ;
	    RECT 195.8000 28.9000 196.5000 29.2000 ;
	    RECT 191.0000 28.5000 191.4000 28.9000 ;
	    RECT 193.8000 28.6000 194.1000 28.9000 ;
	    RECT 191.8000 28.2000 192.2000 28.6000 ;
	    RECT 192.7000 28.3000 194.1000 28.6000 ;
	    RECT 195.8000 28.5000 196.2000 28.9000 ;
	    RECT 192.7000 28.2000 193.1000 28.3000 ;
	    RECT 191.9000 27.2000 192.2000 28.2000 ;
	    RECT 196.7000 27.7000 197.1000 27.8000 ;
	    RECT 198.2000 27.7000 198.6000 29.9000 ;
	    RECT 196.7000 27.4000 198.6000 27.7000 ;
	    RECT 179.8000 25.8000 181.0000 26.1000 ;
	    RECT 183.5000 26.9000 183.9000 27.2000 ;
	    RECT 185.3000 26.9000 185.7000 27.2000 ;
	    RECT 186.9000 26.9000 187.3000 27.2000 ;
	    RECT 183.5000 26.5000 184.8000 26.9000 ;
	    RECT 185.3000 26.5000 186.5000 26.9000 ;
	    RECT 186.9000 26.5000 188.2000 26.9000 ;
	    RECT 183.5000 25.8000 183.9000 26.5000 ;
	    RECT 185.3000 25.8000 185.7000 26.5000 ;
	    RECT 186.9000 25.8000 187.3000 26.5000 ;
	    RECT 188.6000 25.8000 189.0000 27.2000 ;
	    RECT 189.8000 27.1000 190.6000 27.2000 ;
	    RECT 191.8000 27.1000 192.2000 27.2000 ;
	    RECT 194.7000 27.1000 195.4000 27.2000 ;
	    RECT 189.8000 26.8000 195.4000 27.1000 ;
	    RECT 198.2000 27.1000 198.6000 27.4000 ;
	    RECT 199.0000 27.1000 199.4000 27.6000 ;
	    RECT 198.2000 26.8000 199.4000 27.1000 ;
	    RECT 191.3000 26.7000 191.7000 26.8000 ;
	    RECT 190.5000 26.2000 190.9000 26.3000 ;
	    RECT 190.5000 25.9000 193.0000 26.2000 ;
	    RECT 192.6000 25.8000 193.0000 25.9000 ;
	    RECT 179.8000 25.4000 180.2000 25.8000 ;
	    RECT 179.0000 24.7000 179.9000 25.1000 ;
	    RECT 179.5000 24.2000 179.9000 24.7000 ;
	    RECT 179.5000 23.8000 180.2000 24.2000 ;
	    RECT 179.5000 21.1000 179.9000 23.8000 ;
	    RECT 180.6000 21.1000 181.0000 25.8000 ;
	    RECT 183.0000 25.4000 183.9000 25.8000 ;
	    RECT 184.6000 25.4000 185.7000 25.8000 ;
	    RECT 186.2000 25.4000 187.3000 25.8000 ;
	    RECT 187.8000 25.4000 189.0000 25.8000 ;
	    RECT 189.4000 25.5000 192.2000 25.6000 ;
	    RECT 189.4000 25.4000 192.3000 25.5000 ;
	    RECT 183.0000 21.1000 183.4000 25.4000 ;
	    RECT 184.6000 21.1000 185.0000 25.4000 ;
	    RECT 186.2000 21.1000 186.6000 25.4000 ;
	    RECT 187.8000 21.1000 188.2000 25.4000 ;
	    RECT 189.4000 25.3000 194.3000 25.4000 ;
	    RECT 189.4000 21.1000 189.8000 25.3000 ;
	    RECT 191.9000 25.1000 194.3000 25.3000 ;
	    RECT 191.0000 24.5000 193.7000 24.8000 ;
	    RECT 191.0000 24.4000 191.4000 24.5000 ;
	    RECT 193.3000 24.4000 193.7000 24.5000 ;
	    RECT 194.0000 24.5000 194.3000 25.1000 ;
	    RECT 195.0000 25.2000 195.3000 26.8000 ;
	    RECT 195.8000 26.4000 196.2000 26.5000 ;
	    RECT 195.8000 26.1000 197.7000 26.4000 ;
	    RECT 197.3000 26.0000 197.7000 26.1000 ;
	    RECT 196.5000 25.7000 196.9000 25.8000 ;
	    RECT 198.2000 25.7000 198.6000 26.8000 ;
	    RECT 196.5000 25.4000 198.6000 25.7000 ;
	    RECT 195.0000 24.9000 196.2000 25.2000 ;
	    RECT 194.7000 24.5000 195.1000 24.6000 ;
	    RECT 194.0000 24.2000 195.1000 24.5000 ;
	    RECT 195.9000 24.4000 196.2000 24.9000 ;
	    RECT 195.9000 24.0000 196.6000 24.4000 ;
	    RECT 192.7000 23.7000 193.1000 23.8000 ;
	    RECT 194.1000 23.7000 194.5000 23.8000 ;
	    RECT 191.0000 23.1000 191.4000 23.5000 ;
	    RECT 192.7000 23.4000 194.5000 23.7000 ;
	    RECT 193.8000 23.1000 194.1000 23.4000 ;
	    RECT 195.8000 23.1000 196.2000 23.5000 ;
	    RECT 191.0000 22.8000 192.0000 23.1000 ;
	    RECT 191.6000 21.1000 192.0000 22.8000 ;
	    RECT 193.8000 21.1000 194.2000 23.1000 ;
	    RECT 195.9000 21.1000 196.5000 23.1000 ;
	    RECT 198.2000 21.1000 198.6000 25.4000 ;
	    RECT 199.8000 26.1000 200.2000 29.9000 ;
	    RECT 202.5000 28.0000 202.9000 29.5000 ;
	    RECT 204.6000 28.5000 205.0000 29.5000 ;
	    RECT 205.7000 29.2000 206.1000 29.9000 ;
	    RECT 205.4000 28.8000 206.1000 29.2000 ;
	    RECT 202.1000 27.7000 202.9000 28.0000 ;
	    RECT 202.1000 27.5000 202.5000 27.7000 ;
	    RECT 202.1000 27.2000 202.4000 27.5000 ;
	    RECT 204.7000 27.4000 205.0000 28.5000 ;
	    RECT 205.7000 28.4000 206.1000 28.8000 ;
	    RECT 200.6000 27.1000 201.0000 27.2000 ;
	    RECT 201.4000 27.1000 202.4000 27.2000 ;
	    RECT 200.6000 26.8000 202.4000 27.1000 ;
	    RECT 202.9000 27.1000 205.0000 27.4000 ;
	    RECT 205.4000 27.9000 206.1000 28.4000 ;
	    RECT 207.8000 27.9000 208.2000 29.9000 ;
	    RECT 208.6000 28.0000 209.0000 29.9000 ;
	    RECT 210.2000 28.0000 210.6000 29.9000 ;
	    RECT 208.6000 27.9000 210.6000 28.0000 ;
	    RECT 211.0000 27.9000 211.4000 29.9000 ;
	    RECT 202.9000 26.9000 203.4000 27.1000 ;
	    RECT 201.4000 26.1000 201.8000 26.2000 ;
	    RECT 199.8000 25.8000 201.8000 26.1000 ;
	    RECT 199.8000 21.1000 200.2000 25.8000 ;
	    RECT 201.4000 25.4000 201.8000 25.8000 ;
	    RECT 202.1000 24.9000 202.4000 26.8000 ;
	    RECT 202.7000 26.5000 203.4000 26.9000 ;
	    RECT 203.1000 25.5000 203.4000 26.5000 ;
	    RECT 203.8000 25.8000 204.2000 26.6000 ;
	    RECT 204.6000 25.8000 205.0000 26.6000 ;
	    RECT 205.4000 26.2000 205.7000 27.9000 ;
	    RECT 207.8000 27.8000 208.1000 27.9000 ;
	    RECT 207.2000 27.6000 208.1000 27.8000 ;
	    RECT 208.7000 27.7000 210.5000 27.9000 ;
	    RECT 206.0000 27.5000 208.1000 27.6000 ;
	    RECT 206.0000 27.3000 207.5000 27.5000 ;
	    RECT 206.0000 27.2000 206.4000 27.3000 ;
	    RECT 209.0000 27.2000 209.4000 27.4000 ;
	    RECT 211.0000 27.2000 211.3000 27.9000 ;
	    RECT 205.4000 25.8000 205.8000 26.2000 ;
	    RECT 203.1000 25.2000 205.0000 25.5000 ;
	    RECT 202.1000 24.6000 202.9000 24.9000 ;
	    RECT 202.5000 21.1000 202.9000 24.6000 ;
	    RECT 204.7000 23.5000 205.0000 25.2000 ;
	    RECT 204.6000 21.5000 205.0000 23.5000 ;
	    RECT 205.4000 25.1000 205.7000 25.8000 ;
	    RECT 206.1000 25.5000 206.4000 27.2000 ;
	    RECT 206.8000 26.9000 207.2000 27.0000 ;
	    RECT 206.8000 26.6000 207.3000 26.9000 ;
	    RECT 207.0000 26.2000 207.3000 26.6000 ;
	    RECT 207.8000 26.4000 208.2000 27.2000 ;
	    RECT 208.6000 26.9000 209.4000 27.2000 ;
	    RECT 208.6000 26.8000 209.0000 26.9000 ;
	    RECT 210.1000 26.8000 211.4000 27.2000 ;
	    RECT 207.0000 25.8000 207.4000 26.2000 ;
	    RECT 209.4000 25.8000 209.8000 26.6000 ;
	    RECT 206.1000 25.2000 207.3000 25.5000 ;
	    RECT 205.4000 21.1000 205.8000 25.1000 ;
	    RECT 207.0000 23.1000 207.3000 25.2000 ;
	    RECT 210.1000 25.1000 210.4000 26.8000 ;
	    RECT 211.0000 25.1000 211.4000 25.2000 ;
	    RECT 209.9000 24.8000 210.4000 25.1000 ;
	    RECT 210.7000 24.8000 211.4000 25.1000 ;
	    RECT 212.6000 25.1000 213.0000 25.2000 ;
	    RECT 213.4000 25.1000 213.8000 29.9000 ;
	    RECT 215.3000 29.2000 215.7000 29.9000 ;
	    RECT 215.3000 28.8000 216.2000 29.2000 ;
	    RECT 214.2000 27.8000 214.6000 28.6000 ;
	    RECT 215.3000 28.2000 215.7000 28.8000 ;
	    RECT 218.7000 28.2000 219.1000 29.9000 ;
	    RECT 215.3000 27.9000 216.2000 28.2000 ;
	    RECT 212.6000 24.8000 213.8000 25.1000 ;
	    RECT 207.0000 21.1000 207.4000 23.1000 ;
	    RECT 209.9000 21.1000 210.3000 24.8000 ;
	    RECT 210.7000 24.2000 211.0000 24.8000 ;
	    RECT 210.6000 23.8000 211.0000 24.2000 ;
	    RECT 213.4000 21.1000 213.8000 24.8000 ;
	    RECT 215.0000 24.4000 215.4000 25.2000 ;
	    RECT 215.8000 21.1000 216.2000 27.9000 ;
	    RECT 218.2000 27.9000 219.1000 28.2000 ;
	    RECT 216.6000 26.8000 217.0000 27.6000 ;
	    RECT 217.4000 26.8000 217.8000 27.6000 ;
	    RECT 218.2000 26.1000 218.6000 27.9000 ;
	    RECT 219.0000 27.1000 219.4000 27.2000 ;
	    RECT 219.8000 27.1000 220.2000 29.9000 ;
	    RECT 222.7000 29.2000 223.1000 29.9000 ;
	    RECT 222.7000 28.8000 223.4000 29.2000 ;
	    RECT 224.6000 28.9000 225.0000 29.9000 ;
	    RECT 222.7000 28.2000 223.1000 28.8000 ;
	    RECT 222.2000 27.9000 223.1000 28.2000 ;
	    RECT 219.0000 26.8000 220.2000 27.1000 ;
	    RECT 221.4000 26.8000 221.8000 27.6000 ;
	    RECT 219.0000 26.1000 219.4000 26.2000 ;
	    RECT 218.2000 25.8000 219.4000 26.1000 ;
	    RECT 218.2000 21.1000 218.6000 25.8000 ;
	    RECT 219.0000 25.1000 219.4000 25.2000 ;
	    RECT 219.8000 25.1000 220.2000 26.8000 ;
	    RECT 219.0000 24.8000 220.2000 25.1000 ;
	    RECT 219.0000 24.4000 219.4000 24.8000 ;
	    RECT 219.8000 21.1000 220.2000 24.8000 ;
	    RECT 222.2000 21.1000 222.6000 27.9000 ;
	    RECT 224.7000 27.2000 225.0000 28.9000 ;
	    RECT 226.2000 28.0000 226.6000 29.9000 ;
	    RECT 227.8000 28.0000 228.2000 29.9000 ;
	    RECT 226.2000 27.9000 228.2000 28.0000 ;
	    RECT 226.3000 27.7000 228.1000 27.9000 ;
	    RECT 228.6000 27.8000 229.0000 29.9000 ;
	    RECT 231.0000 27.9000 231.4000 29.9000 ;
	    RECT 232.9000 29.2000 233.3000 29.9000 ;
	    RECT 232.6000 28.8000 233.3000 29.2000 ;
	    RECT 231.7000 28.2000 232.1000 28.6000 ;
	    RECT 232.9000 28.2000 233.3000 28.8000 ;
	    RECT 226.6000 27.2000 227.0000 27.4000 ;
	    RECT 228.6000 27.2000 228.9000 27.8000 ;
	    RECT 224.6000 26.8000 225.0000 27.2000 ;
	    RECT 226.2000 26.9000 227.0000 27.2000 ;
	    RECT 226.2000 26.8000 226.6000 26.9000 ;
	    RECT 227.7000 26.8000 229.0000 27.2000 ;
	    RECT 224.7000 26.1000 225.0000 26.8000 ;
	    RECT 223.0000 25.8000 225.0000 26.1000 ;
	    RECT 223.0000 25.2000 223.3000 25.8000 ;
	    RECT 223.0000 24.4000 223.4000 25.2000 ;
	    RECT 224.7000 25.1000 225.0000 25.8000 ;
	    RECT 225.4000 25.4000 225.8000 26.2000 ;
	    RECT 227.0000 25.8000 227.4000 26.6000 ;
	    RECT 227.7000 25.1000 228.0000 26.8000 ;
	    RECT 230.2000 26.4000 230.6000 27.2000 ;
	    RECT 231.0000 27.1000 231.3000 27.9000 ;
	    RECT 231.8000 27.8000 232.2000 28.2000 ;
	    RECT 232.9000 27.9000 233.8000 28.2000 ;
	    RECT 235.0000 27.9000 235.4000 29.9000 ;
	    RECT 235.8000 28.0000 236.2000 29.9000 ;
	    RECT 237.4000 28.0000 237.8000 29.9000 ;
	    RECT 235.8000 27.9000 237.8000 28.0000 ;
	    RECT 239.8000 27.9000 240.2000 29.9000 ;
	    RECT 240.5000 28.2000 240.9000 28.6000 ;
	    RECT 232.6000 27.1000 233.0000 27.2000 ;
	    RECT 231.0000 26.8000 233.0000 27.1000 ;
	    RECT 228.6000 26.1000 229.0000 26.2000 ;
	    RECT 229.4000 26.1000 229.8000 26.2000 ;
	    RECT 231.0000 26.1000 231.3000 26.8000 ;
	    RECT 231.8000 26.1000 232.2000 26.2000 ;
	    RECT 228.6000 25.8000 230.2000 26.1000 ;
	    RECT 231.0000 25.8000 232.2000 26.1000 ;
	    RECT 229.8000 25.6000 230.2000 25.8000 ;
	    RECT 228.6000 25.1000 229.0000 25.2000 ;
	    RECT 231.8000 25.1000 232.1000 25.8000 ;
	    RECT 224.6000 24.7000 225.5000 25.1000 ;
	    RECT 225.1000 21.1000 225.5000 24.7000 ;
	    RECT 227.5000 24.8000 228.0000 25.1000 ;
	    RECT 228.3000 24.8000 229.0000 25.1000 ;
	    RECT 229.4000 24.8000 231.4000 25.1000 ;
	    RECT 227.5000 21.1000 227.9000 24.8000 ;
	    RECT 228.3000 24.2000 228.6000 24.8000 ;
	    RECT 228.2000 23.8000 228.6000 24.2000 ;
	    RECT 229.4000 21.1000 229.8000 24.8000 ;
	    RECT 231.0000 21.1000 231.4000 24.8000 ;
	    RECT 231.8000 21.1000 232.2000 25.1000 ;
	    RECT 232.6000 24.4000 233.0000 25.2000 ;
	    RECT 233.4000 21.1000 233.8000 27.9000 ;
	    RECT 234.2000 26.8000 234.6000 27.6000 ;
	    RECT 235.1000 27.2000 235.4000 27.9000 ;
	    RECT 235.9000 27.7000 237.7000 27.9000 ;
	    RECT 237.0000 27.2000 237.4000 27.4000 ;
	    RECT 235.0000 26.8000 236.3000 27.2000 ;
	    RECT 237.0000 26.9000 237.8000 27.2000 ;
	    RECT 237.4000 26.8000 237.8000 26.9000 ;
	    RECT 236.0000 25.2000 236.3000 26.8000 ;
	    RECT 236.6000 25.8000 237.0000 26.6000 ;
	    RECT 239.0000 26.4000 239.4000 27.2000 ;
	    RECT 238.2000 26.1000 238.6000 26.2000 ;
	    RECT 239.8000 26.1000 240.1000 27.9000 ;
	    RECT 240.6000 27.8000 241.0000 28.2000 ;
	    RECT 240.6000 26.1000 241.0000 26.2000 ;
	    RECT 238.2000 25.8000 239.0000 26.1000 ;
	    RECT 239.8000 25.8000 241.0000 26.1000 ;
	    RECT 238.6000 25.6000 239.0000 25.8000 ;
	    RECT 235.0000 25.1000 235.4000 25.2000 ;
	    RECT 235.0000 24.8000 235.7000 25.1000 ;
	    RECT 236.0000 24.8000 237.0000 25.2000 ;
	    RECT 240.6000 25.1000 240.9000 25.8000 ;
	    RECT 238.2000 24.8000 240.2000 25.1000 ;
	    RECT 235.4000 24.2000 235.7000 24.8000 ;
	    RECT 235.4000 23.8000 235.8000 24.2000 ;
	    RECT 236.1000 21.1000 236.5000 24.8000 ;
	    RECT 238.2000 21.1000 238.6000 24.8000 ;
	    RECT 239.8000 21.1000 240.2000 24.8000 ;
	    RECT 240.6000 21.1000 241.0000 25.1000 ;
	    RECT 242.2000 21.1000 242.6000 29.9000 ;
	    RECT 243.8000 27.9000 244.2000 29.9000 ;
	    RECT 246.0000 28.1000 246.8000 29.9000 ;
	    RECT 243.8000 27.6000 244.9000 27.9000 ;
	    RECT 245.4000 27.7000 246.2000 27.8000 ;
	    RECT 243.0000 26.8000 243.4000 27.6000 ;
	    RECT 244.5000 27.5000 244.9000 27.6000 ;
	    RECT 245.2000 27.4000 246.2000 27.7000 ;
	    RECT 245.2000 27.2000 245.5000 27.4000 ;
	    RECT 243.8000 26.9000 245.5000 27.2000 ;
	    RECT 243.8000 26.8000 244.6000 26.9000 ;
	    RECT 245.8000 26.7000 246.2000 27.1000 ;
	    RECT 245.8000 26.4000 246.1000 26.7000 ;
	    RECT 244.8000 26.1000 246.1000 26.4000 ;
	    RECT 246.5000 26.4000 246.8000 28.1000 ;
	    RECT 248.6000 27.9000 249.0000 29.9000 ;
	    RECT 247.1000 27.4000 247.5000 27.8000 ;
	    RECT 247.8000 27.6000 249.0000 27.9000 ;
	    RECT 247.8000 27.5000 248.2000 27.6000 ;
	    RECT 249.4000 27.5000 249.8000 29.9000 ;
	    RECT 251.6000 29.2000 252.0000 29.9000 ;
	    RECT 251.0000 28.9000 252.0000 29.2000 ;
	    RECT 253.8000 28.9000 254.2000 29.9000 ;
	    RECT 255.9000 29.2000 256.5000 29.9000 ;
	    RECT 255.8000 28.9000 256.5000 29.2000 ;
	    RECT 251.0000 28.5000 251.4000 28.9000 ;
	    RECT 253.8000 28.6000 254.1000 28.9000 ;
	    RECT 251.8000 28.2000 252.2000 28.6000 ;
	    RECT 252.7000 28.3000 254.1000 28.6000 ;
	    RECT 255.8000 28.5000 256.2000 28.9000 ;
	    RECT 252.7000 28.2000 253.1000 28.3000 ;
	    RECT 247.2000 27.2000 247.5000 27.4000 ;
	    RECT 247.2000 26.8000 247.6000 27.2000 ;
	    RECT 248.2000 26.8000 249.0000 27.2000 ;
	    RECT 249.8000 27.1000 250.6000 27.2000 ;
	    RECT 251.9000 27.1000 252.2000 28.2000 ;
	    RECT 255.0000 27.8000 255.4000 28.2000 ;
	    RECT 255.0000 27.2000 255.3000 27.8000 ;
	    RECT 256.7000 27.7000 257.1000 27.8000 ;
	    RECT 258.2000 27.7000 258.6000 29.9000 ;
	    RECT 259.0000 27.8000 259.4000 28.6000 ;
	    RECT 256.7000 27.4000 258.6000 27.7000 ;
	    RECT 254.7000 27.1000 255.3000 27.2000 ;
	    RECT 249.8000 26.8000 255.3000 27.1000 ;
	    RECT 251.3000 26.7000 251.7000 26.8000 ;
	    RECT 246.5000 26.2000 247.0000 26.4000 ;
	    RECT 250.5000 26.2000 250.9000 26.3000 ;
	    RECT 251.8000 26.2000 252.2000 26.3000 ;
	    RECT 246.5000 26.1000 247.4000 26.2000 ;
	    RECT 248.6000 26.1000 249.0000 26.2000 ;
	    RECT 244.8000 26.0000 245.2000 26.1000 ;
	    RECT 246.7000 25.8000 249.0000 26.1000 ;
	    RECT 250.5000 25.9000 253.0000 26.2000 ;
	    RECT 252.6000 25.8000 253.0000 25.9000 ;
	    RECT 245.9000 25.7000 246.3000 25.8000 ;
	    RECT 244.6000 25.4000 246.3000 25.7000 ;
	    RECT 244.6000 25.1000 244.9000 25.4000 ;
	    RECT 246.7000 25.1000 247.0000 25.8000 ;
	    RECT 249.4000 25.5000 252.2000 25.6000 ;
	    RECT 249.4000 25.4000 252.3000 25.5000 ;
	    RECT 249.4000 25.3000 254.3000 25.4000 ;
	    RECT 243.8000 24.8000 244.9000 25.1000 ;
	    RECT 243.8000 21.1000 244.2000 24.8000 ;
	    RECT 244.5000 24.7000 244.9000 24.8000 ;
	    RECT 246.0000 24.8000 247.0000 25.1000 ;
	    RECT 247.8000 24.8000 249.0000 25.1000 ;
	    RECT 246.0000 21.1000 246.8000 24.8000 ;
	    RECT 247.8000 24.7000 248.2000 24.8000 ;
	    RECT 248.6000 21.1000 249.0000 24.8000 ;
	    RECT 249.4000 21.1000 249.8000 25.3000 ;
	    RECT 251.9000 25.1000 254.3000 25.3000 ;
	    RECT 251.0000 24.5000 253.7000 24.8000 ;
	    RECT 251.0000 24.4000 251.4000 24.5000 ;
	    RECT 253.3000 24.4000 253.7000 24.5000 ;
	    RECT 254.0000 24.5000 254.3000 25.1000 ;
	    RECT 255.0000 25.2000 255.3000 26.8000 ;
	    RECT 255.8000 26.4000 256.2000 26.5000 ;
	    RECT 255.8000 26.1000 257.7000 26.4000 ;
	    RECT 257.3000 26.0000 257.7000 26.1000 ;
	    RECT 256.5000 25.7000 256.9000 25.8000 ;
	    RECT 258.2000 25.7000 258.6000 27.4000 ;
	    RECT 256.5000 25.4000 258.6000 25.7000 ;
	    RECT 255.0000 24.9000 256.2000 25.2000 ;
	    RECT 254.7000 24.5000 255.1000 24.6000 ;
	    RECT 254.0000 24.2000 255.1000 24.5000 ;
	    RECT 255.9000 24.4000 256.2000 24.9000 ;
	    RECT 255.9000 24.0000 256.6000 24.4000 ;
	    RECT 252.7000 23.7000 253.1000 23.8000 ;
	    RECT 254.1000 23.7000 254.5000 23.8000 ;
	    RECT 251.0000 23.1000 251.4000 23.5000 ;
	    RECT 252.7000 23.4000 254.5000 23.7000 ;
	    RECT 253.8000 23.1000 254.1000 23.4000 ;
	    RECT 255.8000 23.1000 256.2000 23.5000 ;
	    RECT 251.0000 22.8000 252.0000 23.1000 ;
	    RECT 251.6000 21.1000 252.0000 22.8000 ;
	    RECT 253.8000 21.1000 254.2000 23.1000 ;
	    RECT 255.9000 21.1000 256.5000 23.1000 ;
	    RECT 258.2000 21.1000 258.6000 25.4000 ;
	    RECT 259.8000 21.1000 260.2000 29.9000 ;
	    RECT 260.6000 27.5000 261.0000 29.9000 ;
	    RECT 262.8000 29.2000 263.2000 29.9000 ;
	    RECT 262.2000 28.9000 263.2000 29.2000 ;
	    RECT 265.0000 28.9000 265.4000 29.9000 ;
	    RECT 267.1000 29.2000 267.7000 29.9000 ;
	    RECT 267.0000 28.9000 267.7000 29.2000 ;
	    RECT 262.2000 28.5000 262.6000 28.9000 ;
	    RECT 265.0000 28.6000 265.3000 28.9000 ;
	    RECT 263.0000 28.2000 263.4000 28.6000 ;
	    RECT 263.9000 28.3000 265.3000 28.6000 ;
	    RECT 267.0000 28.5000 267.4000 28.9000 ;
	    RECT 263.9000 28.2000 264.3000 28.3000 ;
	    RECT 261.0000 27.1000 261.8000 27.2000 ;
	    RECT 263.1000 27.1000 263.4000 28.2000 ;
	    RECT 267.9000 27.7000 268.3000 27.8000 ;
	    RECT 269.4000 27.7000 269.8000 29.9000 ;
	    RECT 267.9000 27.4000 269.8000 27.7000 ;
	    RECT 265.9000 27.1000 266.3000 27.2000 ;
	    RECT 261.0000 26.8000 266.5000 27.1000 ;
	    RECT 262.5000 26.7000 262.9000 26.8000 ;
	    RECT 261.7000 26.2000 262.1000 26.3000 ;
	    RECT 261.7000 25.9000 264.2000 26.2000 ;
	    RECT 263.8000 25.8000 264.2000 25.9000 ;
	    RECT 260.6000 25.5000 263.4000 25.6000 ;
	    RECT 260.6000 25.4000 263.5000 25.5000 ;
	    RECT 260.6000 25.3000 265.5000 25.4000 ;
	    RECT 260.6000 21.1000 261.0000 25.3000 ;
	    RECT 263.1000 25.1000 265.5000 25.3000 ;
	    RECT 262.2000 24.5000 264.9000 24.8000 ;
	    RECT 262.2000 24.4000 262.6000 24.5000 ;
	    RECT 264.5000 24.4000 264.9000 24.5000 ;
	    RECT 265.2000 24.5000 265.5000 25.1000 ;
	    RECT 266.2000 25.2000 266.5000 26.8000 ;
	    RECT 267.0000 26.4000 267.4000 26.5000 ;
	    RECT 267.0000 26.1000 268.9000 26.4000 ;
	    RECT 268.5000 26.0000 268.9000 26.1000 ;
	    RECT 267.7000 25.7000 268.1000 25.8000 ;
	    RECT 269.4000 25.7000 269.8000 27.4000 ;
	    RECT 267.7000 25.4000 269.8000 25.7000 ;
	    RECT 266.2000 24.9000 267.4000 25.2000 ;
	    RECT 265.9000 24.5000 266.3000 24.6000 ;
	    RECT 265.2000 24.2000 266.3000 24.5000 ;
	    RECT 267.1000 24.4000 267.4000 24.9000 ;
	    RECT 267.1000 24.0000 267.8000 24.4000 ;
	    RECT 263.9000 23.7000 264.3000 23.8000 ;
	    RECT 265.3000 23.7000 265.7000 23.8000 ;
	    RECT 262.2000 23.1000 262.6000 23.5000 ;
	    RECT 263.9000 23.4000 265.7000 23.7000 ;
	    RECT 265.0000 23.1000 265.3000 23.4000 ;
	    RECT 267.0000 23.1000 267.4000 23.5000 ;
	    RECT 262.2000 22.8000 263.2000 23.1000 ;
	    RECT 262.8000 21.1000 263.2000 22.8000 ;
	    RECT 265.0000 21.1000 265.4000 23.1000 ;
	    RECT 267.1000 21.1000 267.7000 23.1000 ;
	    RECT 269.4000 21.1000 269.8000 25.4000 ;
	    RECT 0.6000 14.1000 1.0000 19.9000 ;
	    RECT 3.5000 16.3000 3.9000 19.9000 ;
	    RECT 3.0000 15.9000 3.9000 16.3000 ;
	    RECT 2.2000 15.1000 2.6000 15.2000 ;
	    RECT 3.1000 15.1000 3.4000 15.9000 ;
	    RECT 4.6000 15.6000 5.0000 19.9000 ;
	    RECT 6.7000 17.9000 7.3000 19.9000 ;
	    RECT 9.0000 17.9000 9.4000 19.9000 ;
	    RECT 11.2000 18.2000 11.6000 19.9000 ;
	    RECT 11.2000 17.9000 12.2000 18.2000 ;
	    RECT 7.0000 17.5000 7.4000 17.9000 ;
	    RECT 9.1000 17.6000 9.4000 17.9000 ;
	    RECT 8.7000 17.3000 10.5000 17.6000 ;
	    RECT 11.8000 17.5000 12.2000 17.9000 ;
	    RECT 8.7000 17.2000 9.1000 17.3000 ;
	    RECT 10.1000 17.2000 10.5000 17.3000 ;
	    RECT 6.6000 16.6000 7.3000 17.0000 ;
	    RECT 7.0000 16.1000 7.3000 16.6000 ;
	    RECT 8.1000 16.5000 9.2000 16.8000 ;
	    RECT 8.1000 16.4000 8.5000 16.5000 ;
	    RECT 7.0000 15.8000 8.2000 16.1000 ;
	    RECT 2.2000 14.8000 3.4000 15.1000 ;
	    RECT 3.8000 14.8000 4.2000 15.6000 ;
	    RECT 4.6000 15.3000 6.7000 15.6000 ;
	    RECT 3.1000 14.2000 3.4000 14.8000 ;
	    RECT 0.6000 13.8000 2.5000 14.1000 ;
	    RECT 3.0000 13.8000 3.4000 14.2000 ;
	    RECT 0.6000 11.1000 1.0000 13.8000 ;
	    RECT 2.2000 13.2000 2.5000 13.8000 ;
	    RECT 1.4000 12.4000 1.8000 13.2000 ;
	    RECT 2.2000 12.4000 2.6000 13.2000 ;
	    RECT 3.1000 12.1000 3.4000 13.8000 ;
	    RECT 3.0000 11.1000 3.4000 12.1000 ;
	    RECT 4.6000 13.6000 5.0000 15.3000 ;
	    RECT 6.3000 15.2000 6.7000 15.3000 ;
	    RECT 5.5000 14.9000 5.9000 15.0000 ;
	    RECT 5.5000 14.6000 7.4000 14.9000 ;
	    RECT 7.0000 14.5000 7.4000 14.6000 ;
	    RECT 7.9000 14.2000 8.2000 15.8000 ;
	    RECT 8.9000 15.9000 9.2000 16.5000 ;
	    RECT 9.5000 16.5000 9.9000 16.6000 ;
	    RECT 11.8000 16.5000 12.2000 16.6000 ;
	    RECT 9.5000 16.2000 12.2000 16.5000 ;
	    RECT 8.9000 15.7000 11.3000 15.9000 ;
	    RECT 13.4000 15.7000 13.8000 19.9000 ;
	    RECT 14.5000 16.3000 14.9000 19.9000 ;
	    RECT 14.5000 15.9000 15.4000 16.3000 ;
	    RECT 8.9000 15.6000 13.8000 15.7000 ;
	    RECT 10.9000 15.5000 13.8000 15.6000 ;
	    RECT 11.0000 15.4000 13.8000 15.5000 ;
	    RECT 10.2000 15.1000 10.6000 15.2000 ;
	    RECT 10.2000 14.8000 12.7000 15.1000 ;
	    RECT 14.2000 14.8000 14.6000 15.6000 ;
	    RECT 15.0000 15.1000 15.3000 15.9000 ;
	    RECT 15.0000 14.8000 16.1000 15.1000 ;
	    RECT 12.3000 14.7000 12.7000 14.8000 ;
	    RECT 11.5000 14.2000 11.9000 14.3000 ;
	    RECT 15.0000 14.2000 15.3000 14.8000 ;
	    RECT 15.8000 14.2000 16.1000 14.8000 ;
	    RECT 7.9000 13.9000 13.4000 14.2000 ;
	    RECT 8.1000 13.8000 8.5000 13.9000 ;
	    RECT 4.6000 13.3000 6.5000 13.6000 ;
	    RECT 4.6000 11.1000 5.0000 13.3000 ;
	    RECT 6.1000 13.2000 6.5000 13.3000 ;
	    RECT 11.0000 12.8000 11.3000 13.9000 ;
	    RECT 12.6000 13.8000 13.4000 13.9000 ;
	    RECT 15.0000 13.8000 15.4000 14.2000 ;
	    RECT 15.8000 13.8000 16.2000 14.2000 ;
	    RECT 10.1000 12.7000 10.5000 12.8000 ;
	    RECT 7.0000 12.1000 7.4000 12.5000 ;
	    RECT 9.1000 12.4000 10.5000 12.7000 ;
	    RECT 11.0000 12.4000 11.4000 12.8000 ;
	    RECT 9.1000 12.1000 9.4000 12.4000 ;
	    RECT 11.8000 12.1000 12.2000 12.5000 ;
	    RECT 6.7000 11.8000 7.4000 12.1000 ;
	    RECT 6.7000 11.1000 7.3000 11.8000 ;
	    RECT 9.0000 11.1000 9.4000 12.1000 ;
	    RECT 11.2000 11.8000 12.2000 12.1000 ;
	    RECT 11.2000 11.1000 11.6000 11.8000 ;
	    RECT 13.4000 11.1000 13.8000 13.5000 ;
	    RECT 15.0000 12.1000 15.3000 13.8000 ;
	    RECT 15.8000 13.1000 16.2000 13.2000 ;
	    RECT 16.6000 13.1000 17.0000 19.9000 ;
	    RECT 18.2000 15.6000 18.6000 19.9000 ;
	    RECT 20.3000 17.9000 20.9000 19.9000 ;
	    RECT 22.6000 17.9000 23.0000 19.9000 ;
	    RECT 24.8000 18.2000 25.2000 19.9000 ;
	    RECT 24.8000 17.9000 25.8000 18.2000 ;
	    RECT 20.6000 17.5000 21.0000 17.9000 ;
	    RECT 22.7000 17.6000 23.0000 17.9000 ;
	    RECT 22.3000 17.3000 24.1000 17.6000 ;
	    RECT 25.4000 17.5000 25.8000 17.9000 ;
	    RECT 22.3000 17.2000 22.7000 17.3000 ;
	    RECT 23.7000 17.2000 24.1000 17.3000 ;
	    RECT 20.2000 16.6000 20.9000 17.0000 ;
	    RECT 20.6000 16.1000 20.9000 16.6000 ;
	    RECT 21.7000 16.5000 22.8000 16.8000 ;
	    RECT 21.7000 16.4000 22.1000 16.5000 ;
	    RECT 20.6000 15.8000 21.8000 16.1000 ;
	    RECT 18.2000 15.3000 20.3000 15.6000 ;
	    RECT 18.2000 13.6000 18.6000 15.3000 ;
	    RECT 19.9000 15.2000 20.3000 15.3000 ;
	    RECT 19.1000 14.9000 19.5000 15.0000 ;
	    RECT 19.1000 14.6000 21.0000 14.9000 ;
	    RECT 20.6000 14.5000 21.0000 14.6000 ;
	    RECT 21.5000 14.2000 21.8000 15.8000 ;
	    RECT 22.5000 15.9000 22.8000 16.5000 ;
	    RECT 23.1000 16.5000 23.5000 16.6000 ;
	    RECT 25.4000 16.5000 25.8000 16.6000 ;
	    RECT 23.1000 16.2000 25.8000 16.5000 ;
	    RECT 22.5000 15.7000 24.9000 15.9000 ;
	    RECT 27.0000 15.7000 27.4000 19.9000 ;
	    RECT 27.8000 16.2000 28.2000 19.9000 ;
	    RECT 27.8000 15.9000 28.9000 16.2000 ;
	    RECT 29.4000 15.9000 29.8000 19.9000 ;
	    RECT 22.5000 15.6000 27.4000 15.7000 ;
	    RECT 24.5000 15.5000 27.4000 15.6000 ;
	    RECT 24.6000 15.4000 27.4000 15.5000 ;
	    RECT 28.6000 15.6000 28.9000 15.9000 ;
	    RECT 28.6000 15.2000 29.2000 15.6000 ;
	    RECT 23.8000 15.1000 24.2000 15.2000 ;
	    RECT 23.8000 14.8000 26.3000 15.1000 ;
	    RECT 25.9000 14.7000 26.3000 14.8000 ;
	    RECT 25.1000 14.2000 25.5000 14.3000 ;
	    RECT 21.5000 13.9000 27.0000 14.2000 ;
	    RECT 21.7000 13.8000 22.1000 13.9000 ;
	    RECT 18.2000 13.3000 20.2000 13.6000 ;
	    RECT 15.8000 12.8000 17.0000 13.1000 ;
	    RECT 15.8000 12.4000 16.2000 12.8000 ;
	    RECT 15.0000 11.1000 15.4000 12.1000 ;
	    RECT 16.6000 11.1000 17.0000 12.8000 ;
	    RECT 17.4000 13.1000 17.8000 13.2000 ;
	    RECT 18.2000 13.1000 18.6000 13.3000 ;
	    RECT 19.7000 13.2000 20.2000 13.3000 ;
	    RECT 17.4000 12.8000 18.6000 13.1000 ;
	    RECT 19.8000 12.8000 20.2000 13.2000 ;
	    RECT 24.6000 12.8000 24.9000 13.9000 ;
	    RECT 26.2000 13.8000 27.0000 13.9000 ;
	    RECT 28.6000 13.7000 28.9000 15.2000 ;
	    RECT 29.5000 14.8000 29.8000 15.9000 ;
	    RECT 30.2000 15.7000 30.6000 19.9000 ;
	    RECT 32.4000 18.2000 32.8000 19.9000 ;
	    RECT 31.8000 17.9000 32.8000 18.2000 ;
	    RECT 34.6000 17.9000 35.0000 19.9000 ;
	    RECT 36.7000 17.9000 37.3000 19.9000 ;
	    RECT 31.8000 17.5000 32.2000 17.9000 ;
	    RECT 34.6000 17.6000 34.9000 17.9000 ;
	    RECT 33.5000 17.3000 35.3000 17.6000 ;
	    RECT 36.6000 17.5000 37.0000 17.9000 ;
	    RECT 33.5000 17.2000 33.9000 17.3000 ;
	    RECT 34.9000 17.2000 35.3000 17.3000 ;
	    RECT 31.8000 16.5000 32.2000 16.6000 ;
	    RECT 34.1000 16.5000 34.5000 16.6000 ;
	    RECT 31.8000 16.2000 34.5000 16.5000 ;
	    RECT 34.8000 16.5000 35.9000 16.8000 ;
	    RECT 34.8000 15.9000 35.1000 16.5000 ;
	    RECT 35.5000 16.4000 35.9000 16.5000 ;
	    RECT 36.7000 16.6000 37.4000 17.0000 ;
	    RECT 36.7000 16.1000 37.0000 16.6000 ;
	    RECT 32.7000 15.7000 35.1000 15.9000 ;
	    RECT 30.2000 15.6000 35.1000 15.7000 ;
	    RECT 35.8000 15.8000 37.0000 16.1000 ;
	    RECT 30.2000 15.5000 33.1000 15.6000 ;
	    RECT 30.2000 15.4000 33.0000 15.5000 ;
	    RECT 35.8000 15.2000 36.1000 15.8000 ;
	    RECT 39.0000 15.6000 39.4000 19.9000 ;
	    RECT 40.1000 16.2000 40.5000 19.9000 ;
	    RECT 37.3000 15.3000 39.4000 15.6000 ;
	    RECT 37.3000 15.2000 37.7000 15.3000 ;
	    RECT 33.4000 15.1000 33.8000 15.2000 ;
	    RECT 17.4000 12.4000 17.8000 12.8000 ;
	    RECT 18.2000 11.1000 18.6000 12.8000 ;
	    RECT 23.7000 12.7000 24.1000 12.8000 ;
	    RECT 20.6000 12.1000 21.0000 12.5000 ;
	    RECT 22.7000 12.4000 24.1000 12.7000 ;
	    RECT 24.6000 12.4000 25.0000 12.8000 ;
	    RECT 22.7000 12.1000 23.0000 12.4000 ;
	    RECT 25.4000 12.1000 25.8000 12.5000 ;
	    RECT 20.3000 11.8000 21.0000 12.1000 ;
	    RECT 20.3000 11.1000 20.9000 11.8000 ;
	    RECT 22.6000 11.1000 23.0000 12.1000 ;
	    RECT 24.8000 11.8000 25.8000 12.1000 ;
	    RECT 24.8000 11.1000 25.2000 11.8000 ;
	    RECT 27.0000 11.1000 27.4000 13.5000 ;
	    RECT 27.8000 13.4000 28.9000 13.7000 ;
	    RECT 27.8000 11.1000 28.2000 13.4000 ;
	    RECT 29.4000 11.1000 29.8000 14.8000 ;
	    RECT 31.3000 14.8000 33.8000 15.1000 ;
	    RECT 35.8000 14.8000 36.2000 15.2000 ;
	    RECT 38.1000 14.9000 38.5000 15.0000 ;
	    RECT 31.3000 14.7000 31.7000 14.8000 ;
	    RECT 32.1000 14.2000 32.5000 14.3000 ;
	    RECT 35.8000 14.2000 36.1000 14.8000 ;
	    RECT 36.6000 14.6000 38.5000 14.9000 ;
	    RECT 36.6000 14.5000 37.0000 14.6000 ;
	    RECT 30.6000 13.9000 36.1000 14.2000 ;
	    RECT 30.6000 13.8000 31.4000 13.9000 ;
	    RECT 30.2000 11.1000 30.6000 13.5000 ;
	    RECT 32.7000 12.8000 33.0000 13.9000 ;
	    RECT 35.5000 13.8000 35.9000 13.9000 ;
	    RECT 39.0000 13.6000 39.4000 15.3000 ;
	    RECT 37.5000 13.3000 39.4000 13.6000 ;
	    RECT 37.5000 13.2000 37.9000 13.3000 ;
	    RECT 31.8000 12.1000 32.2000 12.5000 ;
	    RECT 32.6000 12.4000 33.0000 12.8000 ;
	    RECT 33.5000 12.7000 33.9000 12.8000 ;
	    RECT 33.5000 12.4000 34.9000 12.7000 ;
	    RECT 34.6000 12.1000 34.9000 12.4000 ;
	    RECT 36.6000 12.1000 37.0000 12.5000 ;
	    RECT 31.8000 11.8000 32.8000 12.1000 ;
	    RECT 32.4000 11.1000 32.8000 11.8000 ;
	    RECT 34.6000 11.1000 35.0000 12.1000 ;
	    RECT 36.6000 11.8000 37.3000 12.1000 ;
	    RECT 36.7000 11.1000 37.3000 11.8000 ;
	    RECT 39.0000 11.1000 39.4000 13.3000 ;
	    RECT 39.8000 15.9000 40.5000 16.2000 ;
	    RECT 39.8000 15.2000 40.1000 15.9000 ;
	    RECT 42.2000 15.6000 42.6000 19.9000 ;
	    RECT 43.3000 19.2000 43.7000 19.9000 ;
	    RECT 43.3000 18.8000 44.2000 19.2000 ;
	    RECT 43.3000 16.3000 43.7000 18.8000 ;
	    RECT 43.3000 15.9000 44.2000 16.3000 ;
	    RECT 40.6000 15.4000 42.6000 15.6000 ;
	    RECT 40.5000 15.3000 42.6000 15.4000 ;
	    RECT 39.8000 14.8000 40.2000 15.2000 ;
	    RECT 40.5000 15.0000 40.9000 15.3000 ;
	    RECT 39.8000 13.1000 40.1000 14.8000 ;
	    RECT 40.5000 13.5000 40.8000 15.0000 ;
	    RECT 43.0000 14.8000 43.4000 15.6000 ;
	    RECT 41.2000 14.2000 41.6000 14.6000 ;
	    RECT 43.8000 14.2000 44.1000 15.9000 ;
	    RECT 41.3000 13.8000 41.8000 14.2000 ;
	    RECT 43.8000 13.8000 44.2000 14.2000 ;
	    RECT 40.5000 13.2000 41.7000 13.5000 ;
	    RECT 39.8000 11.1000 40.2000 13.1000 ;
	    RECT 41.4000 12.1000 41.7000 13.2000 ;
	    RECT 42.2000 13.1000 42.6000 13.2000 ;
	    RECT 43.0000 13.1000 43.4000 13.2000 ;
	    RECT 42.2000 12.8000 43.4000 13.1000 ;
	    RECT 42.2000 12.4000 42.6000 12.8000 ;
	    RECT 43.8000 12.1000 44.1000 13.8000 ;
	    RECT 44.6000 13.1000 45.0000 13.2000 ;
	    RECT 45.4000 13.1000 45.8000 19.9000 ;
	    RECT 47.8000 15.1000 48.2000 19.9000 ;
	    RECT 48.9000 16.3000 49.3000 19.9000 ;
	    RECT 48.9000 15.9000 49.8000 16.3000 ;
	    RECT 51.0000 16.2000 51.4000 19.9000 ;
	    RECT 53.2000 17.2000 54.0000 19.9000 ;
	    RECT 53.2000 16.8000 54.6000 17.2000 ;
	    RECT 51.8000 16.2000 52.2000 16.3000 ;
	    RECT 53.2000 16.2000 54.0000 16.8000 ;
	    RECT 51.0000 15.9000 52.2000 16.2000 ;
	    RECT 53.0000 15.9000 54.0000 16.2000 ;
	    RECT 55.1000 16.2000 55.5000 16.3000 ;
	    RECT 55.8000 16.2000 56.2000 19.9000 ;
	    RECT 55.1000 15.9000 56.2000 16.2000 ;
	    RECT 58.2000 15.9000 58.6000 19.9000 ;
	    RECT 59.0000 16.2000 59.4000 19.9000 ;
	    RECT 60.6000 16.2000 61.0000 19.9000 ;
	    RECT 59.0000 15.9000 61.0000 16.2000 ;
	    RECT 48.6000 15.1000 49.0000 15.6000 ;
	    RECT 47.8000 14.8000 49.0000 15.1000 ;
	    RECT 44.6000 12.8000 45.8000 13.1000 ;
	    RECT 44.6000 12.4000 45.0000 12.8000 ;
	    RECT 41.4000 11.1000 41.8000 12.1000 ;
	    RECT 43.8000 11.1000 44.2000 12.1000 ;
	    RECT 45.4000 11.1000 45.8000 12.8000 ;
	    RECT 46.2000 12.4000 46.6000 13.2000 ;
	    RECT 47.0000 12.4000 47.4000 13.2000 ;
	    RECT 47.8000 11.1000 48.2000 14.8000 ;
	    RECT 49.4000 14.2000 49.7000 15.9000 ;
	    RECT 53.0000 15.2000 53.3000 15.9000 ;
	    RECT 55.1000 15.6000 55.4000 15.9000 ;
	    RECT 53.7000 15.3000 55.4000 15.6000 ;
	    RECT 53.7000 15.2000 54.1000 15.3000 ;
	    RECT 58.3000 15.2000 58.6000 15.9000 ;
	    RECT 60.2000 15.2000 60.6000 15.4000 ;
	    RECT 52.6000 14.9000 53.3000 15.2000 ;
	    RECT 54.8000 14.9000 55.2000 15.0000 ;
	    RECT 52.6000 14.8000 53.5000 14.9000 ;
	    RECT 53.0000 14.6000 53.5000 14.8000 ;
	    RECT 49.4000 13.8000 49.8000 14.2000 ;
	    RECT 50.2000 14.1000 50.6000 14.2000 ;
	    RECT 51.0000 14.1000 51.8000 14.2000 ;
	    RECT 50.2000 13.8000 51.8000 14.1000 ;
	    RECT 52.4000 13.8000 52.8000 14.2000 ;
	    RECT 48.6000 13.1000 49.0000 13.2000 ;
	    RECT 49.4000 13.1000 49.7000 13.8000 ;
	    RECT 52.5000 13.6000 52.8000 13.8000 ;
	    RECT 51.8000 13.4000 52.2000 13.5000 ;
	    RECT 48.6000 12.8000 49.7000 13.1000 ;
	    RECT 49.4000 12.1000 49.7000 12.8000 ;
	    RECT 50.2000 12.4000 50.6000 13.2000 ;
	    RECT 51.0000 13.1000 52.2000 13.4000 ;
	    RECT 52.5000 13.2000 52.9000 13.6000 ;
	    RECT 49.4000 11.1000 49.8000 12.1000 ;
	    RECT 51.0000 11.1000 51.4000 13.1000 ;
	    RECT 53.2000 12.9000 53.5000 14.6000 ;
	    RECT 53.9000 14.6000 55.2000 14.9000 ;
	    RECT 58.2000 14.9000 59.4000 15.2000 ;
	    RECT 60.2000 15.1000 61.0000 15.2000 ;
	    RECT 61.4000 15.1000 61.8000 15.2000 ;
	    RECT 60.2000 14.9000 61.8000 15.1000 ;
	    RECT 58.2000 14.8000 58.6000 14.9000 ;
	    RECT 59.0000 14.8000 59.4000 14.9000 ;
	    RECT 60.6000 14.8000 61.8000 14.9000 ;
	    RECT 53.9000 14.3000 54.2000 14.6000 ;
	    RECT 53.8000 13.9000 54.2000 14.3000 ;
	    RECT 55.4000 14.1000 56.2000 14.2000 ;
	    RECT 54.5000 13.8000 56.2000 14.1000 ;
	    RECT 54.5000 13.6000 54.8000 13.8000 ;
	    RECT 53.8000 13.3000 54.8000 13.6000 ;
	    RECT 55.1000 13.4000 55.5000 13.5000 ;
	    RECT 53.8000 13.2000 54.6000 13.3000 ;
	    RECT 55.1000 13.1000 56.2000 13.4000 ;
	    RECT 53.2000 11.1000 54.0000 12.9000 ;
	    RECT 55.8000 11.1000 56.2000 13.1000 ;
	    RECT 57.4000 13.1000 57.8000 13.2000 ;
	    RECT 58.2000 13.1000 58.6000 13.2000 ;
	    RECT 59.1000 13.1000 59.4000 14.8000 ;
	    RECT 59.8000 14.1000 60.2000 14.6000 ;
	    RECT 61.4000 14.1000 61.8000 14.2000 ;
	    RECT 59.8000 13.8000 61.8000 14.1000 ;
	    RECT 61.4000 13.4000 61.8000 13.8000 ;
	    RECT 62.2000 14.1000 62.6000 19.9000 ;
	    RECT 64.9000 19.2000 65.3000 19.9000 ;
	    RECT 64.9000 18.8000 65.8000 19.2000 ;
	    RECT 64.2000 16.8000 64.6000 17.2000 ;
	    RECT 63.0000 15.8000 63.4000 16.6000 ;
	    RECT 64.2000 16.2000 64.5000 16.8000 ;
	    RECT 64.9000 16.2000 65.3000 18.8000 ;
	    RECT 63.8000 15.9000 64.5000 16.2000 ;
	    RECT 64.8000 15.9000 65.3000 16.2000 ;
	    RECT 63.8000 15.8000 64.2000 15.9000 ;
	    RECT 63.0000 14.8000 63.4000 15.2000 ;
	    RECT 63.0000 14.1000 63.3000 14.8000 ;
	    RECT 64.8000 14.2000 65.1000 15.9000 ;
	    RECT 65.4000 14.4000 65.8000 15.2000 ;
	    RECT 67.0000 15.1000 67.4000 15.2000 ;
	    RECT 67.8000 15.1000 68.2000 19.9000 ;
	    RECT 69.9000 16.2000 70.3000 19.9000 ;
	    RECT 70.6000 16.8000 71.0000 17.2000 ;
	    RECT 70.7000 16.2000 71.0000 16.8000 ;
	    RECT 71.8000 16.2000 72.2000 19.9000 ;
	    RECT 73.4000 19.6000 75.4000 19.9000 ;
	    RECT 73.4000 16.2000 73.8000 19.6000 ;
	    RECT 69.4000 15.8000 70.4000 16.2000 ;
	    RECT 70.7000 15.9000 71.4000 16.2000 ;
	    RECT 71.8000 15.9000 73.8000 16.2000 ;
	    RECT 74.2000 15.9000 74.6000 19.3000 ;
	    RECT 75.0000 15.9000 75.4000 19.6000 ;
	    RECT 71.0000 15.8000 71.4000 15.9000 ;
	    RECT 67.0000 14.8000 68.2000 15.1000 ;
	    RECT 68.6000 15.1000 69.0000 15.2000 ;
	    RECT 69.4000 15.1000 69.8000 15.2000 ;
	    RECT 68.6000 14.8000 69.8000 15.1000 ;
	    RECT 62.2000 13.8000 63.3000 14.1000 ;
	    RECT 63.8000 13.8000 65.1000 14.2000 ;
	    RECT 66.2000 14.1000 66.6000 14.2000 ;
	    RECT 65.8000 13.8000 66.6000 14.1000 ;
	    RECT 67.8000 14.1000 68.2000 14.8000 ;
	    RECT 69.4000 14.4000 69.8000 14.8000 ;
	    RECT 70.1000 14.2000 70.4000 15.8000 ;
	    RECT 74.2000 15.6000 74.5000 15.9000 ;
	    RECT 72.2000 15.2000 72.6000 15.4000 ;
	    RECT 73.5000 15.3000 74.5000 15.6000 ;
	    RECT 73.5000 15.2000 73.8000 15.3000 ;
	    RECT 71.0000 15.1000 71.4000 15.2000 ;
	    RECT 71.8000 15.1000 72.6000 15.2000 ;
	    RECT 71.0000 14.9000 72.6000 15.1000 ;
	    RECT 71.0000 14.8000 72.2000 14.9000 ;
	    RECT 73.4000 14.8000 73.8000 15.2000 ;
	    RECT 75.0000 14.8000 75.4000 15.6000 ;
	    RECT 68.6000 14.1000 69.0000 14.2000 ;
	    RECT 67.8000 13.8000 69.4000 14.1000 ;
	    RECT 70.1000 13.8000 71.4000 14.2000 ;
	    RECT 72.6000 13.8000 73.0000 14.6000 ;
	    RECT 57.4000 12.8000 58.6000 13.1000 ;
	    RECT 58.3000 12.4000 58.7000 12.8000 ;
	    RECT 59.0000 11.1000 59.4000 13.1000 ;
	    RECT 62.2000 13.1000 62.6000 13.8000 ;
	    RECT 63.9000 13.1000 64.2000 13.8000 ;
	    RECT 65.8000 13.6000 66.2000 13.8000 ;
	    RECT 64.7000 13.1000 66.5000 13.3000 ;
	    RECT 62.2000 12.8000 63.1000 13.1000 ;
	    RECT 62.7000 11.1000 63.1000 12.8000 ;
	    RECT 63.8000 11.1000 64.2000 13.1000 ;
	    RECT 64.6000 13.0000 66.6000 13.1000 ;
	    RECT 64.6000 11.1000 65.0000 13.0000 ;
	    RECT 66.2000 11.1000 66.6000 13.0000 ;
	    RECT 67.0000 12.4000 67.4000 13.2000 ;
	    RECT 67.8000 11.1000 68.2000 13.8000 ;
	    RECT 69.0000 13.6000 69.4000 13.8000 ;
	    RECT 68.7000 13.1000 70.5000 13.3000 ;
	    RECT 71.0000 13.1000 71.3000 13.8000 ;
	    RECT 73.5000 13.1000 73.8000 14.8000 ;
	    RECT 74.1000 14.4000 74.5000 14.8000 ;
	    RECT 74.2000 14.2000 74.5000 14.4000 ;
	    RECT 74.2000 14.1000 74.6000 14.2000 ;
	    RECT 75.8000 14.1000 76.2000 19.9000 ;
	    RECT 78.2000 15.6000 78.6000 19.9000 ;
	    RECT 79.8000 15.6000 80.2000 19.9000 ;
	    RECT 81.4000 15.6000 81.8000 19.9000 ;
	    RECT 83.0000 15.6000 83.4000 19.9000 ;
	    RECT 84.9000 19.2000 85.3000 19.9000 ;
	    RECT 84.9000 18.8000 85.8000 19.2000 ;
	    RECT 84.9000 16.3000 85.3000 18.8000 ;
	    RECT 84.9000 15.9000 85.8000 16.3000 ;
	    RECT 87.0000 16.2000 87.4000 19.9000 ;
	    RECT 88.6000 16.2000 89.0000 19.9000 ;
	    RECT 87.0000 15.9000 89.0000 16.2000 ;
	    RECT 89.4000 15.9000 89.8000 19.9000 ;
	    RECT 91.3000 19.2000 91.7000 19.9000 ;
	    RECT 93.7000 19.2000 94.1000 19.9000 ;
	    RECT 91.3000 18.8000 92.2000 19.2000 ;
	    RECT 93.7000 18.8000 94.6000 19.2000 ;
	    RECT 90.6000 16.8000 91.0000 17.2000 ;
	    RECT 90.6000 16.2000 90.9000 16.8000 ;
	    RECT 91.3000 16.2000 91.7000 18.8000 ;
	    RECT 90.2000 15.9000 90.9000 16.2000 ;
	    RECT 91.2000 15.9000 91.7000 16.2000 ;
	    RECT 93.7000 16.3000 94.1000 18.8000 ;
	    RECT 96.2000 16.8000 96.6000 17.2000 ;
	    RECT 93.7000 15.9000 94.6000 16.3000 ;
	    RECT 96.2000 16.2000 96.5000 16.8000 ;
	    RECT 96.9000 16.2000 97.3000 19.9000 ;
	    RECT 95.8000 15.9000 96.5000 16.2000 ;
	    RECT 96.8000 15.9000 97.3000 16.2000 ;
	    RECT 74.2000 13.8000 76.2000 14.1000 ;
	    RECT 68.6000 13.0000 70.6000 13.1000 ;
	    RECT 68.6000 11.1000 69.0000 13.0000 ;
	    RECT 70.2000 11.1000 70.6000 13.0000 ;
	    RECT 71.0000 11.1000 71.4000 13.1000 ;
	    RECT 73.3000 12.2000 74.1000 13.1000 ;
	    RECT 73.3000 11.8000 74.6000 12.2000 ;
	    RECT 73.3000 11.1000 74.1000 11.8000 ;
	    RECT 75.8000 11.1000 76.2000 13.8000 ;
	    RECT 77.4000 15.2000 78.6000 15.6000 ;
	    RECT 79.1000 15.2000 80.2000 15.6000 ;
	    RECT 80.7000 15.2000 81.8000 15.6000 ;
	    RECT 82.5000 15.2000 83.4000 15.6000 ;
	    RECT 77.4000 13.8000 77.8000 15.2000 ;
	    RECT 79.1000 14.5000 79.5000 15.2000 ;
	    RECT 80.7000 14.5000 81.1000 15.2000 ;
	    RECT 82.5000 14.5000 82.9000 15.2000 ;
	    RECT 84.6000 14.8000 85.0000 15.6000 ;
	    RECT 78.2000 14.1000 79.5000 14.5000 ;
	    RECT 79.9000 14.1000 81.1000 14.5000 ;
	    RECT 81.6000 14.1000 82.9000 14.5000 ;
	    RECT 79.1000 13.8000 79.5000 14.1000 ;
	    RECT 80.7000 13.8000 81.1000 14.1000 ;
	    RECT 82.5000 13.8000 82.9000 14.1000 ;
	    RECT 85.4000 14.2000 85.7000 15.9000 ;
	    RECT 87.4000 15.2000 87.8000 15.4000 ;
	    RECT 89.4000 15.2000 89.7000 15.9000 ;
	    RECT 90.2000 15.8000 90.6000 15.9000 ;
	    RECT 87.0000 14.9000 87.8000 15.2000 ;
	    RECT 88.6000 14.9000 89.8000 15.2000 ;
	    RECT 87.0000 14.8000 87.4000 14.9000 ;
	    RECT 85.4000 13.8000 85.8000 14.2000 ;
	    RECT 87.8000 13.8000 88.2000 14.6000 ;
	    RECT 77.4000 13.4000 78.6000 13.8000 ;
	    RECT 79.1000 13.4000 80.2000 13.8000 ;
	    RECT 80.7000 13.4000 81.8000 13.8000 ;
	    RECT 82.5000 13.4000 83.4000 13.8000 ;
	    RECT 76.6000 12.4000 77.0000 13.2000 ;
	    RECT 78.2000 11.1000 78.6000 13.4000 ;
	    RECT 79.8000 11.1000 80.2000 13.4000 ;
	    RECT 81.4000 11.1000 81.8000 13.4000 ;
	    RECT 83.0000 11.1000 83.4000 13.4000 ;
	    RECT 85.4000 12.1000 85.7000 13.8000 ;
	    RECT 86.2000 12.4000 86.6000 13.2000 ;
	    RECT 88.6000 13.1000 88.9000 14.9000 ;
	    RECT 89.4000 14.8000 89.8000 14.9000 ;
	    RECT 91.2000 14.2000 91.5000 15.9000 ;
	    RECT 91.8000 14.4000 92.2000 15.2000 ;
	    RECT 93.4000 14.8000 93.8000 15.6000 ;
	    RECT 90.2000 13.8000 91.5000 14.2000 ;
	    RECT 92.6000 14.1000 93.0000 14.2000 ;
	    RECT 93.4000 14.1000 93.7000 14.8000 ;
	    RECT 92.2000 13.8000 93.7000 14.1000 ;
	    RECT 94.2000 14.2000 94.5000 15.9000 ;
	    RECT 95.8000 15.8000 96.2000 15.9000 ;
	    RECT 96.8000 15.1000 97.1000 15.9000 ;
	    RECT 95.0000 14.8000 97.1000 15.1000 ;
	    RECT 95.0000 14.2000 95.3000 14.8000 ;
	    RECT 96.8000 14.2000 97.1000 14.8000 ;
	    RECT 97.4000 15.1000 97.8000 15.2000 ;
	    RECT 99.0000 15.1000 99.4000 19.9000 ;
	    RECT 97.4000 14.8000 99.4000 15.1000 ;
	    RECT 97.4000 14.4000 97.8000 14.8000 ;
	    RECT 94.2000 13.8000 94.6000 14.2000 ;
	    RECT 95.0000 13.8000 95.4000 14.2000 ;
	    RECT 95.8000 13.8000 97.1000 14.2000 ;
	    RECT 98.2000 14.1000 98.6000 14.2000 ;
	    RECT 97.8000 13.8000 98.6000 14.1000 ;
	    RECT 85.4000 11.1000 85.8000 12.1000 ;
	    RECT 88.6000 11.1000 89.0000 13.1000 ;
	    RECT 89.4000 12.8000 89.8000 13.2000 ;
	    RECT 90.3000 13.1000 90.6000 13.8000 ;
	    RECT 92.2000 13.6000 92.6000 13.8000 ;
	    RECT 91.1000 13.1000 92.9000 13.3000 ;
	    RECT 89.3000 12.4000 89.7000 12.8000 ;
	    RECT 90.2000 11.1000 90.6000 13.1000 ;
	    RECT 91.0000 13.0000 93.0000 13.1000 ;
	    RECT 91.0000 11.1000 91.4000 13.0000 ;
	    RECT 92.6000 11.1000 93.0000 13.0000 ;
	    RECT 94.2000 12.1000 94.5000 13.8000 ;
	    RECT 95.0000 12.4000 95.4000 13.2000 ;
	    RECT 95.9000 13.1000 96.2000 13.8000 ;
	    RECT 97.8000 13.6000 98.2000 13.8000 ;
	    RECT 96.7000 13.1000 98.5000 13.3000 ;
	    RECT 94.2000 11.1000 94.6000 12.1000 ;
	    RECT 95.8000 11.1000 96.2000 13.1000 ;
	    RECT 96.6000 13.0000 98.6000 13.1000 ;
	    RECT 96.6000 11.1000 97.0000 13.0000 ;
	    RECT 98.2000 11.1000 98.6000 13.0000 ;
	    RECT 99.0000 11.1000 99.4000 14.8000 ;
	    RECT 101.4000 15.1000 101.8000 19.9000 ;
	    RECT 102.2000 16.2000 102.6000 19.9000 ;
	    RECT 103.8000 16.2000 104.2000 19.9000 ;
	    RECT 102.2000 15.9000 104.2000 16.2000 ;
	    RECT 104.6000 16.1000 105.0000 19.9000 ;
	    RECT 105.4000 16.1000 105.8000 16.6000 ;
	    RECT 104.6000 15.8000 105.8000 16.1000 ;
	    RECT 102.6000 15.2000 103.0000 15.4000 ;
	    RECT 104.6000 15.2000 104.9000 15.8000 ;
	    RECT 102.2000 15.1000 103.0000 15.2000 ;
	    RECT 101.4000 14.9000 103.0000 15.1000 ;
	    RECT 103.8000 14.9000 105.0000 15.2000 ;
	    RECT 101.4000 14.8000 102.6000 14.9000 ;
	    RECT 99.8000 12.4000 100.2000 13.2000 ;
	    RECT 100.6000 12.4000 101.0000 13.2000 ;
	    RECT 101.4000 11.1000 101.8000 14.8000 ;
	    RECT 103.0000 13.8000 103.4000 14.6000 ;
	    RECT 103.8000 13.1000 104.1000 14.9000 ;
	    RECT 104.6000 14.8000 105.0000 14.9000 ;
	    RECT 105.4000 13.8000 105.8000 14.2000 ;
	    RECT 105.4000 13.2000 105.7000 13.8000 ;
	    RECT 106.2000 13.2000 106.6000 19.9000 ;
	    RECT 109.8000 16.8000 110.2000 17.2000 ;
	    RECT 109.8000 16.2000 110.1000 16.8000 ;
	    RECT 110.5000 16.2000 110.9000 19.9000 ;
	    RECT 113.9000 16.3000 114.3000 19.9000 ;
	    RECT 109.4000 15.9000 110.1000 16.2000 ;
	    RECT 110.4000 15.9000 110.9000 16.2000 ;
	    RECT 113.4000 15.9000 114.3000 16.3000 ;
	    RECT 109.4000 15.8000 109.8000 15.9000 ;
	    RECT 110.4000 15.1000 110.7000 15.9000 ;
	    RECT 107.0000 14.8000 110.7000 15.1000 ;
	    RECT 107.0000 14.2000 107.3000 14.8000 ;
	    RECT 110.4000 14.2000 110.7000 14.8000 ;
	    RECT 111.0000 15.1000 111.4000 15.2000 ;
	    RECT 113.5000 15.1000 113.8000 15.9000 ;
	    RECT 111.0000 14.8000 113.8000 15.1000 ;
	    RECT 114.2000 15.1000 114.6000 15.6000 ;
	    RECT 115.0000 15.1000 115.4000 19.9000 ;
	    RECT 117.9000 16.3000 118.3000 19.9000 ;
	    RECT 117.4000 15.9000 118.3000 16.3000 ;
	    RECT 119.8000 16.1000 120.2000 19.9000 ;
	    RECT 120.6000 16.1000 121.0000 16.6000 ;
	    RECT 114.2000 14.8000 115.4000 15.1000 ;
	    RECT 116.6000 15.1000 117.0000 15.2000 ;
	    RECT 117.5000 15.1000 117.8000 15.9000 ;
	    RECT 119.8000 15.8000 121.0000 16.1000 ;
	    RECT 116.6000 14.8000 117.8000 15.1000 ;
	    RECT 118.2000 14.8000 118.6000 15.6000 ;
	    RECT 111.0000 14.4000 111.4000 14.8000 ;
	    RECT 113.5000 14.2000 113.8000 14.8000 ;
	    RECT 107.0000 13.4000 107.4000 14.2000 ;
	    RECT 109.4000 13.8000 110.7000 14.2000 ;
	    RECT 111.8000 14.1000 112.2000 14.2000 ;
	    RECT 111.4000 13.8000 112.2000 14.1000 ;
	    RECT 113.4000 13.8000 113.8000 14.2000 ;
	    RECT 103.8000 11.1000 104.2000 13.1000 ;
	    RECT 104.6000 12.8000 105.0000 13.2000 ;
	    RECT 105.4000 12.8000 106.6000 13.2000 ;
	    RECT 109.5000 13.1000 109.8000 13.8000 ;
	    RECT 111.4000 13.6000 111.8000 13.8000 ;
	    RECT 110.3000 13.1000 112.1000 13.3000 ;
	    RECT 104.5000 12.4000 104.9000 12.8000 ;
	    RECT 105.7000 11.1000 106.1000 12.8000 ;
	    RECT 109.4000 11.1000 109.8000 13.1000 ;
	    RECT 110.2000 13.0000 112.2000 13.1000 ;
	    RECT 110.2000 11.1000 110.6000 13.0000 ;
	    RECT 111.8000 11.1000 112.2000 13.0000 ;
	    RECT 112.6000 12.4000 113.0000 13.2000 ;
	    RECT 113.5000 12.1000 113.8000 13.8000 ;
	    RECT 113.4000 11.1000 113.8000 12.1000 ;
	    RECT 115.0000 11.1000 115.4000 14.8000 ;
	    RECT 117.5000 14.2000 117.8000 14.8000 ;
	    RECT 117.4000 13.8000 117.8000 14.2000 ;
	    RECT 115.8000 12.4000 116.2000 13.2000 ;
	    RECT 116.6000 12.4000 117.0000 13.2000 ;
	    RECT 117.5000 12.1000 117.8000 13.8000 ;
	    RECT 119.0000 12.4000 119.4000 13.2000 ;
	    RECT 117.4000 11.1000 117.8000 12.1000 ;
	    RECT 119.8000 11.1000 120.2000 15.8000 ;
	    RECT 121.4000 13.1000 121.8000 19.9000 ;
	    RECT 122.2000 15.8000 122.6000 16.2000 ;
	    RECT 122.2000 15.1000 122.5000 15.8000 ;
	    RECT 123.0000 15.1000 123.4000 19.9000 ;
	    RECT 122.2000 14.8000 123.4000 15.1000 ;
	    RECT 122.2000 13.4000 122.6000 14.2000 ;
	    RECT 120.9000 12.8000 121.8000 13.1000 ;
	    RECT 120.9000 12.2000 121.3000 12.8000 ;
	    RECT 120.9000 11.8000 121.8000 12.2000 ;
	    RECT 120.9000 11.1000 121.3000 11.8000 ;
	    RECT 123.0000 11.1000 123.4000 14.8000 ;
	    RECT 124.6000 15.6000 125.0000 19.9000 ;
	    RECT 126.7000 17.9000 127.3000 19.9000 ;
	    RECT 129.0000 17.9000 129.4000 19.9000 ;
	    RECT 131.2000 18.2000 131.6000 19.9000 ;
	    RECT 131.2000 17.9000 132.2000 18.2000 ;
	    RECT 127.0000 17.5000 127.4000 17.9000 ;
	    RECT 129.1000 17.6000 129.4000 17.9000 ;
	    RECT 128.7000 17.3000 130.5000 17.6000 ;
	    RECT 131.8000 17.5000 132.2000 17.9000 ;
	    RECT 128.7000 17.2000 129.1000 17.3000 ;
	    RECT 130.1000 17.2000 130.5000 17.3000 ;
	    RECT 126.6000 16.6000 127.3000 17.0000 ;
	    RECT 127.0000 16.1000 127.3000 16.6000 ;
	    RECT 128.1000 16.5000 129.2000 16.8000 ;
	    RECT 128.1000 16.4000 128.5000 16.5000 ;
	    RECT 127.0000 15.8000 128.2000 16.1000 ;
	    RECT 124.6000 15.3000 126.7000 15.6000 ;
	    RECT 124.6000 13.6000 125.0000 15.3000 ;
	    RECT 126.3000 15.2000 126.7000 15.3000 ;
	    RECT 125.5000 14.9000 125.9000 15.0000 ;
	    RECT 125.5000 14.6000 127.4000 14.9000 ;
	    RECT 127.0000 14.5000 127.4000 14.6000 ;
	    RECT 127.9000 14.2000 128.2000 15.8000 ;
	    RECT 128.9000 15.9000 129.2000 16.5000 ;
	    RECT 129.5000 16.5000 129.9000 16.6000 ;
	    RECT 131.8000 16.5000 132.2000 16.6000 ;
	    RECT 129.5000 16.2000 132.2000 16.5000 ;
	    RECT 128.9000 15.7000 131.3000 15.9000 ;
	    RECT 133.4000 15.7000 133.8000 19.9000 ;
	    RECT 128.9000 15.6000 133.8000 15.7000 ;
	    RECT 130.9000 15.5000 133.8000 15.6000 ;
	    RECT 131.0000 15.4000 133.8000 15.5000 ;
	    RECT 130.2000 15.1000 130.6000 15.2000 ;
	    RECT 130.2000 14.8000 132.7000 15.1000 ;
	    RECT 131.0000 14.7000 131.4000 14.8000 ;
	    RECT 132.3000 14.7000 132.7000 14.8000 ;
	    RECT 131.5000 14.2000 131.9000 14.3000 ;
	    RECT 127.9000 13.9000 133.4000 14.2000 ;
	    RECT 128.1000 13.8000 128.5000 13.9000 ;
	    RECT 130.2000 13.8000 130.6000 13.9000 ;
	    RECT 124.6000 13.3000 126.5000 13.6000 ;
	    RECT 123.8000 12.4000 124.2000 13.2000 ;
	    RECT 124.6000 11.1000 125.0000 13.3000 ;
	    RECT 126.1000 13.2000 126.5000 13.3000 ;
	    RECT 131.0000 12.8000 131.3000 13.9000 ;
	    RECT 132.6000 13.8000 133.4000 13.9000 ;
	    RECT 130.1000 12.7000 130.5000 12.8000 ;
	    RECT 127.0000 12.1000 127.4000 12.5000 ;
	    RECT 129.1000 12.4000 130.5000 12.7000 ;
	    RECT 131.0000 12.4000 131.4000 12.8000 ;
	    RECT 129.1000 12.1000 129.4000 12.4000 ;
	    RECT 131.8000 12.1000 132.2000 12.5000 ;
	    RECT 126.7000 11.8000 127.4000 12.1000 ;
	    RECT 126.7000 11.1000 127.3000 11.8000 ;
	    RECT 129.0000 11.1000 129.4000 12.1000 ;
	    RECT 131.2000 11.8000 132.2000 12.1000 ;
	    RECT 131.2000 11.1000 131.6000 11.8000 ;
	    RECT 133.4000 11.1000 133.8000 13.5000 ;
	    RECT 134.2000 12.4000 134.6000 13.2000 ;
	    RECT 135.0000 13.1000 135.4000 19.9000 ;
	    RECT 137.1000 16.3000 137.5000 19.9000 ;
	    RECT 136.6000 15.9000 137.5000 16.3000 ;
	    RECT 138.2000 16.2000 138.6000 19.9000 ;
	    RECT 139.0000 16.2000 139.4000 16.3000 ;
	    RECT 140.4000 16.2000 141.2000 19.9000 ;
	    RECT 138.2000 15.9000 139.4000 16.2000 ;
	    RECT 140.2000 15.9000 141.2000 16.2000 ;
	    RECT 142.3000 16.2000 142.7000 16.3000 ;
	    RECT 143.0000 16.2000 143.4000 19.9000 ;
	    RECT 142.3000 15.9000 143.4000 16.2000 ;
	    RECT 136.6000 15.8000 137.0000 15.9000 ;
	    RECT 136.7000 14.2000 137.0000 15.8000 ;
	    RECT 137.4000 14.8000 137.8000 15.6000 ;
	    RECT 140.2000 15.2000 140.5000 15.9000 ;
	    RECT 142.3000 15.6000 142.6000 15.9000 ;
	    RECT 140.9000 15.3000 142.6000 15.6000 ;
	    RECT 140.9000 15.2000 141.3000 15.3000 ;
	    RECT 139.8000 14.9000 140.5000 15.2000 ;
	    RECT 142.0000 14.9000 142.4000 15.0000 ;
	    RECT 139.8000 14.8000 140.7000 14.9000 ;
	    RECT 140.2000 14.6000 140.7000 14.8000 ;
	    RECT 136.6000 13.8000 137.0000 14.2000 ;
	    RECT 138.2000 13.8000 139.0000 14.2000 ;
	    RECT 139.6000 13.8000 140.0000 14.2000 ;
	    RECT 135.8000 13.1000 136.2000 13.2000 ;
	    RECT 135.0000 12.8000 136.2000 13.1000 ;
	    RECT 135.0000 11.1000 135.4000 12.8000 ;
	    RECT 135.8000 12.4000 136.2000 12.8000 ;
	    RECT 136.7000 12.1000 137.0000 13.8000 ;
	    RECT 139.7000 13.6000 140.0000 13.8000 ;
	    RECT 139.0000 13.4000 139.4000 13.5000 ;
	    RECT 136.6000 11.1000 137.0000 12.1000 ;
	    RECT 138.2000 13.1000 139.4000 13.4000 ;
	    RECT 139.7000 13.2000 140.1000 13.6000 ;
	    RECT 138.2000 11.1000 138.6000 13.1000 ;
	    RECT 140.4000 12.9000 140.7000 14.6000 ;
	    RECT 141.1000 14.6000 142.4000 14.9000 ;
	    RECT 141.1000 14.3000 141.4000 14.6000 ;
	    RECT 141.0000 13.9000 141.4000 14.3000 ;
	    RECT 142.6000 14.1000 143.4000 14.2000 ;
	    RECT 141.7000 13.8000 143.4000 14.1000 ;
	    RECT 141.7000 13.6000 142.0000 13.8000 ;
	    RECT 141.0000 13.3000 142.0000 13.6000 ;
	    RECT 142.3000 13.4000 142.7000 13.5000 ;
	    RECT 141.0000 13.2000 141.8000 13.3000 ;
	    RECT 142.3000 13.1000 143.4000 13.4000 ;
	    RECT 140.4000 11.1000 141.2000 12.9000 ;
	    RECT 143.0000 11.1000 143.4000 13.1000 ;
	    RECT 143.8000 12.4000 144.2000 13.2000 ;
	    RECT 144.6000 13.1000 145.0000 19.9000 ;
	    RECT 146.7000 16.3000 147.1000 19.9000 ;
	    RECT 146.2000 15.9000 147.1000 16.3000 ;
	    RECT 146.3000 14.2000 146.6000 15.9000 ;
	    RECT 148.6000 15.6000 149.0000 19.9000 ;
	    RECT 150.2000 15.6000 150.6000 19.9000 ;
	    RECT 151.8000 15.6000 152.2000 19.9000 ;
	    RECT 153.4000 15.6000 153.8000 19.9000 ;
	    RECT 155.8000 16.4000 156.2000 19.9000 ;
	    RECT 155.7000 15.9000 156.2000 16.4000 ;
	    RECT 157.4000 16.2000 157.8000 19.9000 ;
	    RECT 156.5000 15.9000 157.8000 16.2000 ;
	    RECT 147.0000 14.8000 147.4000 15.6000 ;
	    RECT 148.6000 15.2000 149.5000 15.6000 ;
	    RECT 150.2000 15.2000 151.3000 15.6000 ;
	    RECT 151.8000 15.2000 152.9000 15.6000 ;
	    RECT 153.4000 15.2000 154.6000 15.6000 ;
	    RECT 146.2000 13.8000 146.6000 14.2000 ;
	    RECT 149.1000 14.5000 149.5000 15.2000 ;
	    RECT 150.9000 14.5000 151.3000 15.2000 ;
	    RECT 152.5000 14.5000 152.9000 15.2000 ;
	    RECT 149.1000 14.1000 150.4000 14.5000 ;
	    RECT 150.9000 14.1000 152.1000 14.5000 ;
	    RECT 152.5000 14.1000 153.8000 14.5000 ;
	    RECT 149.1000 13.8000 149.5000 14.1000 ;
	    RECT 150.9000 13.8000 151.3000 14.1000 ;
	    RECT 152.5000 13.8000 152.9000 14.1000 ;
	    RECT 154.2000 13.8000 154.6000 15.2000 ;
	    RECT 155.7000 14.2000 156.0000 15.9000 ;
	    RECT 156.5000 14.9000 156.8000 15.9000 ;
	    RECT 156.3000 14.5000 156.8000 14.9000 ;
	    RECT 155.0000 14.1000 155.4000 14.2000 ;
	    RECT 155.7000 14.1000 156.2000 14.2000 ;
	    RECT 155.0000 13.8000 156.2000 14.1000 ;
	    RECT 145.4000 13.1000 145.8000 13.2000 ;
	    RECT 146.3000 13.1000 146.6000 13.8000 ;
	    RECT 148.6000 13.4000 149.5000 13.8000 ;
	    RECT 150.2000 13.4000 151.3000 13.8000 ;
	    RECT 151.8000 13.4000 152.9000 13.8000 ;
	    RECT 153.4000 13.4000 154.6000 13.8000 ;
	    RECT 147.0000 13.1000 147.4000 13.2000 ;
	    RECT 144.6000 12.8000 145.8000 13.1000 ;
	    RECT 146.2000 12.8000 147.4000 13.1000 ;
	    RECT 144.6000 11.1000 145.0000 12.8000 ;
	    RECT 145.4000 12.4000 145.8000 12.8000 ;
	    RECT 146.3000 12.1000 146.6000 12.8000 ;
	    RECT 146.2000 11.1000 146.6000 12.1000 ;
	    RECT 148.6000 11.1000 149.0000 13.4000 ;
	    RECT 150.2000 11.1000 150.6000 13.4000 ;
	    RECT 151.8000 11.1000 152.2000 13.4000 ;
	    RECT 153.4000 11.1000 153.8000 13.4000 ;
	    RECT 155.7000 13.1000 156.0000 13.8000 ;
	    RECT 156.5000 13.7000 156.8000 14.5000 ;
	    RECT 157.3000 14.8000 157.8000 15.2000 ;
	    RECT 157.3000 14.4000 157.7000 14.8000 ;
	    RECT 156.5000 13.4000 157.8000 13.7000 ;
	    RECT 155.7000 12.8000 156.2000 13.1000 ;
	    RECT 155.8000 11.1000 156.2000 12.8000 ;
	    RECT 157.4000 11.1000 157.8000 13.4000 ;
	    RECT 158.2000 12.4000 158.6000 13.2000 ;
	    RECT 159.0000 13.1000 159.4000 19.9000 ;
	    RECT 162.7000 16.3000 163.1000 19.9000 ;
	    RECT 162.2000 15.9000 163.1000 16.3000 ;
	    RECT 162.3000 14.2000 162.6000 15.9000 ;
	    RECT 164.6000 15.6000 165.0000 19.9000 ;
	    RECT 166.2000 15.6000 166.6000 19.9000 ;
	    RECT 167.8000 15.6000 168.2000 19.9000 ;
	    RECT 169.4000 15.6000 169.8000 19.9000 ;
	    RECT 172.6000 16.2000 173.0000 19.9000 ;
	    RECT 171.9000 15.9000 173.0000 16.2000 ;
	    RECT 171.9000 15.6000 172.2000 15.9000 ;
	    RECT 163.0000 14.8000 163.4000 15.6000 ;
	    RECT 164.6000 15.2000 165.5000 15.6000 ;
	    RECT 166.2000 15.2000 167.3000 15.6000 ;
	    RECT 167.8000 15.2000 168.9000 15.6000 ;
	    RECT 169.4000 15.2000 170.6000 15.6000 ;
	    RECT 171.6000 15.2000 172.2000 15.6000 ;
	    RECT 173.4000 15.6000 173.8000 19.9000 ;
	    RECT 175.5000 17.9000 176.1000 19.9000 ;
	    RECT 177.8000 17.9000 178.2000 19.9000 ;
	    RECT 180.0000 18.2000 180.4000 19.9000 ;
	    RECT 180.0000 17.9000 181.0000 18.2000 ;
	    RECT 175.8000 17.5000 176.2000 17.9000 ;
	    RECT 177.9000 17.6000 178.2000 17.9000 ;
	    RECT 177.5000 17.3000 179.3000 17.6000 ;
	    RECT 180.6000 17.5000 181.0000 17.9000 ;
	    RECT 177.5000 17.2000 177.9000 17.3000 ;
	    RECT 178.9000 17.2000 179.3000 17.3000 ;
	    RECT 175.4000 16.6000 176.1000 17.0000 ;
	    RECT 175.8000 16.1000 176.1000 16.6000 ;
	    RECT 176.9000 16.5000 178.0000 16.8000 ;
	    RECT 176.9000 16.4000 177.3000 16.5000 ;
	    RECT 175.8000 15.8000 177.0000 16.1000 ;
	    RECT 173.4000 15.3000 175.5000 15.6000 ;
	    RECT 162.2000 13.8000 162.6000 14.2000 ;
	    RECT 165.1000 14.5000 165.5000 15.2000 ;
	    RECT 166.9000 14.5000 167.3000 15.2000 ;
	    RECT 168.5000 14.5000 168.9000 15.2000 ;
	    RECT 165.1000 14.1000 166.4000 14.5000 ;
	    RECT 166.9000 14.1000 168.1000 14.5000 ;
	    RECT 168.5000 14.1000 169.8000 14.5000 ;
	    RECT 165.1000 13.8000 165.5000 14.1000 ;
	    RECT 166.9000 13.8000 167.3000 14.1000 ;
	    RECT 168.5000 13.8000 168.9000 14.1000 ;
	    RECT 170.2000 13.8000 170.6000 15.2000 ;
	    RECT 161.4000 13.1000 161.8000 13.2000 ;
	    RECT 162.3000 13.1000 162.6000 13.8000 ;
	    RECT 164.6000 13.4000 165.5000 13.8000 ;
	    RECT 166.2000 13.4000 167.3000 13.8000 ;
	    RECT 167.8000 13.4000 168.9000 13.8000 ;
	    RECT 169.4000 13.4000 170.6000 13.8000 ;
	    RECT 171.9000 13.7000 172.2000 15.2000 ;
	    RECT 172.6000 14.4000 173.0000 15.2000 ;
	    RECT 171.9000 13.4000 173.0000 13.7000 ;
	    RECT 163.0000 13.1000 163.4000 13.2000 ;
	    RECT 159.0000 12.8000 161.8000 13.1000 ;
	    RECT 162.2000 12.8000 163.4000 13.1000 ;
	    RECT 159.0000 11.1000 159.4000 12.8000 ;
	    RECT 161.4000 12.4000 161.8000 12.8000 ;
	    RECT 162.3000 12.1000 162.6000 12.8000 ;
	    RECT 162.2000 11.1000 162.6000 12.1000 ;
	    RECT 164.6000 11.1000 165.0000 13.4000 ;
	    RECT 166.2000 11.1000 166.6000 13.4000 ;
	    RECT 167.8000 11.1000 168.2000 13.4000 ;
	    RECT 169.4000 11.1000 169.8000 13.4000 ;
	    RECT 172.6000 11.1000 173.0000 13.4000 ;
	    RECT 173.4000 13.6000 173.8000 15.3000 ;
	    RECT 175.1000 15.2000 175.5000 15.3000 ;
	    RECT 176.7000 15.2000 177.0000 15.8000 ;
	    RECT 177.7000 15.9000 178.0000 16.5000 ;
	    RECT 178.3000 16.5000 178.7000 16.6000 ;
	    RECT 180.6000 16.5000 181.0000 16.6000 ;
	    RECT 178.3000 16.2000 181.0000 16.5000 ;
	    RECT 177.7000 15.7000 180.1000 15.9000 ;
	    RECT 182.2000 15.7000 182.6000 19.9000 ;
	    RECT 177.7000 15.6000 182.6000 15.7000 ;
	    RECT 179.7000 15.5000 182.6000 15.6000 ;
	    RECT 179.8000 15.4000 182.6000 15.5000 ;
	    RECT 174.3000 14.9000 174.7000 15.0000 ;
	    RECT 174.3000 14.6000 176.2000 14.9000 ;
	    RECT 176.6000 14.8000 177.0000 15.2000 ;
	    RECT 179.0000 15.1000 179.4000 15.2000 ;
	    RECT 179.0000 14.8000 181.5000 15.1000 ;
	    RECT 175.8000 14.5000 176.2000 14.6000 ;
	    RECT 176.7000 14.2000 177.0000 14.8000 ;
	    RECT 179.8000 14.7000 180.2000 14.8000 ;
	    RECT 181.1000 14.7000 181.5000 14.8000 ;
	    RECT 180.3000 14.2000 180.7000 14.3000 ;
	    RECT 176.7000 13.9000 182.2000 14.2000 ;
	    RECT 176.9000 13.8000 177.3000 13.9000 ;
	    RECT 173.4000 13.3000 175.3000 13.6000 ;
	    RECT 173.4000 11.1000 173.8000 13.3000 ;
	    RECT 174.9000 13.2000 175.3000 13.3000 ;
	    RECT 179.8000 12.8000 180.1000 13.9000 ;
	    RECT 181.4000 13.8000 182.2000 13.9000 ;
	    RECT 178.9000 12.7000 179.3000 12.8000 ;
	    RECT 175.8000 12.1000 176.2000 12.5000 ;
	    RECT 177.9000 12.4000 179.3000 12.7000 ;
	    RECT 179.8000 12.4000 180.2000 12.8000 ;
	    RECT 177.9000 12.1000 178.2000 12.4000 ;
	    RECT 180.6000 12.1000 181.0000 12.5000 ;
	    RECT 175.5000 11.8000 176.2000 12.1000 ;
	    RECT 175.5000 11.1000 176.1000 11.8000 ;
	    RECT 177.8000 11.1000 178.2000 12.1000 ;
	    RECT 180.0000 11.8000 181.0000 12.1000 ;
	    RECT 180.0000 11.1000 180.4000 11.8000 ;
	    RECT 182.2000 11.1000 182.6000 13.5000 ;
	    RECT 183.0000 12.4000 183.4000 13.2000 ;
	    RECT 183.8000 13.1000 184.2000 19.9000 ;
	    RECT 185.9000 16.3000 186.3000 19.9000 ;
	    RECT 185.4000 15.9000 186.3000 16.3000 ;
	    RECT 187.3000 16.3000 187.7000 19.9000 ;
	    RECT 190.2000 17.9000 190.6000 19.9000 ;
	    RECT 187.3000 15.9000 188.2000 16.3000 ;
	    RECT 184.6000 14.8000 185.0000 15.2000 ;
	    RECT 184.6000 14.1000 184.9000 14.8000 ;
	    RECT 185.5000 14.2000 185.8000 15.9000 ;
	    RECT 186.2000 14.8000 186.6000 15.6000 ;
	    RECT 187.8000 15.1000 188.1000 15.9000 ;
	    RECT 190.3000 15.8000 190.6000 17.9000 ;
	    RECT 191.8000 15.9000 192.2000 19.9000 ;
	    RECT 193.9000 16.2000 194.3000 19.9000 ;
	    RECT 193.9000 15.9000 194.4000 16.2000 ;
	    RECT 190.3000 15.5000 191.5000 15.8000 ;
	    RECT 187.8000 14.8000 188.9000 15.1000 ;
	    RECT 185.4000 14.1000 185.8000 14.2000 ;
	    RECT 184.6000 13.8000 185.8000 14.1000 ;
	    RECT 184.6000 13.1000 185.0000 13.2000 ;
	    RECT 183.8000 12.8000 185.0000 13.1000 ;
	    RECT 183.8000 11.1000 184.2000 12.8000 ;
	    RECT 184.6000 12.4000 185.0000 12.8000 ;
	    RECT 185.5000 12.1000 185.8000 13.8000 ;
	    RECT 185.4000 11.1000 185.8000 12.1000 ;
	    RECT 187.8000 14.2000 188.1000 14.8000 ;
	    RECT 188.6000 14.2000 188.9000 14.8000 ;
	    RECT 187.8000 13.8000 188.2000 14.2000 ;
	    RECT 188.6000 13.8000 189.0000 14.2000 ;
	    RECT 189.4000 13.8000 189.8000 14.6000 ;
	    RECT 191.2000 13.8000 191.5000 15.5000 ;
	    RECT 191.9000 15.2000 192.2000 15.9000 ;
	    RECT 191.8000 15.1000 192.2000 15.2000 ;
	    RECT 191.8000 14.8000 192.9000 15.1000 ;
	    RECT 187.8000 12.1000 188.1000 13.8000 ;
	    RECT 191.2000 13.7000 191.6000 13.8000 ;
	    RECT 190.1000 13.5000 191.6000 13.7000 ;
	    RECT 189.5000 13.4000 191.6000 13.5000 ;
	    RECT 189.5000 13.2000 190.4000 13.4000 ;
	    RECT 188.6000 12.4000 189.0000 13.2000 ;
	    RECT 189.5000 13.1000 189.8000 13.2000 ;
	    RECT 191.9000 13.1000 192.2000 14.8000 ;
	    RECT 192.6000 14.2000 192.9000 14.8000 ;
	    RECT 193.4000 14.4000 193.8000 15.2000 ;
	    RECT 194.1000 14.2000 194.4000 15.9000 ;
	    RECT 195.8000 15.7000 196.2000 19.9000 ;
	    RECT 198.0000 18.2000 198.4000 19.9000 ;
	    RECT 197.4000 17.9000 198.4000 18.2000 ;
	    RECT 200.2000 17.9000 200.6000 19.9000 ;
	    RECT 202.3000 17.9000 202.9000 19.9000 ;
	    RECT 197.4000 17.5000 197.8000 17.9000 ;
	    RECT 200.2000 17.6000 200.5000 17.9000 ;
	    RECT 199.1000 17.3000 200.9000 17.6000 ;
	    RECT 202.2000 17.5000 202.6000 17.9000 ;
	    RECT 199.1000 17.2000 199.5000 17.3000 ;
	    RECT 200.5000 17.2000 200.9000 17.3000 ;
	    RECT 197.4000 16.5000 197.8000 16.6000 ;
	    RECT 199.7000 16.5000 200.1000 16.6000 ;
	    RECT 197.4000 16.2000 200.1000 16.5000 ;
	    RECT 200.4000 16.5000 201.5000 16.8000 ;
	    RECT 200.4000 15.9000 200.7000 16.5000 ;
	    RECT 201.1000 16.4000 201.5000 16.5000 ;
	    RECT 202.3000 16.6000 203.0000 17.0000 ;
	    RECT 202.3000 16.1000 202.6000 16.6000 ;
	    RECT 198.3000 15.7000 200.7000 15.9000 ;
	    RECT 195.8000 15.6000 200.7000 15.7000 ;
	    RECT 201.4000 15.8000 202.6000 16.1000 ;
	    RECT 195.8000 15.5000 198.7000 15.6000 ;
	    RECT 195.8000 15.4000 198.6000 15.5000 ;
	    RECT 199.0000 15.1000 199.4000 15.2000 ;
	    RECT 196.9000 14.8000 199.4000 15.1000 ;
	    RECT 196.9000 14.7000 197.3000 14.8000 ;
	    RECT 197.7000 14.2000 198.1000 14.3000 ;
	    RECT 201.4000 14.2000 201.7000 15.8000 ;
	    RECT 204.6000 15.6000 205.0000 19.9000 ;
	    RECT 207.3000 16.4000 207.7000 19.9000 ;
	    RECT 209.4000 17.5000 209.8000 19.5000 ;
	    RECT 206.9000 16.1000 207.7000 16.4000 ;
	    RECT 202.9000 15.3000 205.0000 15.6000 ;
	    RECT 202.9000 15.2000 203.3000 15.3000 ;
	    RECT 203.7000 14.9000 204.1000 15.0000 ;
	    RECT 202.2000 14.6000 204.1000 14.9000 ;
	    RECT 202.2000 14.5000 202.6000 14.6000 ;
	    RECT 192.6000 14.1000 193.0000 14.2000 ;
	    RECT 192.6000 13.8000 193.4000 14.1000 ;
	    RECT 194.1000 13.8000 195.4000 14.2000 ;
	    RECT 196.2000 13.9000 201.7000 14.2000 ;
	    RECT 196.2000 13.8000 197.0000 13.9000 ;
	    RECT 198.2000 13.8000 198.6000 13.9000 ;
	    RECT 201.1000 13.8000 201.5000 13.9000 ;
	    RECT 193.0000 13.6000 193.4000 13.8000 ;
	    RECT 192.7000 13.1000 194.5000 13.3000 ;
	    RECT 195.0000 13.1000 195.3000 13.8000 ;
	    RECT 187.8000 11.1000 188.2000 12.1000 ;
	    RECT 189.4000 11.1000 189.8000 13.1000 ;
	    RECT 191.5000 12.6000 192.2000 13.1000 ;
	    RECT 192.6000 13.0000 194.6000 13.1000 ;
	    RECT 191.5000 11.1000 191.9000 12.6000 ;
	    RECT 192.6000 11.1000 193.0000 13.0000 ;
	    RECT 194.2000 11.1000 194.6000 13.0000 ;
	    RECT 195.0000 11.1000 195.4000 13.1000 ;
	    RECT 195.8000 11.1000 196.2000 13.5000 ;
	    RECT 198.3000 12.8000 198.6000 13.8000 ;
	    RECT 204.6000 13.6000 205.0000 15.3000 ;
	    RECT 205.4000 15.1000 205.8000 15.2000 ;
	    RECT 206.2000 15.1000 206.6000 15.6000 ;
	    RECT 205.4000 14.8000 206.6000 15.1000 ;
	    RECT 206.9000 14.2000 207.2000 16.1000 ;
	    RECT 209.5000 15.8000 209.8000 17.5000 ;
	    RECT 207.9000 15.5000 209.8000 15.8000 ;
	    RECT 207.9000 14.5000 208.2000 15.5000 ;
	    RECT 206.2000 13.8000 207.2000 14.2000 ;
	    RECT 207.5000 14.1000 208.2000 14.5000 ;
	    RECT 208.6000 14.4000 209.0000 15.2000 ;
	    RECT 209.4000 14.4000 209.8000 15.2000 ;
	    RECT 210.2000 15.1000 210.6000 15.2000 ;
	    RECT 211.0000 15.1000 211.4000 19.9000 ;
	    RECT 214.5000 19.2000 214.9000 19.9000 ;
	    RECT 214.5000 18.8000 215.4000 19.2000 ;
	    RECT 213.8000 16.8000 214.2000 17.2000 ;
	    RECT 213.8000 16.2000 214.1000 16.8000 ;
	    RECT 214.5000 16.2000 214.9000 18.8000 ;
	    RECT 213.4000 15.9000 214.1000 16.2000 ;
	    RECT 214.4000 15.9000 214.9000 16.2000 ;
	    RECT 213.4000 15.8000 213.8000 15.9000 ;
	    RECT 210.2000 14.8000 211.4000 15.1000 ;
	    RECT 203.1000 13.3000 205.0000 13.6000 ;
	    RECT 203.1000 13.2000 203.5000 13.3000 ;
	    RECT 197.4000 12.1000 197.8000 12.5000 ;
	    RECT 198.2000 12.4000 198.6000 12.8000 ;
	    RECT 199.1000 12.7000 199.5000 12.8000 ;
	    RECT 199.1000 12.4000 200.5000 12.7000 ;
	    RECT 200.2000 12.1000 200.5000 12.4000 ;
	    RECT 202.2000 12.1000 202.6000 12.5000 ;
	    RECT 197.4000 11.8000 198.4000 12.1000 ;
	    RECT 198.0000 11.1000 198.4000 11.8000 ;
	    RECT 200.2000 11.1000 200.6000 12.1000 ;
	    RECT 202.2000 11.8000 202.9000 12.1000 ;
	    RECT 202.3000 11.1000 202.9000 11.8000 ;
	    RECT 204.6000 11.1000 205.0000 13.3000 ;
	    RECT 206.9000 13.5000 207.2000 13.8000 ;
	    RECT 207.7000 13.9000 208.2000 14.1000 ;
	    RECT 207.7000 13.6000 209.8000 13.9000 ;
	    RECT 206.9000 13.3000 207.3000 13.5000 ;
	    RECT 206.9000 13.0000 207.7000 13.3000 ;
	    RECT 207.3000 11.5000 207.7000 13.0000 ;
	    RECT 209.5000 12.5000 209.8000 13.6000 ;
	    RECT 210.2000 13.4000 210.6000 14.2000 ;
	    RECT 209.4000 11.5000 209.8000 12.5000 ;
	    RECT 211.0000 11.1000 211.4000 14.8000 ;
	    RECT 214.4000 14.2000 214.7000 15.9000 ;
	    RECT 217.4000 15.1000 217.8000 19.9000 ;
	    RECT 219.8000 17.9000 220.2000 19.9000 ;
	    RECT 219.9000 15.8000 220.2000 17.9000 ;
	    RECT 221.4000 15.9000 221.8000 19.9000 ;
	    RECT 222.5000 17.2000 222.9000 19.9000 ;
	    RECT 222.2000 16.8000 222.9000 17.2000 ;
	    RECT 222.5000 16.3000 222.9000 16.8000 ;
	    RECT 222.5000 15.9000 223.4000 16.3000 ;
	    RECT 219.9000 15.5000 221.1000 15.8000 ;
	    RECT 217.4000 14.8000 218.5000 15.1000 ;
	    RECT 219.8000 14.8000 220.2000 15.2000 ;
	    RECT 213.4000 13.8000 214.7000 14.2000 ;
	    RECT 215.8000 14.1000 216.2000 14.2000 ;
	    RECT 215.4000 13.8000 216.2000 14.1000 ;
	    RECT 213.5000 13.1000 213.8000 13.8000 ;
	    RECT 215.4000 13.6000 215.8000 13.8000 ;
	    RECT 216.6000 13.4000 217.0000 14.2000 ;
	    RECT 214.3000 13.1000 216.1000 13.3000 ;
	    RECT 217.4000 13.1000 217.8000 14.8000 ;
	    RECT 218.2000 14.2000 218.5000 14.8000 ;
	    RECT 218.2000 13.8000 218.6000 14.2000 ;
	    RECT 219.0000 13.8000 219.4000 14.6000 ;
	    RECT 219.9000 14.4000 220.2000 14.8000 ;
	    RECT 219.9000 14.1000 220.4000 14.4000 ;
	    RECT 220.0000 14.0000 220.4000 14.1000 ;
	    RECT 220.8000 13.8000 221.1000 15.5000 ;
	    RECT 221.5000 15.2000 221.8000 15.9000 ;
	    RECT 221.4000 14.8000 221.8000 15.2000 ;
	    RECT 222.2000 14.8000 222.6000 15.6000 ;
	    RECT 220.8000 13.7000 221.2000 13.8000 ;
	    RECT 219.7000 13.5000 221.2000 13.7000 ;
	    RECT 219.1000 13.4000 221.2000 13.5000 ;
	    RECT 219.1000 13.2000 220.0000 13.4000 ;
	    RECT 219.1000 13.1000 219.4000 13.2000 ;
	    RECT 221.5000 13.1000 221.8000 14.8000 ;
	    RECT 213.4000 11.1000 213.8000 13.1000 ;
	    RECT 214.2000 13.0000 216.2000 13.1000 ;
	    RECT 214.2000 11.1000 214.6000 13.0000 ;
	    RECT 215.8000 11.1000 216.2000 13.0000 ;
	    RECT 217.4000 12.8000 218.3000 13.1000 ;
	    RECT 217.9000 11.1000 218.3000 12.8000 ;
	    RECT 219.0000 11.1000 219.4000 13.1000 ;
	    RECT 221.1000 12.6000 221.8000 13.1000 ;
	    RECT 223.0000 14.2000 223.3000 15.9000 ;
	    RECT 224.6000 15.8000 225.0000 16.6000 ;
	    RECT 224.6000 15.1000 225.0000 15.2000 ;
	    RECT 225.4000 15.1000 225.8000 19.9000 ;
	    RECT 228.3000 17.2000 228.7000 19.9000 ;
	    RECT 228.3000 16.8000 229.0000 17.2000 ;
	    RECT 228.3000 16.3000 228.7000 16.8000 ;
	    RECT 227.8000 15.9000 228.7000 16.3000 ;
	    RECT 224.6000 14.8000 225.8000 15.1000 ;
	    RECT 223.0000 13.8000 223.4000 14.2000 ;
	    RECT 221.1000 12.2000 221.5000 12.6000 ;
	    RECT 221.1000 11.8000 221.8000 12.2000 ;
	    RECT 223.0000 12.1000 223.3000 13.8000 ;
	    RECT 223.8000 12.4000 224.2000 13.2000 ;
	    RECT 225.4000 13.1000 225.8000 14.8000 ;
	    RECT 227.9000 14.2000 228.2000 15.9000 ;
	    RECT 228.6000 14.8000 229.0000 15.6000 ;
	    RECT 226.2000 13.4000 226.6000 14.2000 ;
	    RECT 227.8000 13.8000 228.2000 14.2000 ;
	    RECT 224.9000 12.8000 225.8000 13.1000 ;
	    RECT 221.1000 11.1000 221.5000 11.8000 ;
	    RECT 223.0000 11.1000 223.4000 12.1000 ;
	    RECT 224.9000 11.1000 225.3000 12.8000 ;
	    RECT 227.9000 12.1000 228.2000 13.8000 ;
	    RECT 229.4000 13.4000 229.8000 14.2000 ;
	    RECT 230.2000 13.1000 230.6000 19.9000 ;
	    RECT 231.0000 15.8000 231.4000 16.6000 ;
	    RECT 232.6000 15.1000 233.0000 19.9000 ;
	    RECT 233.4000 19.6000 235.4000 19.9000 ;
	    RECT 233.4000 15.9000 233.8000 19.6000 ;
	    RECT 234.2000 15.9000 234.6000 19.3000 ;
	    RECT 235.0000 16.2000 235.4000 19.6000 ;
	    RECT 236.6000 16.2000 237.0000 19.9000 ;
	    RECT 237.8000 16.8000 238.2000 17.2000 ;
	    RECT 237.8000 16.2000 238.1000 16.8000 ;
	    RECT 238.5000 16.2000 238.9000 19.9000 ;
	    RECT 235.0000 15.9000 237.0000 16.2000 ;
	    RECT 237.4000 15.9000 238.1000 16.2000 ;
	    RECT 238.4000 15.9000 238.9000 16.2000 ;
	    RECT 240.9000 16.3000 241.3000 19.9000 ;
	    RECT 240.9000 15.9000 241.8000 16.3000 ;
	    RECT 234.3000 15.6000 234.6000 15.9000 ;
	    RECT 237.4000 15.8000 237.8000 15.9000 ;
	    RECT 233.4000 15.1000 233.8000 15.6000 ;
	    RECT 234.3000 15.3000 235.3000 15.6000 ;
	    RECT 232.6000 14.8000 233.8000 15.1000 ;
	    RECT 235.0000 15.2000 235.3000 15.3000 ;
	    RECT 236.2000 15.2000 236.6000 15.4000 ;
	    RECT 235.0000 14.8000 235.4000 15.2000 ;
	    RECT 236.2000 14.9000 237.0000 15.2000 ;
	    RECT 236.6000 14.8000 237.0000 14.9000 ;
	    RECT 231.8000 13.1000 232.2000 13.2000 ;
	    RECT 230.2000 12.8000 232.2000 13.1000 ;
	    RECT 227.8000 11.1000 228.2000 12.1000 ;
	    RECT 230.7000 11.1000 231.1000 12.8000 ;
	    RECT 231.8000 12.4000 232.2000 12.8000 ;
	    RECT 232.6000 11.1000 233.0000 14.8000 ;
	    RECT 234.3000 14.4000 234.7000 14.8000 ;
	    RECT 234.3000 14.2000 234.6000 14.4000 ;
	    RECT 234.2000 13.8000 234.6000 14.2000 ;
	    RECT 235.0000 13.1000 235.3000 14.8000 ;
	    RECT 235.8000 14.1000 236.2000 14.6000 ;
	    RECT 238.4000 14.2000 238.7000 15.9000 ;
	    RECT 239.0000 14.4000 239.4000 15.2000 ;
	    RECT 240.6000 14.8000 241.0000 15.6000 ;
	    RECT 241.4000 14.2000 241.7000 15.9000 ;
	    RECT 243.0000 15.8000 243.4000 16.6000 ;
	    RECT 237.4000 14.1000 238.7000 14.2000 ;
	    RECT 239.8000 14.1000 240.2000 14.2000 ;
	    RECT 240.6000 14.1000 241.0000 14.2000 ;
	    RECT 235.8000 13.8000 238.7000 14.1000 ;
	    RECT 239.4000 13.8000 241.0000 14.1000 ;
	    RECT 241.4000 13.8000 241.8000 14.2000 ;
	    RECT 242.2000 13.8000 242.6000 14.2000 ;
	    RECT 237.5000 13.1000 237.8000 13.8000 ;
	    RECT 239.4000 13.6000 239.8000 13.8000 ;
	    RECT 238.3000 13.1000 240.1000 13.3000 ;
	    RECT 234.7000 11.1000 235.5000 13.1000 ;
	    RECT 237.4000 11.1000 237.8000 13.1000 ;
	    RECT 238.2000 13.0000 240.2000 13.1000 ;
	    RECT 238.2000 11.1000 238.6000 13.0000 ;
	    RECT 239.8000 11.1000 240.2000 13.0000 ;
	    RECT 241.4000 12.2000 241.7000 13.8000 ;
	    RECT 242.2000 13.2000 242.5000 13.8000 ;
	    RECT 242.2000 12.4000 242.6000 13.2000 ;
	    RECT 243.8000 13.1000 244.2000 19.9000 ;
	    RECT 246.7000 19.2000 247.1000 19.9000 ;
	    RECT 246.2000 18.8000 247.1000 19.2000 ;
	    RECT 246.7000 16.2000 247.1000 18.8000 ;
	    RECT 247.4000 16.8000 247.8000 17.2000 ;
	    RECT 247.5000 16.2000 247.8000 16.8000 ;
	    RECT 246.7000 15.9000 247.2000 16.2000 ;
	    RECT 247.5000 15.9000 248.2000 16.2000 ;
	    RECT 246.2000 15.1000 246.6000 15.2000 ;
	    RECT 244.6000 14.8000 246.6000 15.1000 ;
	    RECT 244.6000 14.2000 244.9000 14.8000 ;
	    RECT 246.2000 14.4000 246.6000 14.8000 ;
	    RECT 246.9000 14.2000 247.2000 15.9000 ;
	    RECT 247.8000 15.8000 248.2000 15.9000 ;
	    RECT 244.6000 13.4000 245.0000 14.2000 ;
	    RECT 245.4000 14.1000 245.8000 14.2000 ;
	    RECT 245.4000 13.8000 246.2000 14.1000 ;
	    RECT 246.9000 13.8000 248.2000 14.2000 ;
	    RECT 245.8000 13.6000 246.2000 13.8000 ;
	    RECT 245.5000 13.1000 247.3000 13.3000 ;
	    RECT 247.8000 13.1000 248.1000 13.8000 ;
	    RECT 243.3000 12.8000 244.2000 13.1000 ;
	    RECT 245.4000 13.0000 247.4000 13.1000 ;
	    RECT 243.3000 12.2000 243.7000 12.8000 ;
	    RECT 241.4000 11.1000 241.8000 12.2000 ;
	    RECT 243.3000 11.8000 244.2000 12.2000 ;
	    RECT 243.3000 11.1000 243.7000 11.8000 ;
	    RECT 245.4000 11.1000 245.8000 13.0000 ;
	    RECT 247.0000 11.1000 247.4000 13.0000 ;
	    RECT 247.8000 11.1000 248.2000 13.1000 ;
	    RECT 248.6000 11.1000 249.0000 19.9000 ;
	    RECT 250.2000 13.4000 250.6000 14.2000 ;
	    RECT 251.0000 11.1000 251.4000 19.9000 ;
	    RECT 252.1000 16.3000 252.5000 19.9000 ;
	    RECT 252.1000 15.9000 253.0000 16.3000 ;
	    RECT 252.6000 15.8000 253.0000 15.9000 ;
	    RECT 251.8000 14.8000 252.2000 15.6000 ;
	    RECT 252.6000 14.2000 252.9000 15.8000 ;
	    RECT 252.6000 13.8000 253.0000 14.2000 ;
	    RECT 252.6000 12.1000 252.9000 13.8000 ;
	    RECT 253.4000 13.1000 253.8000 13.2000 ;
	    RECT 254.2000 13.1000 254.6000 19.9000 ;
	    RECT 253.4000 12.8000 254.6000 13.1000 ;
	    RECT 253.4000 12.4000 253.8000 12.8000 ;
	    RECT 252.6000 11.1000 253.0000 12.1000 ;
	    RECT 254.2000 11.1000 254.6000 12.8000 ;
	    RECT 255.0000 12.4000 255.4000 13.2000 ;
	    RECT 255.8000 11.1000 256.2000 19.9000 ;
	    RECT 257.4000 15.9000 257.8000 19.9000 ;
	    RECT 258.2000 16.2000 258.6000 19.9000 ;
	    RECT 259.8000 16.2000 260.2000 19.9000 ;
	    RECT 258.2000 15.9000 260.2000 16.2000 ;
	    RECT 257.5000 15.2000 257.8000 15.9000 ;
	    RECT 260.6000 15.7000 261.0000 19.9000 ;
	    RECT 262.8000 18.2000 263.2000 19.9000 ;
	    RECT 262.2000 17.9000 263.2000 18.2000 ;
	    RECT 265.0000 17.9000 265.4000 19.9000 ;
	    RECT 267.1000 17.9000 267.7000 19.9000 ;
	    RECT 262.2000 17.5000 262.6000 17.9000 ;
	    RECT 265.0000 17.6000 265.3000 17.9000 ;
	    RECT 263.9000 17.3000 265.7000 17.6000 ;
	    RECT 267.0000 17.5000 267.4000 17.9000 ;
	    RECT 263.9000 17.2000 264.3000 17.3000 ;
	    RECT 265.3000 17.2000 265.7000 17.3000 ;
	    RECT 262.2000 16.5000 262.6000 16.6000 ;
	    RECT 264.5000 16.5000 264.9000 16.6000 ;
	    RECT 262.2000 16.2000 264.9000 16.5000 ;
	    RECT 265.2000 16.5000 266.3000 16.8000 ;
	    RECT 265.2000 15.9000 265.5000 16.5000 ;
	    RECT 265.9000 16.4000 266.3000 16.5000 ;
	    RECT 267.1000 16.6000 267.8000 17.0000 ;
	    RECT 267.1000 16.1000 267.4000 16.6000 ;
	    RECT 263.1000 15.7000 265.5000 15.9000 ;
	    RECT 260.6000 15.6000 265.5000 15.7000 ;
	    RECT 266.2000 15.8000 267.4000 16.1000 ;
	    RECT 260.6000 15.5000 263.5000 15.6000 ;
	    RECT 260.6000 15.4000 263.4000 15.5000 ;
	    RECT 257.4000 14.9000 258.6000 15.2000 ;
	    RECT 263.8000 15.1000 264.2000 15.2000 ;
	    RECT 257.4000 14.8000 257.8000 14.9000 ;
	    RECT 256.6000 12.4000 257.0000 13.2000 ;
	    RECT 257.4000 12.8000 257.8000 13.2000 ;
	    RECT 258.3000 13.1000 258.6000 14.9000 ;
	    RECT 261.7000 14.8000 264.2000 15.1000 ;
	    RECT 261.7000 14.7000 262.1000 14.8000 ;
	    RECT 259.0000 13.8000 259.4000 14.6000 ;
	    RECT 262.5000 14.2000 262.9000 14.3000 ;
	    RECT 266.2000 14.2000 266.5000 15.8000 ;
	    RECT 269.4000 15.6000 269.8000 19.9000 ;
	    RECT 267.7000 15.3000 269.8000 15.6000 ;
	    RECT 267.7000 15.2000 268.1000 15.3000 ;
	    RECT 268.5000 14.9000 268.9000 15.0000 ;
	    RECT 267.0000 14.6000 268.9000 14.9000 ;
	    RECT 267.0000 14.5000 267.4000 14.6000 ;
	    RECT 261.0000 13.9000 266.5000 14.2000 ;
	    RECT 261.0000 13.8000 261.8000 13.9000 ;
	    RECT 257.5000 12.4000 257.9000 12.8000 ;
	    RECT 258.2000 11.1000 258.6000 13.1000 ;
	    RECT 260.6000 11.1000 261.0000 13.5000 ;
	    RECT 263.1000 12.8000 263.4000 13.9000 ;
	    RECT 265.9000 13.8000 266.3000 13.9000 ;
	    RECT 269.4000 13.6000 269.8000 15.3000 ;
	    RECT 267.9000 13.3000 269.8000 13.6000 ;
	    RECT 267.9000 13.2000 268.3000 13.3000 ;
	    RECT 262.2000 12.1000 262.6000 12.5000 ;
	    RECT 263.0000 12.4000 263.4000 12.8000 ;
	    RECT 263.9000 12.7000 264.3000 12.8000 ;
	    RECT 263.9000 12.4000 265.3000 12.7000 ;
	    RECT 265.0000 12.1000 265.3000 12.4000 ;
	    RECT 267.0000 12.1000 267.4000 12.5000 ;
	    RECT 262.2000 11.8000 263.2000 12.1000 ;
	    RECT 262.8000 11.1000 263.2000 11.8000 ;
	    RECT 265.0000 11.1000 265.4000 12.1000 ;
	    RECT 267.0000 11.8000 267.7000 12.1000 ;
	    RECT 267.1000 11.1000 267.7000 11.8000 ;
	    RECT 269.4000 11.1000 269.8000 13.3000 ;
	    RECT 2.2000 7.6000 2.6000 9.9000 ;
	    RECT 4.6000 7.6000 5.0000 9.9000 ;
	    RECT 5.4000 7.8000 5.8000 8.6000 ;
	    RECT 6.2000 8.1000 6.6000 9.9000 ;
	    RECT 7.8000 8.9000 8.2000 9.9000 ;
	    RECT 7.0000 8.1000 7.4000 8.6000 ;
	    RECT 6.2000 7.8000 7.4000 8.1000 ;
	    RECT 1.5000 7.3000 2.6000 7.6000 ;
	    RECT 3.9000 7.3000 5.0000 7.6000 ;
	    RECT 1.5000 5.8000 1.8000 7.3000 ;
	    RECT 2.2000 5.8000 2.6000 6.6000 ;
	    RECT 3.9000 5.8000 4.2000 7.3000 ;
	    RECT 4.6000 6.1000 5.0000 6.6000 ;
	    RECT 5.4000 6.1000 5.8000 6.2000 ;
	    RECT 4.6000 5.8000 5.8000 6.1000 ;
	    RECT 1.2000 5.4000 1.8000 5.8000 ;
	    RECT 3.6000 5.4000 4.2000 5.8000 ;
	    RECT 1.5000 5.1000 1.8000 5.4000 ;
	    RECT 3.9000 5.1000 4.2000 5.4000 ;
	    RECT 1.5000 4.8000 2.6000 5.1000 ;
	    RECT 3.9000 4.8000 5.0000 5.1000 ;
	    RECT 2.2000 1.1000 2.6000 4.8000 ;
	    RECT 4.6000 1.1000 5.0000 4.8000 ;
	    RECT 6.2000 1.1000 6.6000 7.8000 ;
	    RECT 7.9000 7.2000 8.2000 8.9000 ;
	    RECT 7.8000 6.8000 8.2000 7.2000 ;
	    RECT 7.9000 5.1000 8.2000 6.8000 ;
	    RECT 9.4000 7.7000 9.8000 9.9000 ;
	    RECT 11.5000 9.2000 12.1000 9.9000 ;
	    RECT 11.5000 8.9000 12.2000 9.2000 ;
	    RECT 13.8000 8.9000 14.2000 9.9000 ;
	    RECT 16.0000 9.2000 16.4000 9.9000 ;
	    RECT 16.0000 8.9000 17.0000 9.2000 ;
	    RECT 11.8000 8.5000 12.2000 8.9000 ;
	    RECT 13.9000 8.6000 14.2000 8.9000 ;
	    RECT 13.9000 8.3000 15.3000 8.6000 ;
	    RECT 14.9000 8.2000 15.3000 8.3000 ;
	    RECT 15.8000 7.8000 16.2000 8.6000 ;
	    RECT 16.6000 8.5000 17.0000 8.9000 ;
	    RECT 10.9000 7.7000 11.3000 7.8000 ;
	    RECT 9.4000 7.4000 11.3000 7.7000 ;
	    RECT 8.6000 5.4000 9.0000 6.2000 ;
	    RECT 9.4000 5.7000 9.8000 7.4000 ;
	    RECT 12.9000 7.1000 13.3000 7.2000 ;
	    RECT 15.8000 7.1000 16.1000 7.8000 ;
	    RECT 18.2000 7.5000 18.6000 9.9000 ;
	    RECT 20.6000 7.6000 21.0000 9.9000 ;
	    RECT 19.9000 7.3000 21.0000 7.6000 ;
	    RECT 22.2000 8.9000 22.6000 9.9000 ;
	    RECT 17.4000 7.1000 18.2000 7.2000 ;
	    RECT 12.7000 6.8000 18.2000 7.1000 ;
	    RECT 11.8000 6.4000 12.2000 6.5000 ;
	    RECT 10.3000 6.1000 12.2000 6.4000 ;
	    RECT 10.3000 6.0000 10.7000 6.1000 ;
	    RECT 11.1000 5.7000 11.5000 5.8000 ;
	    RECT 9.4000 5.4000 11.5000 5.7000 ;
	    RECT 7.8000 4.7000 8.7000 5.1000 ;
	    RECT 8.3000 4.2000 8.7000 4.7000 ;
	    RECT 8.3000 3.8000 9.0000 4.2000 ;
	    RECT 8.3000 1.1000 8.7000 3.8000 ;
	    RECT 9.4000 1.1000 9.8000 5.4000 ;
	    RECT 12.7000 5.2000 13.0000 6.8000 ;
	    RECT 16.3000 6.7000 16.7000 6.8000 ;
	    RECT 17.1000 6.2000 17.5000 6.3000 ;
	    RECT 15.0000 5.9000 17.5000 6.2000 ;
	    RECT 15.0000 5.8000 15.4000 5.9000 ;
	    RECT 19.9000 5.8000 20.2000 7.3000 ;
	    RECT 22.2000 7.2000 22.5000 8.9000 ;
	    RECT 23.0000 8.1000 23.4000 8.6000 ;
	    RECT 23.8000 8.1000 24.2000 9.9000 ;
	    RECT 23.0000 7.8000 24.2000 8.1000 ;
	    RECT 22.2000 6.8000 22.6000 7.2000 ;
	    RECT 20.6000 5.8000 21.0000 6.6000 ;
	    RECT 15.8000 5.5000 18.6000 5.6000 ;
	    RECT 15.7000 5.4000 18.6000 5.5000 ;
	    RECT 19.6000 5.4000 20.2000 5.8000 ;
	    RECT 21.4000 5.4000 21.8000 6.2000 ;
	    RECT 11.8000 4.9000 13.0000 5.2000 ;
	    RECT 13.7000 5.3000 18.6000 5.4000 ;
	    RECT 13.7000 5.1000 16.1000 5.3000 ;
	    RECT 11.8000 4.4000 12.1000 4.9000 ;
	    RECT 11.4000 4.0000 12.1000 4.4000 ;
	    RECT 12.9000 4.5000 13.3000 4.6000 ;
	    RECT 13.7000 4.5000 14.0000 5.1000 ;
	    RECT 12.9000 4.2000 14.0000 4.5000 ;
	    RECT 14.3000 4.5000 17.0000 4.8000 ;
	    RECT 14.3000 4.4000 14.7000 4.5000 ;
	    RECT 16.6000 4.4000 17.0000 4.5000 ;
	    RECT 13.5000 3.7000 13.9000 3.8000 ;
	    RECT 14.9000 3.7000 15.3000 3.8000 ;
	    RECT 11.8000 3.1000 12.2000 3.5000 ;
	    RECT 13.5000 3.4000 15.3000 3.7000 ;
	    RECT 13.9000 3.1000 14.2000 3.4000 ;
	    RECT 16.6000 3.1000 17.0000 3.5000 ;
	    RECT 11.5000 1.1000 12.1000 3.1000 ;
	    RECT 13.8000 1.1000 14.2000 3.1000 ;
	    RECT 16.0000 2.8000 17.0000 3.1000 ;
	    RECT 16.0000 1.1000 16.4000 2.8000 ;
	    RECT 18.2000 1.1000 18.6000 5.3000 ;
	    RECT 19.9000 5.1000 20.2000 5.4000 ;
	    RECT 22.2000 5.2000 22.5000 6.8000 ;
	    RECT 22.2000 5.1000 22.6000 5.2000 ;
	    RECT 19.9000 4.8000 21.0000 5.1000 ;
	    RECT 20.6000 1.1000 21.0000 4.8000 ;
	    RECT 21.7000 4.7000 22.6000 5.1000 ;
	    RECT 21.7000 1.1000 22.1000 4.7000 ;
	    RECT 23.8000 1.1000 24.2000 7.8000 ;
	    RECT 24.6000 7.8000 25.0000 8.6000 ;
	    RECT 24.6000 7.2000 24.9000 7.8000 ;
	    RECT 25.4000 7.5000 25.8000 9.9000 ;
	    RECT 27.6000 9.2000 28.0000 9.9000 ;
	    RECT 27.0000 8.9000 28.0000 9.2000 ;
	    RECT 29.8000 8.9000 30.2000 9.9000 ;
	    RECT 31.9000 9.2000 32.5000 9.9000 ;
	    RECT 31.8000 8.9000 32.5000 9.2000 ;
	    RECT 27.0000 8.5000 27.4000 8.9000 ;
	    RECT 29.8000 8.6000 30.1000 8.9000 ;
	    RECT 27.8000 7.8000 28.2000 8.6000 ;
	    RECT 28.7000 8.3000 30.1000 8.6000 ;
	    RECT 31.8000 8.5000 32.2000 8.9000 ;
	    RECT 28.7000 8.2000 29.1000 8.3000 ;
	    RECT 24.6000 6.8000 25.0000 7.2000 ;
	    RECT 25.8000 7.1000 26.6000 7.2000 ;
	    RECT 27.9000 7.1000 28.2000 7.8000 ;
	    RECT 32.7000 7.7000 33.1000 7.8000 ;
	    RECT 34.2000 7.7000 34.6000 9.9000 ;
	    RECT 32.7000 7.4000 34.6000 7.7000 ;
	    RECT 30.7000 7.1000 31.1000 7.2000 ;
	    RECT 25.8000 6.8000 31.3000 7.1000 ;
	    RECT 27.3000 6.7000 27.7000 6.8000 ;
	    RECT 26.5000 6.2000 26.9000 6.3000 ;
	    RECT 27.8000 6.2000 28.2000 6.3000 ;
	    RECT 26.5000 5.9000 29.0000 6.2000 ;
	    RECT 28.6000 5.8000 29.0000 5.9000 ;
	    RECT 25.4000 5.5000 28.2000 5.6000 ;
	    RECT 25.4000 5.4000 28.3000 5.5000 ;
	    RECT 25.4000 5.3000 30.3000 5.4000 ;
	    RECT 25.4000 1.1000 25.8000 5.3000 ;
	    RECT 27.9000 5.1000 30.3000 5.3000 ;
	    RECT 27.0000 4.5000 29.7000 4.8000 ;
	    RECT 27.0000 4.4000 27.4000 4.5000 ;
	    RECT 29.3000 4.4000 29.7000 4.5000 ;
	    RECT 30.0000 4.5000 30.3000 5.1000 ;
	    RECT 31.0000 5.2000 31.3000 6.8000 ;
	    RECT 31.8000 6.4000 32.2000 6.5000 ;
	    RECT 31.8000 6.1000 33.7000 6.4000 ;
	    RECT 33.3000 6.0000 33.7000 6.1000 ;
	    RECT 34.2000 6.1000 34.6000 7.4000 ;
	    RECT 35.0000 7.6000 35.4000 9.9000 ;
	    RECT 38.2000 8.9000 38.6000 9.9000 ;
	    RECT 35.0000 7.3000 36.1000 7.6000 ;
	    RECT 35.0000 6.1000 35.4000 6.6000 ;
	    RECT 34.2000 5.8000 35.4000 6.1000 ;
	    RECT 35.8000 5.8000 36.1000 7.3000 ;
	    RECT 38.2000 7.2000 38.5000 8.9000 ;
	    RECT 39.0000 8.1000 39.4000 8.6000 ;
	    RECT 39.8000 8.1000 40.2000 9.9000 ;
	    RECT 39.0000 7.8000 40.2000 8.1000 ;
	    RECT 38.2000 6.8000 38.6000 7.2000 ;
	    RECT 39.0000 6.8000 39.4000 7.2000 ;
	    RECT 32.5000 5.7000 32.9000 5.8000 ;
	    RECT 34.2000 5.7000 34.6000 5.8000 ;
	    RECT 32.5000 5.4000 34.6000 5.7000 ;
	    RECT 31.0000 4.9000 32.2000 5.2000 ;
	    RECT 30.7000 4.5000 31.1000 4.6000 ;
	    RECT 30.0000 4.2000 31.1000 4.5000 ;
	    RECT 31.9000 4.4000 32.2000 4.9000 ;
	    RECT 31.9000 4.0000 32.6000 4.4000 ;
	    RECT 28.7000 3.7000 29.1000 3.8000 ;
	    RECT 30.1000 3.7000 30.5000 3.8000 ;
	    RECT 27.0000 3.1000 27.4000 3.5000 ;
	    RECT 28.7000 3.4000 30.5000 3.7000 ;
	    RECT 29.8000 3.1000 30.1000 3.4000 ;
	    RECT 31.8000 3.1000 32.2000 3.5000 ;
	    RECT 27.0000 2.8000 28.0000 3.1000 ;
	    RECT 27.6000 1.1000 28.0000 2.8000 ;
	    RECT 29.8000 1.1000 30.2000 3.1000 ;
	    RECT 31.9000 1.1000 32.5000 3.1000 ;
	    RECT 34.2000 1.1000 34.6000 5.4000 ;
	    RECT 35.8000 5.4000 36.4000 5.8000 ;
	    RECT 37.4000 5.4000 37.8000 6.2000 ;
	    RECT 38.2000 6.1000 38.5000 6.8000 ;
	    RECT 39.0000 6.1000 39.3000 6.8000 ;
	    RECT 38.2000 5.8000 39.3000 6.1000 ;
	    RECT 35.8000 5.1000 36.1000 5.4000 ;
	    RECT 38.2000 5.1000 38.5000 5.8000 ;
	    RECT 35.0000 4.8000 36.1000 5.1000 ;
	    RECT 35.0000 1.1000 35.4000 4.8000 ;
	    RECT 37.7000 4.7000 38.6000 5.1000 ;
	    RECT 37.7000 1.1000 38.1000 4.7000 ;
	    RECT 39.8000 1.1000 40.2000 7.8000 ;
	    RECT 40.6000 7.8000 41.0000 8.6000 ;
	    RECT 40.6000 7.2000 40.9000 7.8000 ;
	    RECT 41.4000 7.5000 41.8000 9.9000 ;
	    RECT 43.6000 9.2000 44.0000 9.9000 ;
	    RECT 43.0000 8.9000 44.0000 9.2000 ;
	    RECT 45.8000 8.9000 46.2000 9.9000 ;
	    RECT 47.9000 9.2000 48.5000 9.9000 ;
	    RECT 47.8000 8.9000 48.5000 9.2000 ;
	    RECT 43.0000 8.5000 43.4000 8.9000 ;
	    RECT 45.8000 8.6000 46.1000 8.9000 ;
	    RECT 43.8000 7.8000 44.2000 8.6000 ;
	    RECT 44.7000 8.3000 46.1000 8.6000 ;
	    RECT 47.8000 8.5000 48.2000 8.9000 ;
	    RECT 44.7000 8.2000 45.1000 8.3000 ;
	    RECT 40.6000 6.8000 41.0000 7.2000 ;
	    RECT 41.8000 7.1000 42.6000 7.2000 ;
	    RECT 43.9000 7.1000 44.2000 7.8000 ;
	    RECT 48.7000 7.7000 49.1000 7.8000 ;
	    RECT 50.2000 7.7000 50.6000 9.9000 ;
	    RECT 48.7000 7.4000 50.6000 7.7000 ;
	    RECT 46.7000 7.1000 47.1000 7.2000 ;
	    RECT 41.8000 6.8000 47.3000 7.1000 ;
	    RECT 43.3000 6.7000 43.7000 6.8000 ;
	    RECT 42.5000 6.2000 42.9000 6.3000 ;
	    RECT 43.8000 6.2000 44.2000 6.3000 ;
	    RECT 42.5000 5.9000 45.0000 6.2000 ;
	    RECT 44.6000 5.8000 45.0000 5.9000 ;
	    RECT 41.4000 5.5000 44.2000 5.6000 ;
	    RECT 41.4000 5.4000 44.3000 5.5000 ;
	    RECT 41.4000 5.3000 46.3000 5.4000 ;
	    RECT 41.4000 1.1000 41.8000 5.3000 ;
	    RECT 43.9000 5.1000 46.3000 5.3000 ;
	    RECT 43.0000 4.5000 45.7000 4.8000 ;
	    RECT 43.0000 4.4000 43.4000 4.5000 ;
	    RECT 45.3000 4.4000 45.7000 4.5000 ;
	    RECT 46.0000 4.5000 46.3000 5.1000 ;
	    RECT 47.0000 5.2000 47.3000 6.8000 ;
	    RECT 47.8000 6.4000 48.2000 6.5000 ;
	    RECT 47.8000 6.1000 49.7000 6.4000 ;
	    RECT 49.3000 6.0000 49.7000 6.1000 ;
	    RECT 50.2000 6.1000 50.6000 7.4000 ;
	    RECT 51.0000 7.6000 51.4000 9.9000 ;
	    RECT 53.4000 7.9000 53.8000 9.9000 ;
	    RECT 55.6000 8.1000 56.4000 9.9000 ;
	    RECT 53.4000 7.6000 54.5000 7.9000 ;
	    RECT 55.0000 7.7000 55.8000 7.8000 ;
	    RECT 51.0000 7.3000 52.1000 7.6000 ;
	    RECT 54.1000 7.5000 54.5000 7.6000 ;
	    RECT 51.0000 6.1000 51.4000 6.6000 ;
	    RECT 50.2000 5.8000 51.4000 6.1000 ;
	    RECT 51.8000 5.8000 52.1000 7.3000 ;
	    RECT 54.8000 7.4000 55.8000 7.7000 ;
	    RECT 54.8000 7.2000 55.1000 7.4000 ;
	    RECT 53.4000 6.9000 55.1000 7.2000 ;
	    RECT 53.4000 6.8000 54.2000 6.9000 ;
	    RECT 55.4000 6.7000 55.8000 7.1000 ;
	    RECT 55.4000 6.4000 55.7000 6.7000 ;
	    RECT 54.4000 6.1000 55.7000 6.4000 ;
	    RECT 56.1000 6.4000 56.4000 8.1000 ;
	    RECT 58.2000 7.9000 58.6000 9.9000 ;
	    RECT 61.4000 8.8000 61.8000 9.9000 ;
	    RECT 56.7000 7.4000 57.1000 7.8000 ;
	    RECT 57.4000 7.6000 58.6000 7.9000 ;
	    RECT 60.6000 7.8000 61.0000 8.6000 ;
	    RECT 57.4000 7.5000 57.8000 7.6000 ;
	    RECT 56.8000 7.2000 57.1000 7.4000 ;
	    RECT 61.5000 7.2000 61.8000 8.8000 ;
	    RECT 56.8000 6.8000 57.2000 7.2000 ;
	    RECT 57.8000 6.8000 58.6000 7.2000 ;
	    RECT 61.4000 6.8000 61.8000 7.2000 ;
	    RECT 56.1000 6.2000 56.6000 6.4000 ;
	    RECT 56.1000 6.1000 57.0000 6.2000 ;
	    RECT 59.8000 6.1000 60.2000 6.2000 ;
	    RECT 54.4000 6.0000 54.8000 6.1000 ;
	    RECT 56.3000 5.8000 60.2000 6.1000 ;
	    RECT 48.5000 5.7000 48.9000 5.8000 ;
	    RECT 50.2000 5.7000 50.6000 5.8000 ;
	    RECT 48.5000 5.4000 50.6000 5.7000 ;
	    RECT 47.0000 4.9000 48.2000 5.2000 ;
	    RECT 46.7000 4.5000 47.1000 4.6000 ;
	    RECT 46.0000 4.2000 47.1000 4.5000 ;
	    RECT 47.9000 4.4000 48.2000 4.9000 ;
	    RECT 47.9000 4.0000 48.6000 4.4000 ;
	    RECT 44.7000 3.7000 45.1000 3.8000 ;
	    RECT 46.1000 3.7000 46.5000 3.8000 ;
	    RECT 43.0000 3.1000 43.4000 3.5000 ;
	    RECT 44.7000 3.4000 46.5000 3.7000 ;
	    RECT 45.8000 3.1000 46.1000 3.4000 ;
	    RECT 47.8000 3.1000 48.2000 3.5000 ;
	    RECT 43.0000 2.8000 44.0000 3.1000 ;
	    RECT 43.6000 1.1000 44.0000 2.8000 ;
	    RECT 45.8000 1.1000 46.2000 3.1000 ;
	    RECT 47.9000 1.1000 48.5000 3.1000 ;
	    RECT 50.2000 1.1000 50.6000 5.4000 ;
	    RECT 51.8000 5.4000 52.4000 5.8000 ;
	    RECT 55.5000 5.7000 55.9000 5.8000 ;
	    RECT 54.2000 5.4000 55.9000 5.7000 ;
	    RECT 51.8000 5.1000 52.1000 5.4000 ;
	    RECT 54.2000 5.1000 54.5000 5.4000 ;
	    RECT 56.3000 5.1000 56.6000 5.8000 ;
	    RECT 61.5000 5.1000 61.8000 6.8000 ;
	    RECT 62.2000 6.1000 62.6000 6.2000 ;
	    RECT 63.0000 6.1000 63.4000 9.9000 ;
	    RECT 63.8000 7.8000 64.2000 8.6000 ;
	    RECT 64.6000 7.9000 65.0000 9.9000 ;
	    RECT 66.8000 9.2000 67.6000 9.9000 ;
	    RECT 66.8000 8.8000 68.2000 9.2000 ;
	    RECT 66.8000 8.1000 67.6000 8.8000 ;
	    RECT 64.6000 7.6000 65.8000 7.9000 ;
	    RECT 65.4000 7.5000 65.8000 7.6000 ;
	    RECT 66.1000 7.4000 66.5000 7.8000 ;
	    RECT 66.1000 7.2000 66.4000 7.4000 ;
	    RECT 64.6000 6.8000 65.4000 7.2000 ;
	    RECT 66.0000 6.8000 66.4000 7.2000 ;
	    RECT 66.8000 7.1000 67.1000 8.1000 ;
	    RECT 69.4000 7.9000 69.8000 9.9000 ;
	    RECT 67.4000 7.4000 68.2000 7.8000 ;
	    RECT 68.5000 7.6000 69.8000 7.9000 ;
	    RECT 70.2000 7.9000 70.6000 9.9000 ;
	    RECT 72.4000 8.1000 73.2000 9.9000 ;
	    RECT 70.2000 7.6000 71.5000 7.9000 ;
	    RECT 68.5000 7.5000 68.9000 7.6000 ;
	    RECT 71.1000 7.5000 71.5000 7.6000 ;
	    RECT 71.8000 7.4000 72.6000 7.8000 ;
	    RECT 69.0000 7.1000 69.8000 7.2000 ;
	    RECT 66.8000 6.8000 67.3000 7.1000 ;
	    RECT 68.7000 7.0000 69.8000 7.1000 ;
	    RECT 62.2000 5.8000 63.4000 6.1000 ;
	    RECT 62.2000 5.4000 62.6000 5.8000 ;
	    RECT 51.0000 4.8000 52.1000 5.1000 ;
	    RECT 53.4000 4.8000 54.5000 5.1000 ;
	    RECT 51.0000 1.1000 51.4000 4.8000 ;
	    RECT 53.4000 1.1000 53.8000 4.8000 ;
	    RECT 54.1000 4.7000 54.5000 4.8000 ;
	    RECT 55.6000 4.8000 56.6000 5.1000 ;
	    RECT 57.4000 4.8000 58.6000 5.1000 ;
	    RECT 55.6000 1.1000 56.4000 4.8000 ;
	    RECT 57.4000 4.7000 57.8000 4.8000 ;
	    RECT 58.2000 1.1000 58.6000 4.8000 ;
	    RECT 61.4000 4.7000 62.3000 5.1000 ;
	    RECT 61.9000 1.1000 62.3000 4.7000 ;
	    RECT 63.0000 1.1000 63.4000 5.8000 ;
	    RECT 67.0000 6.2000 67.3000 6.8000 ;
	    RECT 67.6000 6.8000 69.8000 7.0000 ;
	    RECT 70.2000 7.1000 71.0000 7.2000 ;
	    RECT 72.9000 7.1000 73.2000 8.1000 ;
	    RECT 75.0000 7.9000 75.4000 9.9000 ;
	    RECT 73.5000 7.4000 73.9000 7.8000 ;
	    RECT 74.2000 7.6000 75.4000 7.9000 ;
	    RECT 76.6000 8.9000 77.0000 9.9000 ;
	    RECT 74.2000 7.5000 74.6000 7.6000 ;
	    RECT 70.2000 7.0000 71.3000 7.1000 ;
	    RECT 70.2000 6.8000 72.4000 7.0000 ;
	    RECT 67.6000 6.7000 69.0000 6.8000 ;
	    RECT 67.6000 6.6000 68.0000 6.7000 ;
	    RECT 69.4000 6.2000 69.7000 6.8000 ;
	    RECT 71.0000 6.7000 72.4000 6.8000 ;
	    RECT 72.0000 6.6000 72.4000 6.7000 ;
	    RECT 72.7000 6.8000 73.2000 7.1000 ;
	    RECT 73.6000 7.2000 73.9000 7.4000 ;
	    RECT 76.6000 7.2000 76.9000 8.9000 ;
	    RECT 77.4000 7.8000 77.8000 8.6000 ;
	    RECT 78.2000 7.8000 78.6000 8.6000 ;
	    RECT 73.6000 6.8000 74.0000 7.2000 ;
	    RECT 74.6000 6.8000 75.4000 7.2000 ;
	    RECT 76.6000 7.1000 77.0000 7.2000 ;
	    RECT 79.0000 7.1000 79.4000 9.9000 ;
	    RECT 79.8000 8.0000 80.2000 9.9000 ;
	    RECT 81.4000 9.6000 83.4000 9.9000 ;
	    RECT 81.4000 8.0000 81.8000 9.6000 ;
	    RECT 79.8000 7.9000 81.8000 8.0000 ;
	    RECT 82.2000 7.9000 82.6000 9.3000 ;
	    RECT 83.0000 7.9000 83.4000 9.6000 ;
	    RECT 85.3000 7.9000 86.1000 9.9000 ;
	    RECT 79.9000 7.7000 81.7000 7.9000 ;
	    RECT 80.2000 7.2000 80.6000 7.4000 ;
	    RECT 82.3000 7.2000 82.6000 7.9000 ;
	    RECT 79.8000 7.1000 80.6000 7.2000 ;
	    RECT 76.6000 6.8000 78.5000 7.1000 ;
	    RECT 72.7000 6.2000 73.0000 6.8000 ;
	    RECT 67.0000 5.8000 67.4000 6.2000 ;
	    RECT 68.3000 6.1000 68.7000 6.2000 ;
	    RECT 67.9000 5.8000 68.7000 6.1000 ;
	    RECT 69.4000 5.8000 69.8000 6.2000 ;
	    RECT 71.3000 6.1000 71.7000 6.2000 ;
	    RECT 72.6000 6.1000 73.0000 6.2000 ;
	    RECT 75.8000 6.1000 76.2000 6.2000 ;
	    RECT 71.3000 5.8000 72.1000 6.1000 ;
	    RECT 72.6000 5.8000 76.2000 6.1000 ;
	    RECT 67.0000 5.1000 67.3000 5.8000 ;
	    RECT 67.9000 5.7000 68.3000 5.8000 ;
	    RECT 71.7000 5.7000 72.1000 5.8000 ;
	    RECT 72.7000 5.1000 73.0000 5.8000 ;
	    RECT 75.8000 5.4000 76.2000 5.8000 ;
	    RECT 76.6000 5.1000 76.9000 6.8000 ;
	    RECT 78.2000 6.2000 78.5000 6.8000 ;
	    RECT 79.0000 6.9000 80.6000 7.1000 ;
	    RECT 81.4000 6.9000 82.6000 7.2000 ;
	    RECT 79.0000 6.8000 80.2000 6.9000 ;
	    RECT 81.4000 6.8000 81.8000 6.9000 ;
	    RECT 78.2000 5.8000 78.6000 6.2000 ;
	    RECT 64.6000 4.8000 65.8000 5.1000 ;
	    RECT 64.6000 1.1000 65.0000 4.8000 ;
	    RECT 65.4000 4.7000 65.8000 4.8000 ;
	    RECT 66.8000 1.1000 67.6000 5.1000 ;
	    RECT 68.5000 4.8000 69.8000 5.1000 ;
	    RECT 68.5000 4.7000 68.9000 4.8000 ;
	    RECT 69.4000 1.1000 69.8000 4.8000 ;
	    RECT 70.2000 4.8000 71.5000 5.1000 ;
	    RECT 70.2000 1.1000 70.6000 4.8000 ;
	    RECT 71.1000 4.7000 71.5000 4.8000 ;
	    RECT 72.4000 1.1000 73.2000 5.1000 ;
	    RECT 74.2000 4.8000 75.4000 5.1000 ;
	    RECT 74.2000 4.7000 74.6000 4.8000 ;
	    RECT 75.0000 1.1000 75.4000 4.8000 ;
	    RECT 76.1000 4.7000 77.0000 5.1000 ;
	    RECT 76.1000 1.1000 76.5000 4.7000 ;
	    RECT 79.0000 1.1000 79.4000 6.8000 ;
	    RECT 80.6000 5.8000 81.0000 6.6000 ;
	    RECT 81.4000 5.1000 81.7000 6.8000 ;
	    RECT 82.2000 5.8000 82.6000 6.6000 ;
	    RECT 83.0000 6.4000 83.4000 7.2000 ;
	    RECT 84.6000 6.4000 85.0000 7.2000 ;
	    RECT 85.5000 6.2000 85.8000 7.9000 ;
	    RECT 86.2000 6.8000 86.6000 7.2000 ;
	    RECT 86.2000 6.6000 86.5000 6.8000 ;
	    RECT 86.1000 6.2000 86.5000 6.6000 ;
	    RECT 83.8000 6.1000 84.2000 6.2000 ;
	    RECT 83.8000 5.8000 84.6000 6.1000 ;
	    RECT 85.4000 5.8000 85.8000 6.2000 ;
	    RECT 84.2000 5.6000 84.6000 5.8000 ;
	    RECT 85.5000 5.7000 85.8000 5.8000 ;
	    RECT 87.0000 6.1000 87.4000 6.2000 ;
	    RECT 87.8000 6.1000 88.2000 9.9000 ;
	    RECT 89.7000 9.2000 90.1000 9.9000 ;
	    RECT 93.1000 9.2000 93.5000 9.9000 ;
	    RECT 89.4000 8.8000 90.1000 9.2000 ;
	    RECT 92.6000 8.8000 93.5000 9.2000 ;
	    RECT 88.6000 7.8000 89.0000 8.6000 ;
	    RECT 89.7000 8.2000 90.1000 8.8000 ;
	    RECT 93.1000 8.2000 93.5000 8.8000 ;
	    RECT 89.7000 7.9000 90.6000 8.2000 ;
	    RECT 87.0000 5.8000 88.2000 6.1000 ;
	    RECT 85.5000 5.4000 86.5000 5.7000 ;
	    RECT 87.0000 5.4000 87.4000 5.8000 ;
	    RECT 86.2000 5.2000 86.5000 5.4000 ;
	    RECT 81.1000 1.1000 82.1000 5.1000 ;
	    RECT 83.8000 4.8000 85.8000 5.1000 ;
	    RECT 83.8000 1.1000 84.2000 4.8000 ;
	    RECT 85.4000 1.4000 85.8000 4.8000 ;
	    RECT 86.2000 1.7000 86.6000 5.2000 ;
	    RECT 87.0000 1.4000 87.4000 5.1000 ;
	    RECT 85.4000 1.1000 87.4000 1.4000 ;
	    RECT 87.8000 1.1000 88.2000 5.8000 ;
	    RECT 89.4000 4.4000 89.8000 5.2000 ;
	    RECT 90.2000 1.1000 90.6000 7.9000 ;
	    RECT 92.6000 7.9000 93.5000 8.2000 ;
	    RECT 94.2000 7.9000 94.6000 9.9000 ;
	    RECT 96.3000 8.4000 96.7000 9.9000 ;
	    RECT 96.3000 7.9000 97.0000 8.4000 ;
	    RECT 97.5000 8.2000 97.9000 8.6000 ;
	    RECT 91.0000 6.8000 91.4000 7.6000 ;
	    RECT 91.8000 6.8000 92.2000 7.6000 ;
	    RECT 92.6000 1.1000 93.0000 7.9000 ;
	    RECT 94.3000 7.8000 94.6000 7.9000 ;
	    RECT 94.3000 7.6000 95.2000 7.8000 ;
	    RECT 94.3000 7.5000 96.4000 7.6000 ;
	    RECT 94.9000 7.3000 96.4000 7.5000 ;
	    RECT 96.0000 7.2000 96.4000 7.3000 ;
	    RECT 94.2000 6.4000 94.6000 7.2000 ;
	    RECT 95.2000 6.9000 95.6000 7.0000 ;
	    RECT 95.1000 6.6000 95.6000 6.9000 ;
	    RECT 95.1000 6.2000 95.4000 6.6000 ;
	    RECT 95.0000 5.8000 95.4000 6.2000 ;
	    RECT 96.0000 5.5000 96.3000 7.2000 ;
	    RECT 96.7000 6.2000 97.0000 7.9000 ;
	    RECT 97.4000 7.8000 97.8000 8.2000 ;
	    RECT 98.2000 7.9000 98.6000 9.9000 ;
	    RECT 101.4000 8.9000 101.8000 9.9000 ;
	    RECT 101.4000 8.1000 101.7000 8.9000 ;
	    RECT 96.6000 5.8000 97.0000 6.2000 ;
	    RECT 97.4000 6.1000 97.8000 6.2000 ;
	    RECT 98.3000 6.1000 98.6000 7.9000 ;
	    RECT 100.6000 7.8000 101.7000 8.1000 ;
	    RECT 102.2000 7.8000 102.6000 8.6000 ;
	    RECT 103.3000 8.2000 103.7000 9.9000 ;
	    RECT 106.2000 8.9000 106.6000 9.9000 ;
	    RECT 103.3000 7.9000 104.2000 8.2000 ;
	    RECT 100.6000 7.2000 100.9000 7.8000 ;
	    RECT 101.4000 7.2000 101.7000 7.8000 ;
	    RECT 99.0000 6.4000 99.4000 7.2000 ;
	    RECT 100.6000 6.8000 101.0000 7.2000 ;
	    RECT 101.4000 6.8000 101.8000 7.2000 ;
	    RECT 103.0000 7.1000 103.4000 7.2000 ;
	    RECT 103.8000 7.1000 104.2000 7.9000 ;
	    RECT 105.4000 7.8000 105.8000 8.6000 ;
	    RECT 103.0000 6.8000 104.2000 7.1000 ;
	    RECT 104.6000 6.8000 105.0000 7.6000 ;
	    RECT 106.3000 7.2000 106.6000 8.9000 ;
	    RECT 106.2000 7.1000 106.6000 7.2000 ;
	    RECT 105.4000 6.8000 106.6000 7.1000 ;
	    RECT 99.8000 6.1000 100.2000 6.2000 ;
	    RECT 97.4000 5.8000 98.6000 6.1000 ;
	    RECT 99.4000 5.8000 100.2000 6.1000 ;
	    RECT 95.1000 5.2000 96.3000 5.5000 ;
	    RECT 93.4000 4.4000 93.8000 5.2000 ;
	    RECT 95.1000 3.1000 95.4000 5.2000 ;
	    RECT 96.7000 5.1000 97.0000 5.8000 ;
	    RECT 97.5000 5.1000 97.8000 5.8000 ;
	    RECT 99.4000 5.6000 99.8000 5.8000 ;
	    RECT 100.6000 5.4000 101.0000 6.2000 ;
	    RECT 101.4000 5.1000 101.7000 6.8000 ;
	    RECT 95.0000 1.1000 95.4000 3.1000 ;
	    RECT 96.6000 1.1000 97.0000 5.1000 ;
	    RECT 97.4000 1.1000 97.8000 5.1000 ;
	    RECT 98.2000 4.8000 100.2000 5.1000 ;
	    RECT 98.2000 1.1000 98.6000 4.8000 ;
	    RECT 99.8000 1.1000 100.2000 4.8000 ;
	    RECT 100.9000 4.7000 101.8000 5.1000 ;
	    RECT 100.9000 1.1000 101.3000 4.7000 ;
	    RECT 103.0000 4.4000 103.4000 5.2000 ;
	    RECT 103.8000 1.1000 104.2000 6.8000 ;
	    RECT 105.4000 6.2000 105.7000 6.8000 ;
	    RECT 105.4000 5.8000 105.8000 6.2000 ;
	    RECT 106.3000 5.1000 106.6000 6.8000 ;
	    RECT 107.0000 6.1000 107.4000 6.2000 ;
	    RECT 107.8000 6.1000 108.2000 9.9000 ;
	    RECT 108.6000 8.1000 109.0000 8.6000 ;
	    RECT 110.2000 8.1000 110.6000 8.2000 ;
	    RECT 108.6000 7.8000 110.6000 8.1000 ;
	    RECT 111.0000 7.9000 111.4000 9.9000 ;
	    RECT 113.2000 8.1000 114.0000 9.9000 ;
	    RECT 111.0000 7.6000 112.2000 7.9000 ;
	    RECT 111.8000 7.5000 112.2000 7.6000 ;
	    RECT 112.5000 7.4000 112.9000 7.8000 ;
	    RECT 112.5000 7.2000 112.8000 7.4000 ;
	    RECT 111.0000 6.8000 111.8000 7.2000 ;
	    RECT 112.4000 6.8000 112.8000 7.2000 ;
	    RECT 113.2000 6.4000 113.5000 8.1000 ;
	    RECT 115.8000 7.9000 116.2000 9.9000 ;
	    RECT 116.9000 9.2000 117.3000 9.9000 ;
	    RECT 116.9000 8.8000 117.8000 9.2000 ;
	    RECT 116.9000 8.2000 117.3000 8.8000 ;
	    RECT 116.9000 7.9000 117.8000 8.2000 ;
	    RECT 113.8000 7.7000 114.6000 7.8000 ;
	    RECT 113.8000 7.4000 114.8000 7.7000 ;
	    RECT 115.1000 7.6000 116.2000 7.9000 ;
	    RECT 115.1000 7.5000 115.5000 7.6000 ;
	    RECT 114.5000 7.2000 114.8000 7.4000 ;
	    RECT 113.8000 6.7000 114.2000 7.1000 ;
	    RECT 114.5000 6.9000 116.2000 7.2000 ;
	    RECT 115.4000 6.8000 116.2000 6.9000 ;
	    RECT 113.0000 6.2000 113.5000 6.4000 ;
	    RECT 107.0000 5.8000 108.2000 6.1000 ;
	    RECT 112.6000 6.1000 113.5000 6.2000 ;
	    RECT 113.9000 6.4000 114.2000 6.7000 ;
	    RECT 113.9000 6.1000 115.2000 6.4000 ;
	    RECT 112.6000 5.8000 113.3000 6.1000 ;
	    RECT 114.8000 6.0000 115.2000 6.1000 ;
	    RECT 107.0000 5.4000 107.4000 5.8000 ;
	    RECT 106.2000 4.7000 107.1000 5.1000 ;
	    RECT 106.7000 1.1000 107.1000 4.7000 ;
	    RECT 107.8000 1.1000 108.2000 5.8000 ;
	    RECT 113.0000 5.2000 113.3000 5.8000 ;
	    RECT 113.7000 5.7000 114.1000 5.8000 ;
	    RECT 113.7000 5.4000 115.4000 5.7000 ;
	    RECT 112.6000 5.1000 113.3000 5.2000 ;
	    RECT 115.1000 5.1000 115.4000 5.4000 ;
	    RECT 111.0000 4.8000 112.2000 5.1000 ;
	    RECT 112.6000 4.8000 114.0000 5.1000 ;
	    RECT 111.0000 1.1000 111.4000 4.8000 ;
	    RECT 111.8000 4.7000 112.2000 4.8000 ;
	    RECT 113.2000 1.1000 114.0000 4.8000 ;
	    RECT 115.1000 4.8000 116.2000 5.1000 ;
	    RECT 115.1000 4.7000 115.5000 4.8000 ;
	    RECT 115.8000 1.1000 116.2000 4.8000 ;
	    RECT 116.6000 4.4000 117.0000 5.2000 ;
	    RECT 117.4000 1.1000 117.8000 7.9000 ;
	    RECT 118.2000 6.8000 118.6000 7.6000 ;
	    RECT 118.2000 5.1000 118.6000 5.2000 ;
	    RECT 119.0000 5.1000 119.4000 9.9000 ;
	    RECT 121.4000 8.9000 121.8000 9.9000 ;
	    RECT 123.3000 9.2000 123.7000 9.9000 ;
	    RECT 119.8000 8.1000 120.2000 8.6000 ;
	    RECT 120.6000 8.1000 121.0000 8.6000 ;
	    RECT 121.5000 8.1000 121.8000 8.9000 ;
	    RECT 123.0000 8.8000 123.7000 9.2000 ;
	    RECT 123.3000 8.2000 123.7000 8.8000 ;
	    RECT 122.2000 8.1000 122.6000 8.2000 ;
	    RECT 119.8000 7.8000 121.0000 8.1000 ;
	    RECT 121.4000 7.8000 122.6000 8.1000 ;
	    RECT 123.3000 7.9000 124.2000 8.2000 ;
	    RECT 121.5000 7.2000 121.8000 7.8000 ;
	    RECT 121.4000 6.8000 121.8000 7.2000 ;
	    RECT 121.5000 5.1000 121.8000 6.8000 ;
	    RECT 122.2000 5.4000 122.6000 6.2000 ;
	    RECT 118.2000 4.8000 119.4000 5.1000 ;
	    RECT 119.0000 1.1000 119.4000 4.8000 ;
	    RECT 121.4000 4.7000 122.3000 5.1000 ;
	    RECT 121.9000 1.1000 122.3000 4.7000 ;
	    RECT 123.0000 4.4000 123.4000 5.2000 ;
	    RECT 123.8000 1.1000 124.2000 7.9000 ;
	    RECT 125.4000 7.9000 125.8000 9.9000 ;
	    RECT 127.6000 8.1000 128.4000 9.9000 ;
	    RECT 125.4000 7.6000 126.6000 7.9000 ;
	    RECT 124.6000 6.8000 125.0000 7.6000 ;
	    RECT 126.2000 7.5000 126.6000 7.6000 ;
	    RECT 126.9000 7.4000 127.3000 7.8000 ;
	    RECT 126.9000 7.2000 127.2000 7.4000 ;
	    RECT 125.4000 6.8000 126.2000 7.2000 ;
	    RECT 126.8000 6.8000 127.2000 7.2000 ;
	    RECT 127.6000 7.1000 127.9000 8.1000 ;
	    RECT 130.2000 7.9000 130.6000 9.9000 ;
	    RECT 128.2000 7.4000 129.0000 7.8000 ;
	    RECT 129.3000 7.6000 130.6000 7.9000 ;
	    RECT 132.6000 7.9000 133.0000 9.9000 ;
	    RECT 135.0000 8.9000 135.4000 9.9000 ;
	    RECT 133.3000 8.2000 133.7000 8.6000 ;
	    RECT 129.3000 7.5000 129.7000 7.6000 ;
	    RECT 129.8000 7.1000 130.6000 7.2000 ;
	    RECT 127.6000 6.8000 128.1000 7.1000 ;
	    RECT 129.5000 7.0000 130.6000 7.1000 ;
	    RECT 127.8000 6.2000 128.1000 6.8000 ;
	    RECT 128.4000 6.8000 130.6000 7.0000 ;
	    RECT 128.4000 6.7000 129.8000 6.8000 ;
	    RECT 128.4000 6.6000 128.8000 6.7000 ;
	    RECT 131.8000 6.4000 132.2000 7.2000 ;
	    RECT 127.0000 5.8000 127.4000 6.2000 ;
	    RECT 127.8000 5.8000 128.2000 6.2000 ;
	    RECT 129.1000 6.1000 129.5000 6.2000 ;
	    RECT 128.7000 5.8000 129.5000 6.1000 ;
	    RECT 131.0000 6.1000 131.4000 6.2000 ;
	    RECT 132.6000 6.1000 132.9000 7.9000 ;
	    RECT 133.4000 7.8000 133.8000 8.2000 ;
	    RECT 134.2000 7.8000 134.6000 8.6000 ;
	    RECT 133.4000 7.1000 133.7000 7.8000 ;
	    RECT 135.1000 7.2000 135.4000 8.9000 ;
	    RECT 137.9000 8.2000 138.3000 9.9000 ;
	    RECT 137.4000 7.9000 138.3000 8.2000 ;
	    RECT 135.0000 7.1000 135.4000 7.2000 ;
	    RECT 133.4000 6.8000 135.4000 7.1000 ;
	    RECT 136.6000 6.8000 137.0000 7.6000 ;
	    RECT 137.4000 7.1000 137.8000 7.9000 ;
	    RECT 138.2000 7.1000 138.6000 7.2000 ;
	    RECT 137.4000 6.8000 138.6000 7.1000 ;
	    RECT 133.4000 6.1000 133.8000 6.2000 ;
	    RECT 131.0000 5.8000 131.8000 6.1000 ;
	    RECT 132.6000 5.8000 133.8000 6.1000 ;
	    RECT 127.0000 5.2000 127.3000 5.8000 ;
	    RECT 127.8000 5.2000 128.1000 5.8000 ;
	    RECT 128.7000 5.7000 129.1000 5.8000 ;
	    RECT 131.4000 5.6000 131.8000 5.8000 ;
	    RECT 127.0000 5.1000 128.1000 5.2000 ;
	    RECT 133.4000 5.1000 133.7000 5.8000 ;
	    RECT 135.1000 5.1000 135.4000 6.8000 ;
	    RECT 135.8000 5.4000 136.2000 6.2000 ;
	    RECT 125.4000 4.8000 126.6000 5.1000 ;
	    RECT 127.0000 4.8000 128.4000 5.1000 ;
	    RECT 125.4000 1.1000 125.8000 4.8000 ;
	    RECT 126.2000 4.7000 126.6000 4.8000 ;
	    RECT 127.6000 1.1000 128.4000 4.8000 ;
	    RECT 129.3000 4.8000 130.6000 5.1000 ;
	    RECT 129.3000 4.7000 129.7000 4.8000 ;
	    RECT 130.2000 1.1000 130.6000 4.8000 ;
	    RECT 131.0000 4.8000 133.0000 5.1000 ;
	    RECT 131.0000 1.1000 131.4000 4.8000 ;
	    RECT 132.6000 1.1000 133.0000 4.8000 ;
	    RECT 133.4000 1.1000 133.8000 5.1000 ;
	    RECT 135.0000 4.7000 135.9000 5.1000 ;
	    RECT 135.5000 1.1000 135.9000 4.7000 ;
	    RECT 137.4000 1.1000 137.8000 6.8000 ;
	    RECT 138.2000 5.8000 138.6000 6.2000 ;
	    RECT 138.2000 5.2000 138.5000 5.8000 ;
	    RECT 138.2000 5.1000 138.6000 5.2000 ;
	    RECT 139.0000 5.1000 139.4000 9.9000 ;
	    RECT 140.9000 9.2000 141.3000 9.9000 ;
	    RECT 140.9000 8.8000 141.8000 9.2000 ;
	    RECT 139.8000 7.8000 140.2000 8.6000 ;
	    RECT 140.9000 8.2000 141.3000 8.8000 ;
	    RECT 140.9000 7.9000 141.8000 8.2000 ;
	    RECT 138.2000 4.8000 139.4000 5.1000 ;
	    RECT 138.2000 4.4000 138.6000 4.8000 ;
	    RECT 139.0000 1.1000 139.4000 4.8000 ;
	    RECT 140.6000 4.4000 141.0000 5.2000 ;
	    RECT 141.4000 1.1000 141.8000 7.9000 ;
	    RECT 143.0000 7.7000 143.4000 9.9000 ;
	    RECT 145.1000 9.2000 145.7000 9.9000 ;
	    RECT 145.1000 8.9000 145.8000 9.2000 ;
	    RECT 147.4000 8.9000 147.8000 9.9000 ;
	    RECT 149.6000 9.2000 150.0000 9.9000 ;
	    RECT 149.6000 8.9000 150.6000 9.2000 ;
	    RECT 145.4000 8.5000 145.8000 8.9000 ;
	    RECT 147.5000 8.6000 147.8000 8.9000 ;
	    RECT 147.5000 8.3000 148.9000 8.6000 ;
	    RECT 148.5000 8.2000 148.9000 8.3000 ;
	    RECT 149.4000 8.2000 149.8000 8.6000 ;
	    RECT 150.2000 8.5000 150.6000 8.9000 ;
	    RECT 144.5000 7.7000 144.9000 7.8000 ;
	    RECT 142.2000 6.8000 142.6000 7.6000 ;
	    RECT 143.0000 7.4000 144.9000 7.7000 ;
	    RECT 143.0000 5.7000 143.4000 7.4000 ;
	    RECT 146.5000 7.1000 146.9000 7.2000 ;
	    RECT 149.4000 7.1000 149.7000 8.2000 ;
	    RECT 151.8000 7.5000 152.2000 9.9000 ;
	    RECT 152.6000 7.9000 153.0000 9.9000 ;
	    RECT 154.8000 8.1000 155.6000 9.9000 ;
	    RECT 152.6000 7.6000 153.8000 7.9000 ;
	    RECT 153.4000 7.5000 153.8000 7.6000 ;
	    RECT 154.1000 7.4000 154.5000 7.8000 ;
	    RECT 154.1000 7.2000 154.4000 7.4000 ;
	    RECT 151.0000 7.1000 151.8000 7.2000 ;
	    RECT 146.3000 6.8000 151.8000 7.1000 ;
	    RECT 152.6000 6.8000 153.4000 7.2000 ;
	    RECT 154.0000 6.8000 154.4000 7.2000 ;
	    RECT 145.4000 6.4000 145.8000 6.5000 ;
	    RECT 143.9000 6.1000 145.8000 6.4000 ;
	    RECT 143.9000 6.0000 144.3000 6.1000 ;
	    RECT 144.7000 5.7000 145.1000 5.8000 ;
	    RECT 143.0000 5.4000 145.1000 5.7000 ;
	    RECT 143.0000 1.1000 143.4000 5.4000 ;
	    RECT 146.3000 5.2000 146.6000 6.8000 ;
	    RECT 149.9000 6.7000 150.3000 6.8000 ;
	    RECT 154.8000 6.4000 155.1000 8.1000 ;
	    RECT 157.4000 7.9000 157.8000 9.9000 ;
	    RECT 158.2000 9.1000 158.6000 9.2000 ;
	    RECT 159.8000 9.1000 160.2000 9.9000 ;
	    RECT 158.2000 8.8000 160.2000 9.1000 ;
	    RECT 161.9000 9.2000 162.5000 9.9000 ;
	    RECT 161.9000 8.9000 162.6000 9.2000 ;
	    RECT 164.2000 8.9000 164.6000 9.9000 ;
	    RECT 166.4000 9.2000 166.8000 9.9000 ;
	    RECT 166.4000 8.9000 167.4000 9.2000 ;
	    RECT 155.4000 7.7000 156.2000 7.8000 ;
	    RECT 155.4000 7.4000 156.4000 7.7000 ;
	    RECT 156.7000 7.6000 157.8000 7.9000 ;
	    RECT 159.8000 7.7000 160.2000 8.8000 ;
	    RECT 162.2000 8.5000 162.6000 8.9000 ;
	    RECT 164.3000 8.6000 164.6000 8.9000 ;
	    RECT 164.3000 8.3000 165.7000 8.6000 ;
	    RECT 165.3000 8.2000 165.7000 8.3000 ;
	    RECT 166.2000 8.2000 166.6000 8.6000 ;
	    RECT 167.0000 8.5000 167.4000 8.9000 ;
	    RECT 161.3000 7.7000 161.7000 7.8000 ;
	    RECT 156.7000 7.5000 157.1000 7.6000 ;
	    RECT 156.1000 7.2000 156.4000 7.4000 ;
	    RECT 159.8000 7.4000 161.7000 7.7000 ;
	    RECT 156.1000 7.1000 157.8000 7.2000 ;
	    RECT 159.8000 7.1000 160.2000 7.4000 ;
	    RECT 163.3000 7.1000 163.7000 7.2000 ;
	    RECT 164.6000 7.1000 165.0000 7.2000 ;
	    RECT 166.2000 7.1000 166.5000 8.2000 ;
	    RECT 168.6000 7.5000 169.0000 9.9000 ;
	    RECT 170.2000 8.9000 170.6000 9.9000 ;
	    RECT 169.4000 7.8000 169.8000 8.6000 ;
	    RECT 170.3000 7.8000 170.6000 8.9000 ;
	    RECT 171.8000 7.9000 172.2000 9.9000 ;
	    RECT 170.3000 7.5000 171.5000 7.8000 ;
	    RECT 167.8000 7.1000 168.6000 7.2000 ;
	    RECT 155.4000 6.7000 155.8000 7.1000 ;
	    RECT 156.1000 6.9000 160.2000 7.1000 ;
	    RECT 157.0000 6.8000 160.2000 6.9000 ;
	    RECT 150.7000 6.2000 151.1000 6.3000 ;
	    RECT 154.6000 6.2000 155.1000 6.4000 ;
	    RECT 147.0000 6.1000 147.4000 6.2000 ;
	    RECT 148.6000 6.1000 151.1000 6.2000 ;
	    RECT 147.0000 5.9000 151.1000 6.1000 ;
	    RECT 154.2000 6.1000 155.1000 6.2000 ;
	    RECT 155.5000 6.4000 155.8000 6.7000 ;
	    RECT 155.5000 6.1000 156.8000 6.4000 ;
	    RECT 147.0000 5.8000 149.0000 5.9000 ;
	    RECT 154.2000 5.8000 154.9000 6.1000 ;
	    RECT 156.4000 6.0000 156.8000 6.1000 ;
	    RECT 149.4000 5.5000 152.2000 5.6000 ;
	    RECT 149.3000 5.4000 152.2000 5.5000 ;
	    RECT 145.4000 4.9000 146.6000 5.2000 ;
	    RECT 147.3000 5.3000 152.2000 5.4000 ;
	    RECT 147.3000 5.1000 149.7000 5.3000 ;
	    RECT 145.4000 4.4000 145.7000 4.9000 ;
	    RECT 145.0000 4.0000 145.7000 4.4000 ;
	    RECT 146.5000 4.5000 146.9000 4.6000 ;
	    RECT 147.3000 4.5000 147.6000 5.1000 ;
	    RECT 146.5000 4.2000 147.6000 4.5000 ;
	    RECT 147.9000 4.5000 150.6000 4.8000 ;
	    RECT 147.9000 4.4000 148.3000 4.5000 ;
	    RECT 150.2000 4.4000 150.6000 4.5000 ;
	    RECT 147.1000 3.7000 147.5000 3.8000 ;
	    RECT 148.5000 3.7000 148.9000 3.8000 ;
	    RECT 145.4000 3.1000 145.8000 3.5000 ;
	    RECT 147.1000 3.4000 148.9000 3.7000 ;
	    RECT 147.5000 3.1000 147.8000 3.4000 ;
	    RECT 150.2000 3.1000 150.6000 3.5000 ;
	    RECT 145.1000 1.1000 145.7000 3.1000 ;
	    RECT 147.4000 1.1000 147.8000 3.1000 ;
	    RECT 149.6000 2.8000 150.6000 3.1000 ;
	    RECT 149.6000 1.1000 150.0000 2.8000 ;
	    RECT 151.8000 1.1000 152.2000 5.3000 ;
	    RECT 154.6000 5.2000 154.9000 5.8000 ;
	    RECT 155.3000 5.7000 155.7000 5.8000 ;
	    RECT 159.8000 5.7000 160.2000 6.8000 ;
	    RECT 163.1000 6.8000 168.6000 7.1000 ;
	    RECT 170.2000 6.8000 170.7000 7.2000 ;
	    RECT 162.2000 6.4000 162.6000 6.5000 ;
	    RECT 160.7000 6.1000 162.6000 6.4000 ;
	    RECT 160.7000 6.0000 161.1000 6.1000 ;
	    RECT 161.5000 5.7000 161.9000 5.8000 ;
	    RECT 155.3000 5.4000 157.0000 5.7000 ;
	    RECT 154.2000 5.1000 154.9000 5.2000 ;
	    RECT 156.7000 5.1000 157.0000 5.4000 ;
	    RECT 159.8000 5.4000 161.9000 5.7000 ;
	    RECT 152.6000 4.8000 153.8000 5.1000 ;
	    RECT 154.2000 4.8000 155.6000 5.1000 ;
	    RECT 152.6000 1.1000 153.0000 4.8000 ;
	    RECT 153.4000 4.7000 153.8000 4.8000 ;
	    RECT 154.8000 1.1000 155.6000 4.8000 ;
	    RECT 156.7000 4.8000 157.8000 5.1000 ;
	    RECT 156.7000 4.7000 157.1000 4.8000 ;
	    RECT 157.4000 1.1000 157.8000 4.8000 ;
	    RECT 159.8000 1.1000 160.2000 5.4000 ;
	    RECT 163.1000 5.2000 163.4000 6.8000 ;
	    RECT 166.7000 6.7000 167.1000 6.8000 ;
	    RECT 170.4000 6.4000 170.8000 6.8000 ;
	    RECT 167.5000 6.2000 167.9000 6.3000 ;
	    RECT 163.8000 6.1000 164.2000 6.2000 ;
	    RECT 165.4000 6.1000 167.9000 6.2000 ;
	    RECT 163.8000 5.9000 167.9000 6.1000 ;
	    RECT 171.2000 6.0000 171.5000 7.5000 ;
	    RECT 171.9000 6.2000 172.2000 7.9000 ;
	    RECT 163.8000 5.8000 165.8000 5.9000 ;
	    RECT 171.1000 5.7000 171.5000 6.0000 ;
	    RECT 171.8000 5.8000 172.2000 6.2000 ;
	    RECT 169.4000 5.6000 171.5000 5.7000 ;
	    RECT 166.2000 5.5000 169.0000 5.6000 ;
	    RECT 166.1000 5.4000 169.0000 5.5000 ;
	    RECT 162.2000 4.9000 163.4000 5.2000 ;
	    RECT 164.1000 5.3000 169.0000 5.4000 ;
	    RECT 164.1000 5.1000 166.5000 5.3000 ;
	    RECT 162.2000 4.4000 162.5000 4.9000 ;
	    RECT 161.8000 4.0000 162.5000 4.4000 ;
	    RECT 163.3000 4.5000 163.7000 4.6000 ;
	    RECT 164.1000 4.5000 164.4000 5.1000 ;
	    RECT 163.3000 4.2000 164.4000 4.5000 ;
	    RECT 164.7000 4.5000 167.4000 4.8000 ;
	    RECT 164.7000 4.4000 165.1000 4.5000 ;
	    RECT 167.0000 4.4000 167.4000 4.5000 ;
	    RECT 163.9000 3.7000 164.3000 3.8000 ;
	    RECT 165.3000 3.7000 165.7000 3.8000 ;
	    RECT 162.2000 3.1000 162.6000 3.5000 ;
	    RECT 163.9000 3.4000 165.7000 3.7000 ;
	    RECT 164.3000 3.1000 164.6000 3.4000 ;
	    RECT 167.0000 3.1000 167.4000 3.5000 ;
	    RECT 161.9000 1.1000 162.5000 3.1000 ;
	    RECT 164.2000 1.1000 164.6000 3.1000 ;
	    RECT 166.4000 2.8000 167.4000 3.1000 ;
	    RECT 166.4000 1.1000 166.8000 2.8000 ;
	    RECT 168.6000 1.1000 169.0000 5.3000 ;
	    RECT 169.4000 5.4000 171.4000 5.6000 ;
	    RECT 169.4000 1.1000 169.8000 5.4000 ;
	    RECT 171.9000 5.1000 172.2000 5.8000 ;
	    RECT 171.5000 4.8000 172.2000 5.1000 ;
	    RECT 172.6000 7.7000 173.0000 9.9000 ;
	    RECT 174.7000 9.2000 175.3000 9.9000 ;
	    RECT 174.7000 8.9000 175.4000 9.2000 ;
	    RECT 177.0000 8.9000 177.4000 9.9000 ;
	    RECT 179.2000 9.2000 179.6000 9.9000 ;
	    RECT 179.2000 8.9000 180.2000 9.2000 ;
	    RECT 175.0000 8.5000 175.4000 8.9000 ;
	    RECT 177.1000 8.6000 177.4000 8.9000 ;
	    RECT 177.1000 8.3000 178.5000 8.6000 ;
	    RECT 178.1000 8.2000 178.5000 8.3000 ;
	    RECT 179.0000 8.2000 179.4000 8.6000 ;
	    RECT 179.8000 8.5000 180.2000 8.9000 ;
	    RECT 174.1000 7.7000 174.5000 7.8000 ;
	    RECT 172.6000 7.4000 174.5000 7.7000 ;
	    RECT 172.6000 5.7000 173.0000 7.4000 ;
	    RECT 176.1000 7.1000 176.5000 7.2000 ;
	    RECT 179.0000 7.1000 179.3000 8.2000 ;
	    RECT 181.4000 7.5000 181.8000 9.9000 ;
	    RECT 183.8000 7.6000 184.2000 9.9000 ;
	    RECT 183.1000 7.3000 184.2000 7.6000 ;
	    RECT 184.6000 7.7000 185.0000 9.9000 ;
	    RECT 186.7000 9.2000 187.3000 9.9000 ;
	    RECT 186.7000 8.9000 187.4000 9.2000 ;
	    RECT 189.0000 8.9000 189.4000 9.9000 ;
	    RECT 191.2000 9.2000 191.6000 9.9000 ;
	    RECT 191.2000 8.9000 192.2000 9.2000 ;
	    RECT 187.0000 8.5000 187.4000 8.9000 ;
	    RECT 189.1000 8.6000 189.4000 8.9000 ;
	    RECT 189.1000 8.3000 190.5000 8.6000 ;
	    RECT 190.1000 8.2000 190.5000 8.3000 ;
	    RECT 191.0000 7.8000 191.4000 8.6000 ;
	    RECT 191.8000 8.5000 192.2000 8.9000 ;
	    RECT 186.1000 7.7000 186.5000 7.8000 ;
	    RECT 184.6000 7.4000 186.5000 7.7000 ;
	    RECT 180.6000 7.1000 181.4000 7.2000 ;
	    RECT 175.9000 6.8000 181.4000 7.1000 ;
	    RECT 175.0000 6.4000 175.4000 6.5000 ;
	    RECT 173.5000 6.1000 175.4000 6.4000 ;
	    RECT 175.9000 6.2000 176.2000 6.8000 ;
	    RECT 179.5000 6.7000 179.9000 6.8000 ;
	    RECT 180.3000 6.2000 180.7000 6.3000 ;
	    RECT 173.5000 6.0000 173.9000 6.1000 ;
	    RECT 175.8000 5.8000 176.2000 6.2000 ;
	    RECT 178.2000 5.9000 180.7000 6.2000 ;
	    RECT 178.2000 5.8000 178.6000 5.9000 ;
	    RECT 183.1000 5.8000 183.4000 7.3000 ;
	    RECT 183.8000 6.1000 184.2000 6.6000 ;
	    RECT 184.6000 6.1000 185.0000 7.4000 ;
	    RECT 188.1000 7.1000 188.5000 7.2000 ;
	    RECT 191.0000 7.1000 191.3000 7.8000 ;
	    RECT 193.4000 7.5000 193.8000 9.9000 ;
	    RECT 194.2000 7.8000 194.6000 8.6000 ;
	    RECT 195.0000 8.1000 195.4000 9.9000 ;
	    RECT 196.6000 8.9000 197.0000 9.9000 ;
	    RECT 195.8000 8.1000 196.2000 8.6000 ;
	    RECT 195.0000 7.8000 196.2000 8.1000 ;
	    RECT 194.2000 7.2000 194.5000 7.8000 ;
	    RECT 192.6000 7.1000 193.4000 7.2000 ;
	    RECT 187.9000 6.8000 193.4000 7.1000 ;
	    RECT 194.2000 6.8000 194.6000 7.2000 ;
	    RECT 187.0000 6.4000 187.4000 6.5000 ;
	    RECT 183.8000 5.8000 185.0000 6.1000 ;
	    RECT 185.5000 6.1000 187.4000 6.4000 ;
	    RECT 185.5000 6.0000 185.9000 6.1000 ;
	    RECT 174.3000 5.7000 174.7000 5.8000 ;
	    RECT 172.6000 5.4000 174.7000 5.7000 ;
	    RECT 171.5000 1.1000 171.9000 4.8000 ;
	    RECT 172.6000 1.1000 173.0000 5.4000 ;
	    RECT 175.9000 5.2000 176.2000 5.8000 ;
	    RECT 179.0000 5.5000 181.8000 5.6000 ;
	    RECT 178.9000 5.4000 181.8000 5.5000 ;
	    RECT 182.8000 5.4000 183.4000 5.8000 ;
	    RECT 175.0000 4.9000 176.2000 5.2000 ;
	    RECT 176.9000 5.3000 181.8000 5.4000 ;
	    RECT 176.9000 5.1000 179.3000 5.3000 ;
	    RECT 175.0000 4.4000 175.3000 4.9000 ;
	    RECT 174.6000 4.0000 175.3000 4.4000 ;
	    RECT 176.1000 4.5000 176.5000 4.6000 ;
	    RECT 176.9000 4.5000 177.2000 5.1000 ;
	    RECT 176.1000 4.2000 177.2000 4.5000 ;
	    RECT 177.5000 4.5000 180.2000 4.8000 ;
	    RECT 177.5000 4.4000 177.9000 4.5000 ;
	    RECT 179.8000 4.4000 180.2000 4.5000 ;
	    RECT 176.7000 3.7000 177.1000 3.8000 ;
	    RECT 178.1000 3.7000 178.5000 3.8000 ;
	    RECT 175.0000 3.1000 175.4000 3.5000 ;
	    RECT 176.7000 3.4000 178.5000 3.7000 ;
	    RECT 177.1000 3.1000 177.4000 3.4000 ;
	    RECT 179.8000 3.1000 180.2000 3.5000 ;
	    RECT 174.7000 1.1000 175.3000 3.1000 ;
	    RECT 177.0000 1.1000 177.4000 3.1000 ;
	    RECT 179.2000 2.8000 180.2000 3.1000 ;
	    RECT 179.2000 1.1000 179.6000 2.8000 ;
	    RECT 181.4000 1.1000 181.8000 5.3000 ;
	    RECT 183.1000 5.1000 183.4000 5.4000 ;
	    RECT 184.6000 5.7000 185.0000 5.8000 ;
	    RECT 186.3000 5.7000 186.7000 5.8000 ;
	    RECT 184.6000 5.4000 186.7000 5.7000 ;
	    RECT 183.1000 4.8000 184.2000 5.1000 ;
	    RECT 183.8000 1.1000 184.2000 4.8000 ;
	    RECT 184.6000 1.1000 185.0000 5.4000 ;
	    RECT 187.9000 5.2000 188.2000 6.8000 ;
	    RECT 191.5000 6.7000 191.9000 6.8000 ;
	    RECT 191.0000 6.2000 191.4000 6.3000 ;
	    RECT 192.3000 6.2000 192.7000 6.3000 ;
	    RECT 190.2000 5.9000 192.7000 6.2000 ;
	    RECT 190.2000 5.8000 190.6000 5.9000 ;
	    RECT 191.0000 5.5000 193.8000 5.6000 ;
	    RECT 190.9000 5.4000 193.8000 5.5000 ;
	    RECT 187.0000 4.9000 188.2000 5.2000 ;
	    RECT 188.9000 5.3000 193.8000 5.4000 ;
	    RECT 188.9000 5.1000 191.3000 5.3000 ;
	    RECT 187.0000 4.4000 187.3000 4.9000 ;
	    RECT 186.6000 4.0000 187.3000 4.4000 ;
	    RECT 188.1000 4.5000 188.5000 4.6000 ;
	    RECT 188.9000 4.5000 189.2000 5.1000 ;
	    RECT 188.1000 4.2000 189.2000 4.5000 ;
	    RECT 189.5000 4.5000 192.2000 4.8000 ;
	    RECT 189.5000 4.4000 189.9000 4.5000 ;
	    RECT 191.8000 4.4000 192.2000 4.5000 ;
	    RECT 188.7000 3.7000 189.1000 3.8000 ;
	    RECT 190.1000 3.7000 190.5000 3.8000 ;
	    RECT 187.0000 3.1000 187.4000 3.5000 ;
	    RECT 188.7000 3.4000 190.5000 3.7000 ;
	    RECT 189.1000 3.1000 189.4000 3.4000 ;
	    RECT 191.8000 3.1000 192.2000 3.5000 ;
	    RECT 186.7000 1.1000 187.3000 3.1000 ;
	    RECT 189.0000 1.1000 189.4000 3.1000 ;
	    RECT 191.2000 2.8000 192.2000 3.1000 ;
	    RECT 191.2000 1.1000 191.6000 2.8000 ;
	    RECT 193.4000 1.1000 193.8000 5.3000 ;
	    RECT 195.0000 1.1000 195.4000 7.8000 ;
	    RECT 196.7000 7.2000 197.0000 8.9000 ;
	    RECT 198.2000 7.6000 198.6000 9.9000 ;
	    RECT 201.4000 8.9000 201.8000 9.9000 ;
	    RECT 198.2000 7.3000 199.3000 7.6000 ;
	    RECT 195.8000 6.8000 196.2000 7.2000 ;
	    RECT 196.6000 6.8000 197.0000 7.2000 ;
	    RECT 195.8000 6.1000 196.1000 6.8000 ;
	    RECT 196.7000 6.1000 197.0000 6.8000 ;
	    RECT 195.8000 5.8000 197.0000 6.1000 ;
	    RECT 196.7000 5.1000 197.0000 5.8000 ;
	    RECT 197.4000 5.4000 197.8000 6.2000 ;
	    RECT 198.2000 5.8000 198.6000 6.6000 ;
	    RECT 199.0000 5.8000 199.3000 7.3000 ;
	    RECT 201.4000 7.2000 201.7000 8.9000 ;
	    RECT 202.2000 8.1000 202.6000 8.6000 ;
	    RECT 203.0000 8.1000 203.4000 9.9000 ;
	    RECT 202.2000 7.8000 203.4000 8.1000 ;
	    RECT 203.8000 7.8000 204.2000 8.6000 ;
	    RECT 201.4000 6.8000 201.8000 7.2000 ;
	    RECT 202.2000 6.8000 202.6000 7.2000 ;
	    RECT 199.0000 5.4000 199.6000 5.8000 ;
	    RECT 200.6000 5.4000 201.0000 6.2000 ;
	    RECT 201.4000 6.1000 201.7000 6.8000 ;
	    RECT 202.2000 6.1000 202.5000 6.8000 ;
	    RECT 201.4000 5.8000 202.5000 6.1000 ;
	    RECT 199.0000 5.1000 199.3000 5.4000 ;
	    RECT 201.4000 5.1000 201.7000 5.8000 ;
	    RECT 196.6000 4.7000 197.5000 5.1000 ;
	    RECT 197.1000 1.1000 197.5000 4.7000 ;
	    RECT 198.2000 4.8000 199.3000 5.1000 ;
	    RECT 198.2000 1.1000 198.6000 4.8000 ;
	    RECT 200.9000 4.7000 201.8000 5.1000 ;
	    RECT 200.9000 1.1000 201.3000 4.7000 ;
	    RECT 203.0000 1.1000 203.4000 7.8000 ;
	    RECT 204.6000 7.5000 205.0000 9.9000 ;
	    RECT 206.8000 9.2000 207.2000 9.9000 ;
	    RECT 206.2000 8.9000 207.2000 9.2000 ;
	    RECT 209.0000 8.9000 209.4000 9.9000 ;
	    RECT 211.1000 9.2000 211.7000 9.9000 ;
	    RECT 211.0000 8.9000 211.7000 9.2000 ;
	    RECT 206.2000 8.5000 206.6000 8.9000 ;
	    RECT 209.0000 8.6000 209.3000 8.9000 ;
	    RECT 207.0000 8.2000 207.4000 8.6000 ;
	    RECT 207.9000 8.3000 209.3000 8.6000 ;
	    RECT 211.0000 8.5000 211.4000 8.9000 ;
	    RECT 207.9000 8.2000 208.3000 8.3000 ;
	    RECT 205.0000 7.1000 205.8000 7.2000 ;
	    RECT 207.1000 7.1000 207.4000 8.2000 ;
	    RECT 211.9000 7.7000 212.3000 7.8000 ;
	    RECT 213.4000 7.7000 213.8000 9.9000 ;
	    RECT 214.2000 9.1000 214.6000 9.2000 ;
	    RECT 215.8000 9.1000 216.2000 9.9000 ;
	    RECT 214.2000 8.8000 216.2000 9.1000 ;
	    RECT 211.9000 7.4000 213.8000 7.7000 ;
	    RECT 209.9000 7.1000 210.3000 7.2000 ;
	    RECT 205.0000 6.8000 210.5000 7.1000 ;
	    RECT 206.5000 6.7000 206.9000 6.8000 ;
	    RECT 205.7000 6.2000 206.1000 6.3000 ;
	    RECT 207.0000 6.2000 207.4000 6.3000 ;
	    RECT 205.7000 5.9000 208.2000 6.2000 ;
	    RECT 207.8000 5.8000 208.2000 5.9000 ;
	    RECT 204.6000 5.5000 207.4000 5.6000 ;
	    RECT 204.6000 5.4000 207.5000 5.5000 ;
	    RECT 204.6000 5.3000 209.5000 5.4000 ;
	    RECT 204.6000 1.1000 205.0000 5.3000 ;
	    RECT 207.1000 5.1000 209.5000 5.3000 ;
	    RECT 206.2000 4.5000 208.9000 4.8000 ;
	    RECT 206.2000 4.4000 206.6000 4.5000 ;
	    RECT 208.5000 4.4000 208.9000 4.5000 ;
	    RECT 209.2000 4.5000 209.5000 5.1000 ;
	    RECT 210.2000 5.2000 210.5000 6.8000 ;
	    RECT 211.0000 6.4000 211.4000 6.5000 ;
	    RECT 211.0000 6.1000 212.9000 6.4000 ;
	    RECT 212.5000 6.0000 212.9000 6.1000 ;
	    RECT 211.7000 5.7000 212.1000 5.8000 ;
	    RECT 213.4000 5.7000 213.8000 7.4000 ;
	    RECT 211.7000 5.4000 213.8000 5.7000 ;
	    RECT 210.2000 4.9000 211.4000 5.2000 ;
	    RECT 209.9000 4.5000 210.3000 4.6000 ;
	    RECT 209.2000 4.2000 210.3000 4.5000 ;
	    RECT 211.1000 4.4000 211.4000 4.9000 ;
	    RECT 211.1000 4.0000 211.8000 4.4000 ;
	    RECT 207.9000 3.7000 208.3000 3.8000 ;
	    RECT 209.3000 3.7000 209.7000 3.8000 ;
	    RECT 206.2000 3.1000 206.6000 3.5000 ;
	    RECT 207.9000 3.4000 209.7000 3.7000 ;
	    RECT 209.0000 3.1000 209.3000 3.4000 ;
	    RECT 211.0000 3.1000 211.4000 3.5000 ;
	    RECT 206.2000 2.8000 207.2000 3.1000 ;
	    RECT 206.8000 1.1000 207.2000 2.8000 ;
	    RECT 209.0000 1.1000 209.4000 3.1000 ;
	    RECT 211.1000 1.1000 211.7000 3.1000 ;
	    RECT 213.4000 1.1000 213.8000 5.4000 ;
	    RECT 215.8000 6.1000 216.2000 8.8000 ;
	    RECT 217.4000 7.7000 217.8000 9.9000 ;
	    RECT 219.5000 9.2000 220.1000 9.9000 ;
	    RECT 219.5000 8.9000 220.2000 9.2000 ;
	    RECT 221.8000 8.9000 222.2000 9.9000 ;
	    RECT 224.0000 9.2000 224.4000 9.9000 ;
	    RECT 224.0000 8.9000 225.0000 9.2000 ;
	    RECT 219.8000 8.5000 220.2000 8.9000 ;
	    RECT 221.9000 8.6000 222.2000 8.9000 ;
	    RECT 221.9000 8.3000 223.3000 8.6000 ;
	    RECT 222.9000 8.2000 223.3000 8.3000 ;
	    RECT 223.8000 8.2000 224.2000 8.6000 ;
	    RECT 224.6000 8.5000 225.0000 8.9000 ;
	    RECT 218.9000 7.7000 219.3000 7.8000 ;
	    RECT 217.4000 7.4000 219.3000 7.7000 ;
	    RECT 216.6000 6.1000 217.0000 6.2000 ;
	    RECT 215.8000 5.8000 217.0000 6.1000 ;
	    RECT 215.8000 1.1000 216.2000 5.8000 ;
	    RECT 217.4000 5.7000 217.8000 7.4000 ;
	    RECT 220.9000 7.1000 221.3000 7.2000 ;
	    RECT 222.2000 7.1000 222.6000 7.2000 ;
	    RECT 223.8000 7.1000 224.1000 8.2000 ;
	    RECT 226.2000 7.5000 226.6000 9.9000 ;
	    RECT 227.0000 7.8000 227.4000 8.6000 ;
	    RECT 225.4000 7.1000 226.2000 7.2000 ;
	    RECT 220.7000 6.8000 226.2000 7.1000 ;
	    RECT 227.8000 7.1000 228.2000 9.9000 ;
	    RECT 230.5000 8.0000 230.9000 9.5000 ;
	    RECT 232.6000 8.5000 233.0000 9.5000 ;
	    RECT 230.1000 7.7000 230.9000 8.0000 ;
	    RECT 230.1000 7.5000 230.5000 7.7000 ;
	    RECT 230.1000 7.2000 230.4000 7.5000 ;
	    RECT 232.7000 7.4000 233.0000 8.5000 ;
	    RECT 233.4000 7.8000 233.8000 8.6000 ;
	    RECT 228.6000 7.1000 229.0000 7.2000 ;
	    RECT 227.8000 6.8000 229.0000 7.1000 ;
	    RECT 229.4000 6.8000 230.4000 7.2000 ;
	    RECT 230.9000 7.1000 233.0000 7.4000 ;
	    RECT 230.9000 6.9000 231.4000 7.1000 ;
	    RECT 219.8000 6.4000 220.2000 6.5000 ;
	    RECT 218.3000 6.1000 220.2000 6.4000 ;
	    RECT 218.3000 6.0000 218.7000 6.1000 ;
	    RECT 219.1000 5.7000 219.5000 5.8000 ;
	    RECT 217.4000 5.4000 219.5000 5.7000 ;
	    RECT 217.4000 1.1000 217.8000 5.4000 ;
	    RECT 220.7000 5.2000 221.0000 6.8000 ;
	    RECT 224.3000 6.7000 224.7000 6.8000 ;
	    RECT 223.8000 6.2000 224.2000 6.3000 ;
	    RECT 225.1000 6.2000 225.5000 6.3000 ;
	    RECT 223.0000 5.9000 225.5000 6.2000 ;
	    RECT 223.0000 5.8000 223.4000 5.9000 ;
	    RECT 223.8000 5.5000 226.6000 5.6000 ;
	    RECT 223.7000 5.4000 226.6000 5.5000 ;
	    RECT 219.8000 4.9000 221.0000 5.2000 ;
	    RECT 221.7000 5.3000 226.6000 5.4000 ;
	    RECT 221.7000 5.1000 224.1000 5.3000 ;
	    RECT 219.8000 4.4000 220.1000 4.9000 ;
	    RECT 219.4000 4.0000 220.1000 4.4000 ;
	    RECT 220.9000 4.5000 221.3000 4.6000 ;
	    RECT 221.7000 4.5000 222.0000 5.1000 ;
	    RECT 220.9000 4.2000 222.0000 4.5000 ;
	    RECT 222.3000 4.5000 225.0000 4.8000 ;
	    RECT 222.3000 4.4000 222.7000 4.5000 ;
	    RECT 224.6000 4.4000 225.0000 4.5000 ;
	    RECT 221.5000 3.7000 221.9000 3.8000 ;
	    RECT 222.9000 3.7000 223.3000 3.8000 ;
	    RECT 219.8000 3.1000 220.2000 3.5000 ;
	    RECT 221.5000 3.4000 223.3000 3.7000 ;
	    RECT 221.9000 3.1000 222.2000 3.4000 ;
	    RECT 224.6000 3.1000 225.0000 3.5000 ;
	    RECT 219.5000 1.1000 220.1000 3.1000 ;
	    RECT 221.8000 1.1000 222.2000 3.1000 ;
	    RECT 224.0000 2.8000 225.0000 3.1000 ;
	    RECT 224.0000 1.1000 224.4000 2.8000 ;
	    RECT 226.2000 1.1000 226.6000 5.3000 ;
	    RECT 227.8000 1.1000 228.2000 6.8000 ;
	    RECT 229.4000 5.4000 229.8000 6.2000 ;
	    RECT 230.1000 4.9000 230.4000 6.8000 ;
	    RECT 230.7000 6.5000 231.4000 6.9000 ;
	    RECT 231.1000 5.5000 231.4000 6.5000 ;
	    RECT 231.8000 5.8000 232.2000 6.6000 ;
	    RECT 232.6000 5.8000 233.0000 6.6000 ;
	    RECT 234.2000 6.1000 234.6000 9.9000 ;
	    RECT 235.8000 8.9000 236.2000 9.9000 ;
	    RECT 235.8000 7.2000 236.1000 8.9000 ;
	    RECT 236.6000 8.1000 237.0000 8.6000 ;
	    RECT 237.4000 8.1000 237.8000 9.9000 ;
	    RECT 239.8000 8.9000 240.2000 9.9000 ;
	    RECT 236.6000 7.8000 237.8000 8.1000 ;
	    RECT 238.2000 8.1000 238.6000 8.6000 ;
	    RECT 239.8000 8.1000 240.1000 8.9000 ;
	    RECT 238.2000 7.8000 240.1000 8.1000 ;
	    RECT 241.4000 7.8000 241.8000 8.6000 ;
	    RECT 235.8000 6.8000 236.2000 7.2000 ;
	    RECT 235.0000 6.1000 235.4000 6.2000 ;
	    RECT 234.2000 5.8000 235.4000 6.1000 ;
	    RECT 231.1000 5.2000 233.0000 5.5000 ;
	    RECT 230.1000 4.6000 230.9000 4.9000 ;
	    RECT 230.5000 1.1000 230.9000 4.6000 ;
	    RECT 232.7000 3.5000 233.0000 5.2000 ;
	    RECT 232.6000 1.5000 233.0000 3.5000 ;
	    RECT 234.2000 1.1000 234.6000 5.8000 ;
	    RECT 235.0000 5.4000 235.4000 5.8000 ;
	    RECT 235.8000 6.1000 236.1000 6.8000 ;
	    RECT 236.6000 6.1000 237.0000 6.2000 ;
	    RECT 235.8000 5.8000 237.0000 6.1000 ;
	    RECT 235.8000 5.1000 236.1000 5.8000 ;
	    RECT 235.3000 4.7000 236.2000 5.1000 ;
	    RECT 235.3000 1.1000 235.7000 4.7000 ;
	    RECT 237.4000 1.1000 237.8000 7.8000 ;
	    RECT 239.8000 7.2000 240.1000 7.8000 ;
	    RECT 239.8000 6.8000 240.2000 7.2000 ;
	    RECT 242.2000 7.1000 242.6000 9.9000 ;
	    RECT 243.0000 9.6000 245.0000 9.9000 ;
	    RECT 243.0000 7.9000 243.4000 9.6000 ;
	    RECT 243.8000 7.9000 244.2000 9.3000 ;
	    RECT 244.6000 8.0000 245.0000 9.6000 ;
	    RECT 246.2000 8.0000 246.6000 9.9000 ;
	    RECT 244.6000 7.9000 246.6000 8.0000 ;
	    RECT 247.3000 8.2000 247.7000 9.9000 ;
	    RECT 247.3000 7.9000 248.2000 8.2000 ;
	    RECT 243.8000 7.2000 244.1000 7.9000 ;
	    RECT 244.7000 7.7000 246.5000 7.9000 ;
	    RECT 245.8000 7.2000 246.2000 7.4000 ;
	    RECT 243.0000 7.1000 243.4000 7.2000 ;
	    RECT 242.2000 6.8000 243.4000 7.1000 ;
	    RECT 243.8000 6.9000 245.0000 7.2000 ;
	    RECT 245.8000 7.1000 246.6000 7.2000 ;
	    RECT 247.8000 7.1000 248.2000 7.9000 ;
	    RECT 249.4000 7.8000 249.8000 8.6000 ;
	    RECT 245.8000 6.9000 248.2000 7.1000 ;
	    RECT 244.6000 6.8000 245.0000 6.9000 ;
	    RECT 246.2000 6.8000 248.2000 6.9000 ;
	    RECT 248.6000 6.8000 249.0000 7.6000 ;
	    RECT 239.0000 5.4000 239.4000 6.2000 ;
	    RECT 239.8000 5.2000 240.1000 6.8000 ;
	    RECT 239.8000 5.1000 240.2000 5.2000 ;
	    RECT 239.3000 4.7000 240.2000 5.1000 ;
	    RECT 239.3000 1.1000 239.7000 4.7000 ;
	    RECT 242.2000 1.1000 242.6000 6.8000 ;
	    RECT 243.0000 5.8000 243.4000 6.8000 ;
	    RECT 243.8000 5.8000 244.2000 6.6000 ;
	    RECT 244.7000 5.1000 245.0000 6.8000 ;
	    RECT 245.4000 5.8000 245.8000 6.6000 ;
	    RECT 247.8000 6.1000 248.2000 6.8000 ;
	    RECT 249.4000 6.1000 249.8000 6.2000 ;
	    RECT 247.8000 5.8000 249.8000 6.1000 ;
	    RECT 250.2000 6.1000 250.6000 9.9000 ;
	    RECT 252.6000 7.9000 253.0000 9.9000 ;
	    RECT 255.0000 8.8000 255.4000 9.9000 ;
	    RECT 253.3000 8.2000 253.7000 8.6000 ;
	    RECT 251.8000 6.4000 252.2000 7.2000 ;
	    RECT 251.0000 6.1000 251.4000 6.2000 ;
	    RECT 252.6000 6.1000 252.9000 7.9000 ;
	    RECT 253.4000 7.8000 253.8000 8.2000 ;
	    RECT 255.0000 7.2000 255.3000 8.8000 ;
	    RECT 255.8000 7.8000 256.2000 8.6000 ;
	    RECT 255.0000 6.8000 255.4000 7.2000 ;
	    RECT 255.8000 6.8000 256.2000 7.2000 ;
	    RECT 253.4000 6.1000 253.8000 6.2000 ;
	    RECT 250.2000 5.8000 251.8000 6.1000 ;
	    RECT 252.6000 5.8000 253.8000 6.1000 ;
	    RECT 244.3000 1.1000 245.3000 5.1000 ;
	    RECT 247.0000 4.4000 247.4000 5.2000 ;
	    RECT 247.8000 1.1000 248.2000 5.8000 ;
	    RECT 250.2000 1.1000 250.6000 5.8000 ;
	    RECT 251.4000 5.6000 251.8000 5.8000 ;
	    RECT 253.4000 5.1000 253.7000 5.8000 ;
	    RECT 254.2000 5.4000 254.6000 6.2000 ;
	    RECT 255.0000 5.1000 255.3000 6.8000 ;
	    RECT 255.8000 6.1000 256.1000 6.8000 ;
	    RECT 256.6000 6.1000 257.0000 9.9000 ;
	    RECT 259.0000 8.9000 259.4000 9.9000 ;
	    RECT 261.9000 9.2000 262.3000 9.9000 ;
	    RECT 257.4000 7.8000 257.8000 8.6000 ;
	    RECT 259.1000 8.1000 259.4000 8.9000 ;
	    RECT 261.4000 8.8000 262.3000 9.2000 ;
	    RECT 261.9000 8.2000 262.3000 8.8000 ;
	    RECT 259.8000 8.1000 260.2000 8.2000 ;
	    RECT 259.0000 7.8000 260.2000 8.1000 ;
	    RECT 261.4000 7.9000 262.3000 8.2000 ;
	    RECT 264.6000 7.9000 265.0000 9.9000 ;
	    RECT 265.3000 8.2000 265.7000 8.6000 ;
	    RECT 259.1000 7.2000 259.4000 7.8000 ;
	    RECT 259.0000 6.8000 259.4000 7.2000 ;
	    RECT 255.8000 5.8000 257.0000 6.1000 ;
	    RECT 251.0000 4.8000 253.0000 5.1000 ;
	    RECT 251.0000 1.1000 251.4000 4.8000 ;
	    RECT 252.6000 1.1000 253.0000 4.8000 ;
	    RECT 253.4000 1.1000 253.8000 5.1000 ;
	    RECT 254.5000 4.7000 255.4000 5.1000 ;
	    RECT 254.5000 1.1000 254.9000 4.7000 ;
	    RECT 256.6000 1.1000 257.0000 5.8000 ;
	    RECT 259.1000 5.1000 259.4000 6.8000 ;
	    RECT 259.8000 6.1000 260.2000 6.2000 ;
	    RECT 260.6000 6.1000 261.0000 6.2000 ;
	    RECT 259.8000 5.8000 261.0000 6.1000 ;
	    RECT 259.8000 5.4000 260.2000 5.8000 ;
	    RECT 259.0000 4.7000 259.9000 5.1000 ;
	    RECT 259.5000 1.1000 259.9000 4.7000 ;
	    RECT 261.4000 1.1000 261.8000 7.9000 ;
	    RECT 263.8000 6.4000 264.2000 7.2000 ;
	    RECT 263.0000 6.1000 263.4000 6.2000 ;
	    RECT 264.6000 6.1000 264.9000 7.9000 ;
	    RECT 265.4000 7.8000 265.8000 8.2000 ;
	    RECT 267.8000 7.6000 268.2000 9.9000 ;
	    RECT 268.6000 7.8000 269.0000 8.6000 ;
	    RECT 267.1000 7.3000 268.2000 7.6000 ;
	    RECT 265.4000 6.1000 265.8000 6.2000 ;
	    RECT 263.0000 5.8000 263.8000 6.1000 ;
	    RECT 264.6000 5.8000 265.8000 6.1000 ;
	    RECT 267.1000 5.8000 267.4000 7.3000 ;
	    RECT 267.8000 5.8000 268.2000 6.6000 ;
	    RECT 263.4000 5.6000 263.8000 5.8000 ;
	    RECT 262.2000 4.4000 262.6000 5.2000 ;
	    RECT 265.4000 5.1000 265.7000 5.8000 ;
	    RECT 266.8000 5.4000 267.4000 5.8000 ;
	    RECT 267.1000 5.1000 267.4000 5.4000 ;
	    RECT 263.0000 4.8000 265.0000 5.1000 ;
	    RECT 263.0000 1.1000 263.4000 4.8000 ;
	    RECT 264.6000 1.1000 265.0000 4.8000 ;
	    RECT 265.4000 1.1000 265.8000 5.1000 ;
	    RECT 267.1000 4.8000 268.2000 5.1000 ;
	    RECT 267.8000 1.1000 268.2000 4.8000 ;
	    RECT 269.4000 1.1000 269.8000 9.9000 ;
         LAYER metal2 ;
	    RECT 10.2000 176.8000 10.6000 177.2000 ;
	    RECT 10.2000 176.2000 10.5000 176.8000 ;
	    RECT 0.6000 176.1000 1.0000 176.2000 ;
	    RECT 1.4000 176.1000 1.8000 176.2000 ;
	    RECT 0.6000 175.8000 1.8000 176.1000 ;
	    RECT 5.4000 176.1000 5.8000 176.2000 ;
	    RECT 6.2000 176.1000 6.6000 176.2000 ;
	    RECT 5.4000 175.8000 6.6000 176.1000 ;
	    RECT 8.6000 176.1000 9.0000 176.2000 ;
	    RECT 9.4000 176.1000 9.8000 176.2000 ;
	    RECT 8.6000 175.8000 9.8000 176.1000 ;
	    RECT 10.2000 175.8000 10.6000 176.2000 ;
	    RECT 8.6000 174.2000 8.9000 175.8000 ;
	    RECT 49.4000 174.8000 49.8000 175.2000 ;
	    RECT 3.8000 173.8000 4.2000 174.2000 ;
	    RECT 5.4000 174.1000 5.8000 174.2000 ;
	    RECT 6.2000 174.1000 6.6000 174.2000 ;
	    RECT 5.4000 173.8000 6.6000 174.1000 ;
	    RECT 8.6000 173.8000 9.0000 174.2000 ;
	    RECT 25.4000 174.1000 25.8000 174.2000 ;
	    RECT 26.2000 174.1000 26.6000 174.2000 ;
	    RECT 25.4000 173.8000 26.6000 174.1000 ;
	    RECT 30.2000 174.1000 30.6000 174.2000 ;
	    RECT 31.0000 174.1000 31.4000 174.2000 ;
	    RECT 30.2000 173.8000 31.4000 174.1000 ;
	    RECT 3.0000 165.1000 3.4000 165.2000 ;
	    RECT 3.8000 165.1000 4.1000 173.8000 ;
	    RECT 30.2000 172.8000 30.6000 173.2000 ;
	    RECT 30.2000 172.2000 30.5000 172.8000 ;
	    RECT 49.4000 172.2000 49.7000 174.8000 ;
	    RECT 7.0000 171.8000 7.4000 172.2000 ;
	    RECT 8.6000 171.8000 9.0000 172.2000 ;
	    RECT 13.4000 172.1000 13.8000 172.2000 ;
	    RECT 14.2000 172.1000 14.6000 172.2000 ;
	    RECT 13.4000 171.8000 14.6000 172.1000 ;
	    RECT 19.8000 172.1000 20.2000 172.2000 ;
	    RECT 20.6000 172.1000 21.0000 172.2000 ;
	    RECT 19.8000 171.8000 21.0000 172.1000 ;
	    RECT 27.0000 171.8000 27.4000 172.2000 ;
	    RECT 27.8000 171.8000 28.2000 172.2000 ;
	    RECT 30.2000 171.8000 30.6000 172.2000 ;
	    RECT 32.6000 171.8000 33.0000 172.2000 ;
	    RECT 35.0000 171.8000 35.4000 172.2000 ;
	    RECT 39.0000 171.8000 39.4000 172.2000 ;
	    RECT 43.8000 171.8000 44.2000 172.2000 ;
	    RECT 47.0000 171.8000 47.4000 172.2000 ;
	    RECT 49.4000 171.8000 49.8000 172.2000 ;
	    RECT 51.8000 172.1000 52.2000 172.2000 ;
	    RECT 52.6000 172.1000 53.0000 172.2000 ;
	    RECT 54.2000 172.1000 54.6000 177.9000 ;
	    RECT 58.2000 174.7000 58.6000 175.1000 ;
	    RECT 58.2000 174.2000 58.5000 174.7000 ;
	    RECT 58.2000 173.8000 58.6000 174.2000 ;
	    RECT 59.0000 172.1000 59.4000 177.9000 ;
	    RECT 60.6000 173.1000 61.0000 175.9000 ;
	    RECT 63.0000 173.1000 63.4000 175.9000 ;
	    RECT 51.8000 171.8000 53.0000 172.1000 ;
	    RECT 62.2000 171.8000 62.6000 172.2000 ;
	    RECT 64.6000 172.1000 65.0000 177.9000 ;
	    RECT 65.4000 174.8000 65.8000 175.2000 ;
	    RECT 67.8000 174.8000 68.2000 175.2000 ;
	    RECT 7.0000 168.1000 7.3000 171.8000 ;
	    RECT 7.0000 167.8000 8.1000 168.1000 ;
	    RECT 6.2000 167.1000 6.6000 167.2000 ;
	    RECT 7.0000 167.1000 7.4000 167.2000 ;
	    RECT 6.2000 166.8000 7.4000 167.1000 ;
	    RECT 3.0000 164.8000 4.1000 165.1000 ;
	    RECT 7.8000 165.2000 8.1000 167.8000 ;
	    RECT 8.6000 166.2000 8.9000 171.8000 ;
	    RECT 11.0000 166.8000 11.4000 167.2000 ;
	    RECT 25.4000 166.8000 25.8000 167.2000 ;
	    RECT 11.0000 166.2000 11.3000 166.8000 ;
	    RECT 25.4000 166.2000 25.7000 166.8000 ;
	    RECT 8.6000 165.8000 9.0000 166.2000 ;
	    RECT 11.0000 165.8000 11.4000 166.2000 ;
	    RECT 23.0000 166.1000 23.4000 166.2000 ;
	    RECT 23.8000 166.1000 24.2000 166.2000 ;
	    RECT 23.0000 165.8000 24.2000 166.1000 ;
	    RECT 25.4000 165.8000 25.8000 166.2000 ;
	    RECT 7.8000 164.8000 8.2000 165.2000 ;
	    RECT 13.4000 164.8000 13.8000 165.2000 ;
	    RECT 13.4000 164.2000 13.7000 164.8000 ;
	    RECT 27.0000 164.2000 27.3000 171.8000 ;
	    RECT 27.8000 165.2000 28.1000 171.8000 ;
	    RECT 31.8000 167.8000 32.2000 168.2000 ;
	    RECT 32.6000 168.1000 32.9000 171.8000 ;
	    RECT 35.0000 168.2000 35.3000 171.8000 ;
	    RECT 32.6000 167.8000 33.7000 168.1000 ;
	    RECT 35.0000 167.8000 35.4000 168.2000 ;
	    RECT 28.6000 166.1000 29.0000 166.2000 ;
	    RECT 29.4000 166.1000 29.8000 166.2000 ;
	    RECT 28.6000 165.8000 29.8000 166.1000 ;
	    RECT 27.8000 164.8000 28.2000 165.2000 ;
	    RECT 9.4000 164.1000 9.8000 164.2000 ;
	    RECT 10.2000 164.1000 10.6000 164.2000 ;
	    RECT 9.4000 163.8000 10.6000 164.1000 ;
	    RECT 13.4000 163.8000 13.8000 164.2000 ;
	    RECT 27.0000 163.8000 27.4000 164.2000 ;
	    RECT 4.6000 161.8000 5.0000 162.2000 ;
	    RECT 8.6000 161.8000 9.0000 162.2000 ;
	    RECT 16.6000 161.8000 17.0000 162.2000 ;
	    RECT 20.6000 161.8000 21.0000 162.2000 ;
	    RECT 24.6000 161.8000 25.0000 162.2000 ;
	    RECT 28.6000 161.8000 29.0000 162.2000 ;
	    RECT 4.6000 156.2000 4.9000 161.8000 ;
	    RECT 4.6000 155.8000 5.0000 156.2000 ;
	    RECT 3.0000 152.1000 3.4000 152.2000 ;
	    RECT 3.8000 152.1000 4.2000 152.2000 ;
	    RECT 3.0000 151.8000 4.2000 152.1000 ;
	    RECT 6.2000 151.8000 6.6000 152.2000 ;
	    RECT 5.4000 149.8000 5.8000 150.2000 ;
	    RECT 5.4000 149.2000 5.7000 149.8000 ;
	    RECT 0.6000 148.8000 1.0000 149.2000 ;
	    RECT 5.4000 148.8000 5.8000 149.2000 ;
	    RECT 0.6000 148.2000 0.9000 148.8000 ;
	    RECT 0.6000 147.8000 1.0000 148.2000 ;
	    RECT 6.2000 147.2000 6.5000 151.8000 ;
	    RECT 8.6000 149.2000 8.9000 161.8000 ;
	    RECT 16.6000 159.2000 16.9000 161.8000 ;
	    RECT 13.4000 158.8000 13.8000 159.2000 ;
	    RECT 16.6000 158.8000 17.0000 159.2000 ;
	    RECT 13.4000 156.2000 13.7000 158.8000 ;
	    RECT 20.6000 157.2000 20.9000 161.8000 ;
	    RECT 14.2000 156.8000 14.6000 157.2000 ;
	    RECT 15.8000 157.1000 16.2000 157.2000 ;
	    RECT 16.6000 157.1000 17.0000 157.2000 ;
	    RECT 15.8000 156.8000 17.0000 157.1000 ;
	    RECT 20.6000 156.8000 21.0000 157.2000 ;
	    RECT 14.2000 156.2000 14.5000 156.8000 ;
	    RECT 13.4000 155.8000 13.8000 156.2000 ;
	    RECT 14.2000 155.8000 14.6000 156.2000 ;
	    RECT 13.4000 154.8000 13.8000 155.2000 ;
	    RECT 14.2000 155.1000 14.6000 155.2000 ;
	    RECT 15.0000 155.1000 15.4000 155.2000 ;
	    RECT 20.6000 155.1000 20.9000 156.8000 ;
	    RECT 24.6000 155.2000 24.9000 161.8000 ;
	    RECT 26.2000 157.8000 26.6000 158.2000 ;
	    RECT 25.4000 155.8000 25.8000 156.2000 ;
	    RECT 14.2000 154.8000 15.4000 155.1000 ;
	    RECT 19.8000 154.8000 20.9000 155.1000 ;
	    RECT 21.4000 154.8000 21.8000 155.2000 ;
	    RECT 24.6000 154.8000 25.0000 155.2000 ;
	    RECT 13.4000 154.2000 13.7000 154.8000 ;
	    RECT 9.4000 153.8000 9.8000 154.2000 ;
	    RECT 13.4000 153.8000 13.8000 154.2000 ;
	    RECT 19.0000 153.8000 19.4000 154.2000 ;
	    RECT 8.6000 148.8000 9.0000 149.2000 ;
	    RECT 9.4000 147.2000 9.7000 153.8000 ;
	    RECT 19.0000 153.2000 19.3000 153.8000 ;
	    RECT 19.8000 153.2000 20.1000 154.8000 ;
	    RECT 20.6000 154.1000 21.0000 154.2000 ;
	    RECT 21.4000 154.1000 21.7000 154.8000 ;
	    RECT 20.6000 153.8000 21.7000 154.1000 ;
	    RECT 23.0000 154.1000 23.4000 154.2000 ;
	    RECT 23.8000 154.1000 24.2000 154.2000 ;
	    RECT 23.0000 153.8000 24.2000 154.1000 ;
	    RECT 25.4000 153.2000 25.7000 155.8000 ;
	    RECT 26.2000 153.2000 26.5000 157.8000 ;
	    RECT 27.8000 155.1000 28.2000 155.2000 ;
	    RECT 28.6000 155.1000 28.9000 161.8000 ;
	    RECT 29.4000 156.8000 29.8000 157.2000 ;
	    RECT 29.4000 156.2000 29.7000 156.8000 ;
	    RECT 29.4000 155.8000 29.8000 156.2000 ;
	    RECT 31.0000 156.1000 31.4000 156.2000 ;
	    RECT 31.8000 156.1000 32.1000 167.8000 ;
	    RECT 32.6000 166.8000 33.0000 167.2000 ;
	    RECT 32.6000 166.2000 32.9000 166.8000 ;
	    RECT 32.6000 165.8000 33.0000 166.2000 ;
	    RECT 33.4000 166.1000 33.7000 167.8000 ;
	    RECT 35.0000 167.1000 35.4000 167.2000 ;
	    RECT 35.8000 167.1000 36.2000 167.2000 ;
	    RECT 35.0000 166.8000 36.2000 167.1000 ;
	    RECT 34.2000 166.1000 34.6000 166.2000 ;
	    RECT 33.4000 165.8000 34.6000 166.1000 ;
	    RECT 35.0000 158.2000 35.3000 166.8000 ;
	    RECT 37.4000 165.1000 37.8000 165.2000 ;
	    RECT 38.2000 165.1000 38.6000 165.2000 ;
	    RECT 37.4000 164.8000 38.6000 165.1000 ;
	    RECT 39.0000 163.1000 39.3000 171.8000 ;
	    RECT 43.0000 167.8000 43.4000 168.2000 ;
	    RECT 41.4000 167.1000 41.8000 167.2000 ;
	    RECT 42.2000 167.1000 42.6000 167.2000 ;
	    RECT 41.4000 166.8000 42.6000 167.1000 ;
	    RECT 43.0000 166.2000 43.3000 167.8000 ;
	    RECT 43.0000 165.8000 43.4000 166.2000 ;
	    RECT 43.8000 165.2000 44.1000 171.8000 ;
	    RECT 47.0000 168.2000 47.3000 171.8000 ;
	    RECT 62.2000 168.2000 62.5000 171.8000 ;
	    RECT 65.4000 169.2000 65.7000 174.8000 ;
	    RECT 66.2000 173.8000 66.6000 174.2000 ;
	    RECT 65.4000 168.8000 65.8000 169.2000 ;
	    RECT 47.0000 167.8000 47.4000 168.2000 ;
	    RECT 51.0000 168.1000 51.4000 168.2000 ;
	    RECT 51.8000 168.1000 52.2000 168.2000 ;
	    RECT 51.0000 167.8000 52.2000 168.1000 ;
	    RECT 56.6000 167.8000 57.0000 168.2000 ;
	    RECT 62.2000 167.8000 62.6000 168.2000 ;
	    RECT 56.6000 167.2000 56.9000 167.8000 ;
	    RECT 51.8000 167.1000 52.2000 167.2000 ;
	    RECT 52.6000 167.1000 53.0000 167.2000 ;
	    RECT 51.8000 166.8000 53.0000 167.1000 ;
	    RECT 55.0000 166.8000 55.4000 167.2000 ;
	    RECT 56.6000 166.8000 57.0000 167.2000 ;
	    RECT 58.2000 166.8000 58.6000 167.2000 ;
	    RECT 60.6000 167.1000 61.0000 167.2000 ;
	    RECT 61.4000 167.1000 61.8000 167.2000 ;
	    RECT 60.6000 166.8000 61.8000 167.1000 ;
	    RECT 64.6000 166.8000 65.0000 167.2000 ;
	    RECT 55.0000 166.2000 55.3000 166.8000 ;
	    RECT 58.2000 166.2000 58.5000 166.8000 ;
	    RECT 50.2000 166.1000 50.6000 166.2000 ;
	    RECT 51.0000 166.1000 51.4000 166.2000 ;
	    RECT 50.2000 165.8000 51.4000 166.1000 ;
	    RECT 53.4000 166.1000 53.8000 166.2000 ;
	    RECT 54.2000 166.1000 54.6000 166.2000 ;
	    RECT 53.4000 165.8000 54.6000 166.1000 ;
	    RECT 55.0000 165.8000 55.4000 166.2000 ;
	    RECT 58.2000 165.8000 58.6000 166.2000 ;
	    RECT 43.8000 164.8000 44.2000 165.2000 ;
	    RECT 55.0000 164.8000 55.4000 165.2000 ;
	    RECT 61.4000 165.1000 61.8000 165.2000 ;
	    RECT 62.2000 165.1000 62.6000 165.2000 ;
	    RECT 61.4000 164.8000 62.6000 165.1000 ;
	    RECT 55.0000 164.2000 55.3000 164.8000 ;
	    RECT 64.6000 164.2000 64.9000 166.8000 ;
	    RECT 42.2000 164.1000 42.6000 164.2000 ;
	    RECT 43.0000 164.1000 43.4000 164.2000 ;
	    RECT 42.2000 163.8000 43.4000 164.1000 ;
	    RECT 47.0000 164.1000 47.4000 164.2000 ;
	    RECT 47.8000 164.1000 48.2000 164.2000 ;
	    RECT 47.0000 163.8000 48.2000 164.1000 ;
	    RECT 55.0000 163.8000 55.4000 164.2000 ;
	    RECT 61.4000 163.8000 61.8000 164.2000 ;
	    RECT 64.6000 163.8000 65.0000 164.2000 ;
	    RECT 38.2000 162.8000 39.3000 163.1000 ;
	    RECT 35.8000 161.8000 36.2000 162.2000 ;
	    RECT 35.0000 157.8000 35.4000 158.2000 ;
	    RECT 35.8000 157.2000 36.1000 161.8000 ;
	    RECT 35.8000 156.8000 36.2000 157.2000 ;
	    RECT 31.0000 155.8000 32.1000 156.1000 ;
	    RECT 33.4000 155.8000 33.8000 156.2000 ;
	    RECT 35.0000 155.8000 35.4000 156.2000 ;
	    RECT 33.4000 155.2000 33.7000 155.8000 ;
	    RECT 35.0000 155.2000 35.3000 155.8000 ;
	    RECT 27.8000 154.8000 28.9000 155.1000 ;
	    RECT 30.2000 154.8000 30.6000 155.2000 ;
	    RECT 31.8000 155.1000 32.2000 155.2000 ;
	    RECT 32.6000 155.1000 33.0000 155.2000 ;
	    RECT 31.8000 154.8000 33.0000 155.1000 ;
	    RECT 33.4000 154.8000 33.8000 155.2000 ;
	    RECT 35.0000 154.8000 35.4000 155.2000 ;
	    RECT 35.8000 155.1000 36.2000 155.2000 ;
	    RECT 36.6000 155.1000 37.0000 155.2000 ;
	    RECT 35.8000 154.8000 37.0000 155.1000 ;
	    RECT 30.2000 154.2000 30.5000 154.8000 ;
	    RECT 38.2000 154.2000 38.5000 162.8000 ;
	    RECT 39.0000 161.8000 39.4000 162.2000 ;
	    RECT 40.6000 161.8000 41.0000 162.2000 ;
	    RECT 39.0000 156.2000 39.3000 161.8000 ;
	    RECT 39.0000 155.8000 39.4000 156.2000 ;
	    RECT 40.6000 155.2000 40.9000 161.8000 ;
	    RECT 47.0000 157.8000 47.4000 158.2000 ;
	    RECT 50.2000 158.1000 50.6000 158.2000 ;
	    RECT 51.0000 158.1000 51.4000 158.2000 ;
	    RECT 50.2000 157.8000 51.4000 158.1000 ;
	    RECT 43.8000 155.8000 44.2000 156.2000 ;
	    RECT 40.6000 154.8000 41.0000 155.2000 ;
	    RECT 40.6000 154.2000 40.9000 154.8000 ;
	    RECT 27.8000 153.8000 28.2000 154.2000 ;
	    RECT 30.2000 153.8000 30.6000 154.2000 ;
	    RECT 38.2000 153.8000 38.6000 154.2000 ;
	    RECT 39.0000 153.8000 39.4000 154.2000 ;
	    RECT 40.6000 153.8000 41.0000 154.2000 ;
	    RECT 43.0000 153.8000 43.4000 154.2000 ;
	    RECT 27.8000 153.2000 28.1000 153.8000 ;
	    RECT 38.2000 153.2000 38.5000 153.8000 ;
	    RECT 39.0000 153.2000 39.3000 153.8000 ;
	    RECT 43.0000 153.2000 43.3000 153.8000 ;
	    RECT 19.0000 152.8000 19.4000 153.2000 ;
	    RECT 19.8000 152.8000 20.2000 153.2000 ;
	    RECT 25.4000 152.8000 25.8000 153.2000 ;
	    RECT 26.2000 152.8000 26.6000 153.2000 ;
	    RECT 27.8000 152.8000 28.2000 153.2000 ;
	    RECT 38.2000 152.8000 38.6000 153.2000 ;
	    RECT 39.0000 152.8000 39.4000 153.2000 ;
	    RECT 40.6000 153.1000 41.0000 153.2000 ;
	    RECT 41.4000 153.1000 41.8000 153.2000 ;
	    RECT 40.6000 152.8000 41.8000 153.1000 ;
	    RECT 43.0000 152.8000 43.4000 153.2000 ;
	    RECT 10.2000 151.8000 10.6000 152.2000 ;
	    RECT 15.8000 151.8000 16.2000 152.2000 ;
	    RECT 18.2000 151.8000 18.6000 152.2000 ;
	    RECT 25.4000 151.8000 25.8000 152.2000 ;
	    RECT 27.0000 151.8000 27.4000 152.2000 ;
	    RECT 10.2000 149.2000 10.5000 151.8000 ;
	    RECT 10.2000 148.8000 10.6000 149.2000 ;
	    RECT 6.2000 146.8000 6.6000 147.2000 ;
	    RECT 9.4000 146.8000 9.8000 147.2000 ;
	    RECT 2.2000 145.8000 2.6000 146.2000 ;
	    RECT 3.8000 146.1000 4.2000 146.2000 ;
	    RECT 4.6000 146.1000 5.0000 146.2000 ;
	    RECT 3.8000 145.8000 5.0000 146.1000 ;
	    RECT 7.8000 146.1000 8.2000 146.2000 ;
	    RECT 8.6000 146.1000 9.0000 146.2000 ;
	    RECT 7.8000 145.8000 9.0000 146.1000 ;
	    RECT 1.4000 141.8000 1.8000 142.2000 ;
	    RECT 1.4000 138.2000 1.7000 141.8000 ;
	    RECT 2.2000 139.2000 2.5000 145.8000 ;
	    RECT 5.4000 145.1000 5.8000 145.2000 ;
	    RECT 6.2000 145.1000 6.6000 145.2000 ;
	    RECT 5.4000 144.8000 6.6000 145.1000 ;
	    RECT 7.8000 144.8000 8.2000 145.2000 ;
	    RECT 8.6000 145.1000 9.0000 145.2000 ;
	    RECT 9.4000 145.1000 9.8000 145.2000 ;
	    RECT 8.6000 144.8000 9.8000 145.1000 ;
	    RECT 10.2000 145.1000 10.6000 145.2000 ;
	    RECT 11.0000 145.1000 11.4000 145.2000 ;
	    RECT 10.2000 144.8000 11.4000 145.1000 ;
	    RECT 13.4000 145.1000 13.8000 145.2000 ;
	    RECT 14.2000 145.1000 14.6000 145.2000 ;
	    RECT 13.4000 144.8000 14.6000 145.1000 ;
	    RECT 2.2000 138.8000 2.6000 139.2000 ;
	    RECT 1.4000 137.8000 1.8000 138.2000 ;
	    RECT 1.4000 136.8000 1.8000 137.2000 ;
	    RECT 1.4000 129.2000 1.7000 136.8000 ;
	    RECT 7.0000 135.8000 7.4000 136.2000 ;
	    RECT 7.0000 135.2000 7.3000 135.8000 ;
	    RECT 2.2000 134.8000 2.6000 135.2000 ;
	    RECT 7.0000 135.1000 7.4000 135.2000 ;
	    RECT 6.2000 134.8000 7.4000 135.1000 ;
	    RECT 2.2000 133.2000 2.5000 134.8000 ;
	    RECT 6.2000 133.2000 6.5000 134.8000 ;
	    RECT 7.0000 133.8000 7.4000 134.2000 ;
	    RECT 7.0000 133.2000 7.3000 133.8000 ;
	    RECT 2.2000 132.8000 2.6000 133.2000 ;
	    RECT 6.2000 132.8000 6.6000 133.2000 ;
	    RECT 7.0000 132.8000 7.4000 133.2000 ;
	    RECT 7.8000 129.2000 8.1000 144.8000 ;
	    RECT 15.8000 144.2000 16.1000 151.8000 ;
	    RECT 16.6000 148.8000 17.0000 149.2000 ;
	    RECT 16.6000 146.2000 16.9000 148.8000 ;
	    RECT 18.2000 148.2000 18.5000 151.8000 ;
	    RECT 24.6000 149.8000 25.0000 150.2000 ;
	    RECT 18.2000 147.8000 18.6000 148.2000 ;
	    RECT 23.8000 147.8000 24.2000 148.2000 ;
	    RECT 20.6000 146.8000 21.0000 147.2000 ;
	    RECT 21.4000 146.8000 21.8000 147.2000 ;
	    RECT 23.0000 146.8000 23.4000 147.2000 ;
	    RECT 16.6000 145.8000 17.0000 146.2000 ;
	    RECT 17.4000 145.1000 17.8000 145.2000 ;
	    RECT 18.2000 145.1000 18.6000 145.2000 ;
	    RECT 17.4000 144.8000 18.6000 145.1000 ;
	    RECT 20.6000 145.1000 20.9000 146.8000 ;
	    RECT 21.4000 146.2000 21.7000 146.8000 ;
	    RECT 23.0000 146.2000 23.3000 146.8000 ;
	    RECT 23.8000 146.2000 24.1000 147.8000 ;
	    RECT 24.6000 147.2000 24.9000 149.8000 ;
	    RECT 25.4000 148.1000 25.7000 151.8000 ;
	    RECT 26.2000 148.1000 26.6000 148.2000 ;
	    RECT 25.4000 147.8000 26.6000 148.1000 ;
	    RECT 24.6000 146.8000 25.0000 147.2000 ;
	    RECT 27.0000 146.2000 27.3000 151.8000 ;
	    RECT 43.8000 150.2000 44.1000 155.8000 ;
	    RECT 47.0000 155.2000 47.3000 157.8000 ;
	    RECT 49.4000 156.8000 49.8000 157.2000 ;
	    RECT 49.4000 156.2000 49.7000 156.8000 ;
	    RECT 49.4000 155.8000 49.8000 156.2000 ;
	    RECT 47.0000 154.8000 47.4000 155.2000 ;
	    RECT 50.2000 155.1000 50.6000 155.2000 ;
	    RECT 51.0000 155.1000 51.4000 155.2000 ;
	    RECT 50.2000 154.8000 51.4000 155.1000 ;
	    RECT 47.0000 153.2000 47.3000 154.8000 ;
	    RECT 47.0000 152.8000 47.4000 153.2000 ;
	    RECT 53.4000 152.1000 53.8000 157.9000 ;
	    RECT 56.6000 155.8000 57.0000 156.2000 ;
	    RECT 56.6000 155.2000 56.9000 155.8000 ;
	    RECT 56.6000 154.8000 57.0000 155.2000 ;
	    RECT 58.2000 152.1000 58.6000 157.9000 ;
	    RECT 59.8000 153.1000 60.2000 155.9000 ;
	    RECT 60.6000 151.8000 61.0000 152.2000 ;
	    RECT 43.8000 149.8000 44.2000 150.2000 ;
	    RECT 53.4000 149.8000 53.8000 150.2000 ;
	    RECT 29.4000 148.8000 29.8000 149.2000 ;
	    RECT 29.4000 148.2000 29.7000 148.8000 ;
	    RECT 27.8000 147.8000 28.2000 148.2000 ;
	    RECT 29.4000 147.8000 29.8000 148.2000 ;
	    RECT 27.8000 147.2000 28.1000 147.8000 ;
	    RECT 27.8000 146.8000 28.2000 147.2000 ;
	    RECT 21.4000 145.8000 21.8000 146.2000 ;
	    RECT 23.0000 145.8000 23.4000 146.2000 ;
	    RECT 23.8000 145.8000 24.2000 146.2000 ;
	    RECT 27.0000 145.8000 27.4000 146.2000 ;
	    RECT 20.6000 144.8000 21.7000 145.1000 ;
	    RECT 15.8000 143.8000 16.2000 144.2000 ;
	    RECT 16.6000 141.8000 17.0000 142.2000 ;
	    RECT 16.6000 137.2000 16.9000 141.8000 ;
	    RECT 21.4000 139.2000 21.7000 144.8000 ;
	    RECT 23.0000 144.8000 23.4000 145.2000 ;
	    RECT 21.4000 138.8000 21.8000 139.2000 ;
	    RECT 15.0000 136.8000 15.4000 137.2000 ;
	    RECT 16.6000 136.8000 17.0000 137.2000 ;
	    RECT 22.2000 136.8000 22.6000 137.2000 ;
	    RECT 15.0000 136.2000 15.3000 136.8000 ;
	    RECT 15.0000 135.8000 15.4000 136.2000 ;
	    RECT 15.8000 136.1000 16.2000 136.2000 ;
	    RECT 16.6000 136.1000 17.0000 136.2000 ;
	    RECT 15.8000 135.8000 17.0000 136.1000 ;
	    RECT 17.4000 135.8000 17.8000 136.2000 ;
	    RECT 9.4000 135.1000 9.8000 135.2000 ;
	    RECT 10.2000 135.1000 10.6000 135.2000 ;
	    RECT 9.4000 134.8000 10.6000 135.1000 ;
	    RECT 11.8000 135.1000 12.2000 135.2000 ;
	    RECT 12.6000 135.1000 13.0000 135.2000 ;
	    RECT 11.8000 134.8000 13.0000 135.1000 ;
	    RECT 16.6000 134.8000 17.0000 135.2000 ;
	    RECT 16.6000 134.2000 16.9000 134.8000 ;
	    RECT 16.6000 133.8000 17.0000 134.2000 ;
	    RECT 17.4000 133.2000 17.7000 135.8000 ;
	    RECT 20.6000 135.1000 21.0000 135.2000 ;
	    RECT 21.4000 135.1000 21.8000 135.2000 ;
	    RECT 20.6000 134.8000 21.8000 135.1000 ;
	    RECT 22.2000 134.1000 22.5000 136.8000 ;
	    RECT 21.4000 133.8000 22.5000 134.1000 ;
	    RECT 9.4000 132.8000 9.8000 133.2000 ;
	    RECT 10.2000 132.8000 10.6000 133.2000 ;
	    RECT 17.4000 132.8000 17.8000 133.2000 ;
	    RECT 9.4000 131.1000 9.7000 132.8000 ;
	    RECT 8.6000 130.8000 9.7000 131.1000 ;
	    RECT 1.4000 128.8000 1.8000 129.2000 ;
	    RECT 3.8000 129.1000 4.2000 129.2000 ;
	    RECT 4.6000 129.1000 5.0000 129.2000 ;
	    RECT 3.8000 128.8000 5.0000 129.1000 ;
	    RECT 7.0000 128.8000 7.4000 129.2000 ;
	    RECT 7.8000 128.8000 8.2000 129.2000 ;
	    RECT 1.3000 127.5000 1.7000 127.9000 ;
	    RECT 4.6000 127.5000 5.0000 127.9000 ;
	    RECT 1.3000 125.1000 1.6000 127.5000 ;
	    RECT 4.7000 127.1000 5.0000 127.5000 ;
	    RECT 2.6000 126.8000 5.0000 127.1000 ;
	    RECT 7.0000 127.2000 7.3000 128.8000 ;
	    RECT 7.0000 126.8000 7.4000 127.2000 ;
	    RECT 2.6000 126.7000 3.0000 126.8000 ;
	    RECT 4.7000 125.1000 5.0000 126.8000 ;
	    RECT 8.6000 126.2000 8.9000 130.8000 ;
	    RECT 6.2000 126.1000 6.6000 126.2000 ;
	    RECT 7.0000 126.1000 7.4000 126.2000 ;
	    RECT 6.2000 125.8000 7.4000 126.1000 ;
	    RECT 8.6000 125.8000 9.0000 126.2000 ;
	    RECT 1.3000 124.7000 1.7000 125.1000 ;
	    RECT 4.6000 124.7000 5.0000 125.1000 ;
	    RECT 5.4000 114.1000 5.8000 114.2000 ;
	    RECT 6.2000 114.1000 6.6000 114.2000 ;
	    RECT 5.4000 113.8000 6.6000 114.1000 ;
	    RECT 3.0000 108.8000 3.4000 109.2000 ;
	    RECT 3.0000 108.2000 3.3000 108.8000 ;
	    RECT 5.4000 108.2000 5.7000 113.8000 ;
	    RECT 6.2000 111.8000 6.6000 112.2000 ;
	    RECT 3.0000 107.8000 3.4000 108.2000 ;
	    RECT 3.8000 107.8000 4.2000 108.2000 ;
	    RECT 5.4000 107.8000 5.8000 108.2000 ;
	    RECT 3.8000 107.2000 4.1000 107.8000 ;
	    RECT 0.6000 107.1000 1.0000 107.2000 ;
	    RECT 1.4000 107.1000 1.8000 107.2000 ;
	    RECT 0.6000 106.8000 1.8000 107.1000 ;
	    RECT 3.8000 106.8000 4.2000 107.2000 ;
	    RECT 4.6000 107.1000 5.0000 107.2000 ;
	    RECT 5.4000 107.1000 5.8000 107.2000 ;
	    RECT 4.6000 106.8000 5.8000 107.1000 ;
	    RECT 6.2000 106.2000 6.5000 111.8000 ;
	    RECT 10.2000 109.2000 10.5000 132.8000 ;
	    RECT 19.8000 130.8000 20.2000 131.2000 ;
	    RECT 14.1000 127.5000 14.5000 127.9000 ;
	    RECT 17.4000 127.5000 17.8000 127.9000 ;
	    RECT 14.1000 125.1000 14.4000 127.5000 ;
	    RECT 17.5000 127.1000 17.8000 127.5000 ;
	    RECT 15.4000 126.8000 17.8000 127.1000 ;
	    RECT 15.4000 126.7000 15.8000 126.8000 ;
	    RECT 16.6000 125.8000 17.0000 126.2000 ;
	    RECT 16.6000 125.2000 16.9000 125.8000 ;
	    RECT 14.1000 124.7000 14.5000 125.1000 ;
	    RECT 16.6000 124.8000 17.0000 125.2000 ;
	    RECT 17.5000 125.1000 17.8000 126.8000 ;
	    RECT 18.2000 126.1000 18.6000 126.2000 ;
	    RECT 19.0000 126.1000 19.4000 126.2000 ;
	    RECT 18.2000 125.8000 19.4000 126.1000 ;
	    RECT 17.4000 124.7000 17.8000 125.1000 ;
	    RECT 18.2000 122.8000 18.6000 123.2000 ;
	    RECT 18.2000 119.2000 18.5000 122.8000 ;
	    RECT 18.2000 118.8000 18.6000 119.2000 ;
	    RECT 12.6000 115.9000 13.0000 116.3000 ;
	    RECT 15.9000 115.9000 16.3000 116.3000 ;
	    RECT 11.0000 114.8000 11.4000 115.2000 ;
	    RECT 11.0000 114.2000 11.3000 114.8000 ;
	    RECT 12.6000 114.2000 12.9000 115.9000 ;
	    RECT 14.6000 114.2000 15.0000 114.3000 ;
	    RECT 11.0000 113.8000 11.4000 114.2000 ;
	    RECT 12.6000 113.9000 15.0000 114.2000 ;
	    RECT 12.6000 113.5000 12.9000 113.9000 ;
	    RECT 16.0000 113.5000 16.3000 115.9000 ;
	    RECT 19.8000 116.2000 20.1000 130.8000 ;
	    RECT 21.4000 127.2000 21.7000 133.8000 ;
	    RECT 22.2000 129.8000 22.6000 130.2000 ;
	    RECT 21.4000 126.8000 21.8000 127.2000 ;
	    RECT 21.4000 125.2000 21.7000 126.8000 ;
	    RECT 21.4000 124.8000 21.8000 125.2000 ;
	    RECT 22.2000 116.2000 22.5000 129.8000 ;
	    RECT 23.0000 129.2000 23.3000 144.8000 ;
	    RECT 23.8000 135.2000 24.1000 145.8000 ;
	    RECT 26.2000 141.8000 26.6000 142.2000 ;
	    RECT 26.2000 139.2000 26.5000 141.8000 ;
	    RECT 26.2000 138.8000 26.6000 139.2000 ;
	    RECT 27.0000 137.2000 27.3000 145.8000 ;
	    RECT 30.2000 145.1000 30.6000 147.9000 ;
	    RECT 31.8000 143.1000 32.2000 148.9000 ;
	    RECT 32.6000 145.9000 33.0000 146.3000 ;
	    RECT 29.4000 141.8000 29.8000 142.2000 ;
	    RECT 28.6000 137.8000 29.0000 138.2000 ;
	    RECT 25.4000 136.8000 25.8000 137.2000 ;
	    RECT 27.0000 136.8000 27.4000 137.2000 ;
	    RECT 23.8000 134.8000 24.2000 135.2000 ;
	    RECT 25.4000 133.2000 25.7000 136.8000 ;
	    RECT 27.0000 135.1000 27.4000 135.2000 ;
	    RECT 27.8000 135.1000 28.2000 135.2000 ;
	    RECT 27.0000 134.8000 28.2000 135.1000 ;
	    RECT 28.6000 134.2000 28.9000 137.8000 ;
	    RECT 29.4000 136.2000 29.7000 141.8000 ;
	    RECT 31.0000 137.8000 31.4000 138.2000 ;
	    RECT 31.0000 136.2000 31.3000 137.8000 ;
	    RECT 29.4000 135.8000 29.8000 136.2000 ;
	    RECT 31.0000 135.8000 31.4000 136.2000 ;
	    RECT 29.4000 134.8000 29.8000 135.2000 ;
	    RECT 29.4000 134.2000 29.7000 134.8000 ;
	    RECT 28.6000 133.8000 29.0000 134.2000 ;
	    RECT 29.4000 133.8000 29.8000 134.2000 ;
	    RECT 31.8000 133.8000 32.2000 134.2000 ;
	    RECT 31.8000 133.2000 32.1000 133.8000 ;
	    RECT 25.4000 132.8000 25.8000 133.2000 ;
	    RECT 31.8000 132.8000 32.2000 133.2000 ;
	    RECT 24.6000 131.8000 25.0000 132.2000 ;
	    RECT 26.2000 131.8000 26.6000 132.2000 ;
	    RECT 30.2000 131.8000 30.6000 132.2000 ;
	    RECT 24.6000 130.2000 24.9000 131.8000 ;
	    RECT 26.2000 131.2000 26.5000 131.8000 ;
	    RECT 26.2000 130.8000 26.6000 131.2000 ;
	    RECT 24.6000 129.8000 25.0000 130.2000 ;
	    RECT 23.0000 128.8000 23.4000 129.2000 ;
	    RECT 23.8000 128.8000 24.2000 129.2000 ;
	    RECT 23.8000 128.2000 24.1000 128.8000 ;
	    RECT 30.2000 128.2000 30.5000 131.8000 ;
	    RECT 32.6000 129.2000 32.9000 145.9000 ;
	    RECT 35.8000 145.8000 36.2000 146.2000 ;
	    RECT 35.8000 144.2000 36.1000 145.8000 ;
	    RECT 35.8000 143.8000 36.2000 144.2000 ;
	    RECT 36.6000 143.1000 37.0000 148.9000 ;
	    RECT 43.8000 148.8000 44.2000 149.2000 ;
	    RECT 51.0000 149.1000 51.4000 149.2000 ;
	    RECT 51.8000 149.1000 52.2000 149.2000 ;
	    RECT 51.0000 148.8000 52.2000 149.1000 ;
	    RECT 43.8000 148.2000 44.1000 148.8000 ;
	    RECT 43.8000 147.8000 44.2000 148.2000 ;
	    RECT 46.2000 147.8000 46.6000 148.2000 ;
	    RECT 50.2000 148.1000 50.6000 148.2000 ;
	    RECT 51.0000 148.1000 51.4000 148.2000 ;
	    RECT 50.2000 147.8000 51.4000 148.1000 ;
	    RECT 43.8000 146.8000 44.2000 147.2000 ;
	    RECT 43.8000 146.2000 44.1000 146.8000 ;
	    RECT 42.2000 145.8000 42.6000 146.2000 ;
	    RECT 43.8000 145.8000 44.2000 146.2000 ;
	    RECT 40.6000 143.8000 41.0000 144.2000 ;
	    RECT 39.0000 141.8000 39.4000 142.2000 ;
	    RECT 39.0000 141.2000 39.3000 141.8000 ;
	    RECT 39.0000 140.8000 39.4000 141.2000 ;
	    RECT 34.2000 138.8000 34.6000 139.2000 ;
	    RECT 34.2000 136.2000 34.5000 138.8000 ;
	    RECT 33.4000 135.8000 33.8000 136.2000 ;
	    RECT 34.2000 135.8000 34.6000 136.2000 ;
	    RECT 32.6000 128.8000 33.0000 129.2000 ;
	    RECT 23.8000 127.8000 24.2000 128.2000 ;
	    RECT 26.2000 127.8000 26.6000 128.2000 ;
	    RECT 28.6000 127.8000 29.0000 128.2000 ;
	    RECT 30.2000 127.8000 30.6000 128.2000 ;
	    RECT 32.6000 127.8000 33.0000 128.2000 ;
	    RECT 26.2000 127.2000 26.5000 127.8000 ;
	    RECT 28.6000 127.2000 28.9000 127.8000 ;
	    RECT 32.6000 127.2000 32.9000 127.8000 ;
	    RECT 26.2000 126.8000 26.6000 127.2000 ;
	    RECT 28.6000 126.8000 29.0000 127.2000 ;
	    RECT 30.2000 126.8000 30.6000 127.2000 ;
	    RECT 31.0000 126.8000 31.4000 127.2000 ;
	    RECT 32.6000 126.8000 33.0000 127.2000 ;
	    RECT 30.2000 126.2000 30.5000 126.8000 ;
	    RECT 27.8000 125.8000 28.2000 126.2000 ;
	    RECT 30.2000 125.8000 30.6000 126.2000 ;
	    RECT 27.0000 124.8000 27.4000 125.2000 ;
	    RECT 23.8000 123.8000 24.2000 124.2000 ;
	    RECT 19.8000 115.8000 20.2000 116.2000 ;
	    RECT 22.2000 115.8000 22.6000 116.2000 ;
	    RECT 18.2000 114.8000 18.6000 115.2000 ;
	    RECT 20.6000 114.8000 21.0000 115.2000 ;
	    RECT 12.6000 113.1000 13.0000 113.5000 ;
	    RECT 15.9000 113.1000 16.3000 113.5000 ;
	    RECT 17.4000 113.8000 17.8000 114.2000 ;
	    RECT 17.4000 113.2000 17.7000 113.8000 ;
	    RECT 17.4000 112.8000 17.8000 113.2000 ;
	    RECT 13.4000 111.8000 13.8000 112.2000 ;
	    RECT 13.4000 109.2000 13.7000 111.8000 ;
	    RECT 18.2000 109.2000 18.5000 114.8000 ;
	    RECT 20.6000 114.2000 20.9000 114.8000 ;
	    RECT 22.2000 114.2000 22.5000 115.8000 ;
	    RECT 23.8000 115.2000 24.1000 123.8000 ;
	    RECT 27.0000 119.2000 27.3000 124.8000 ;
	    RECT 27.0000 118.8000 27.4000 119.2000 ;
	    RECT 23.8000 114.8000 24.2000 115.2000 ;
	    RECT 27.0000 114.8000 27.4000 115.2000 ;
	    RECT 27.0000 114.2000 27.3000 114.8000 ;
	    RECT 20.6000 113.8000 21.0000 114.2000 ;
	    RECT 21.4000 113.8000 21.8000 114.2000 ;
	    RECT 22.2000 113.8000 22.6000 114.2000 ;
	    RECT 26.2000 113.8000 26.6000 114.2000 ;
	    RECT 27.0000 113.8000 27.4000 114.2000 ;
	    RECT 21.4000 113.2000 21.7000 113.8000 ;
	    RECT 26.2000 113.2000 26.5000 113.8000 ;
	    RECT 21.4000 112.8000 21.8000 113.2000 ;
	    RECT 26.2000 112.8000 26.6000 113.2000 ;
	    RECT 27.8000 112.2000 28.1000 125.8000 ;
	    RECT 31.0000 125.2000 31.3000 126.8000 ;
	    RECT 31.8000 125.8000 32.2000 126.2000 ;
	    RECT 31.0000 124.8000 31.4000 125.2000 ;
	    RECT 30.2000 117.8000 30.6000 118.2000 ;
	    RECT 30.2000 117.2000 30.5000 117.8000 ;
	    RECT 30.2000 116.8000 30.6000 117.2000 ;
	    RECT 28.6000 116.1000 29.0000 116.2000 ;
	    RECT 29.4000 116.1000 29.8000 116.2000 ;
	    RECT 28.6000 115.8000 29.8000 116.1000 ;
	    RECT 31.0000 116.1000 31.3000 124.8000 ;
	    RECT 31.8000 123.2000 32.1000 125.8000 ;
	    RECT 31.8000 122.8000 32.2000 123.2000 ;
	    RECT 33.4000 116.2000 33.7000 135.8000 ;
	    RECT 34.2000 128.2000 34.5000 135.8000 ;
	    RECT 35.8000 135.1000 36.2000 135.2000 ;
	    RECT 36.6000 135.1000 37.0000 135.2000 ;
	    RECT 35.8000 134.8000 37.0000 135.1000 ;
	    RECT 37.4000 133.8000 37.8000 134.2000 ;
	    RECT 39.0000 133.8000 39.4000 134.2000 ;
	    RECT 34.2000 127.8000 34.6000 128.2000 ;
	    RECT 35.0000 127.8000 35.4000 128.2000 ;
	    RECT 35.8000 127.8000 36.2000 128.2000 ;
	    RECT 34.2000 126.8000 34.6000 127.2000 ;
	    RECT 34.2000 126.2000 34.5000 126.8000 ;
	    RECT 35.0000 126.2000 35.3000 127.8000 ;
	    RECT 35.8000 127.2000 36.1000 127.8000 ;
	    RECT 37.4000 127.2000 37.7000 133.8000 ;
	    RECT 39.0000 133.2000 39.3000 133.8000 ;
	    RECT 39.0000 132.8000 39.4000 133.2000 ;
	    RECT 39.8000 133.1000 40.2000 135.9000 ;
	    RECT 40.6000 134.2000 40.9000 143.8000 ;
	    RECT 40.6000 133.8000 41.0000 134.2000 ;
	    RECT 41.4000 132.1000 41.8000 137.9000 ;
	    RECT 42.2000 137.1000 42.5000 145.8000 ;
	    RECT 46.2000 144.2000 46.5000 147.8000 ;
	    RECT 50.2000 146.1000 50.6000 146.2000 ;
	    RECT 51.0000 146.1000 51.4000 146.2000 ;
	    RECT 50.2000 145.8000 51.4000 146.1000 ;
	    RECT 53.4000 145.2000 53.7000 149.8000 ;
	    RECT 60.6000 148.2000 60.9000 151.8000 ;
	    RECT 57.4000 147.8000 57.8000 148.2000 ;
	    RECT 60.6000 147.8000 61.0000 148.2000 ;
	    RECT 57.4000 147.2000 57.7000 147.8000 ;
	    RECT 61.4000 147.2000 61.7000 163.8000 ;
	    RECT 62.2000 153.1000 62.6000 155.9000 ;
	    RECT 63.0000 154.8000 63.4000 155.2000 ;
	    RECT 63.0000 149.2000 63.3000 154.8000 ;
	    RECT 63.8000 152.1000 64.2000 157.9000 ;
	    RECT 64.6000 155.8000 65.0000 156.2000 ;
	    RECT 64.6000 155.1000 64.9000 155.8000 ;
	    RECT 64.6000 154.7000 65.0000 155.1000 ;
	    RECT 66.2000 154.2000 66.5000 173.8000 ;
	    RECT 67.8000 169.2000 68.1000 174.8000 ;
	    RECT 69.4000 172.1000 69.8000 177.9000 ;
	    RECT 75.0000 174.8000 75.4000 175.2000 ;
	    RECT 77.4000 174.8000 77.8000 175.2000 ;
	    RECT 71.8000 172.1000 72.2000 172.2000 ;
	    RECT 71.0000 171.8000 72.2000 172.1000 ;
	    RECT 67.8000 168.8000 68.2000 169.2000 ;
	    RECT 71.0000 168.2000 71.3000 171.8000 ;
	    RECT 67.0000 168.1000 67.4000 168.2000 ;
	    RECT 67.8000 168.1000 68.2000 168.2000 ;
	    RECT 67.0000 167.8000 68.2000 168.1000 ;
	    RECT 71.0000 167.8000 71.4000 168.2000 ;
	    RECT 71.8000 168.1000 72.2000 168.2000 ;
	    RECT 72.6000 168.1000 73.0000 168.2000 ;
	    RECT 71.8000 167.8000 73.0000 168.1000 ;
	    RECT 65.4000 153.8000 65.8000 154.2000 ;
	    RECT 66.2000 153.8000 66.6000 154.2000 ;
	    RECT 63.0000 148.8000 63.4000 149.2000 ;
	    RECT 63.0000 148.1000 63.4000 148.2000 ;
	    RECT 63.8000 148.1000 64.2000 148.2000 ;
	    RECT 63.0000 147.8000 64.2000 148.1000 ;
	    RECT 57.4000 146.8000 57.8000 147.2000 ;
	    RECT 61.4000 146.8000 61.8000 147.2000 ;
	    RECT 63.0000 146.8000 63.4000 147.2000 ;
	    RECT 55.0000 145.8000 55.4000 146.2000 ;
	    RECT 55.8000 145.8000 56.2000 146.2000 ;
	    RECT 53.4000 145.1000 53.8000 145.2000 ;
	    RECT 54.2000 145.1000 54.6000 145.2000 ;
	    RECT 53.4000 144.8000 54.6000 145.1000 ;
	    RECT 55.0000 144.2000 55.3000 145.8000 ;
	    RECT 46.2000 143.8000 46.6000 144.2000 ;
	    RECT 55.0000 143.8000 55.4000 144.2000 ;
	    RECT 55.8000 139.2000 56.1000 145.8000 ;
	    RECT 62.2000 143.8000 62.6000 144.2000 ;
	    RECT 62.2000 139.2000 62.5000 143.8000 ;
	    RECT 55.8000 138.8000 56.2000 139.2000 ;
	    RECT 62.2000 138.8000 62.6000 139.2000 ;
	    RECT 42.2000 136.8000 43.3000 137.1000 ;
	    RECT 42.2000 135.8000 42.6000 136.2000 ;
	    RECT 42.2000 135.1000 42.5000 135.8000 ;
	    RECT 42.2000 134.7000 42.6000 135.1000 ;
	    RECT 39.0000 130.8000 39.4000 131.2000 ;
	    RECT 38.2000 128.8000 38.6000 129.2000 ;
	    RECT 38.2000 128.2000 38.5000 128.8000 ;
	    RECT 38.2000 127.8000 38.6000 128.2000 ;
	    RECT 39.0000 127.2000 39.3000 130.8000 ;
	    RECT 42.2000 128.8000 42.6000 129.2000 ;
	    RECT 42.2000 127.2000 42.5000 128.8000 ;
	    RECT 35.8000 126.8000 36.2000 127.2000 ;
	    RECT 37.4000 126.8000 37.8000 127.2000 ;
	    RECT 39.0000 126.8000 39.4000 127.2000 ;
	    RECT 42.2000 126.8000 42.6000 127.2000 ;
	    RECT 34.2000 125.8000 34.6000 126.2000 ;
	    RECT 35.0000 125.8000 35.4000 126.2000 ;
	    RECT 39.0000 125.1000 39.4000 125.2000 ;
	    RECT 39.8000 125.1000 40.2000 125.2000 ;
	    RECT 39.0000 124.8000 40.2000 125.1000 ;
	    RECT 41.4000 124.8000 41.8000 125.2000 ;
	    RECT 41.4000 124.2000 41.7000 124.8000 ;
	    RECT 41.4000 123.8000 41.8000 124.2000 ;
	    RECT 35.0000 122.8000 35.4000 123.2000 ;
	    RECT 35.0000 117.2000 35.3000 122.8000 ;
	    RECT 43.0000 122.2000 43.3000 136.8000 ;
	    RECT 45.4000 134.8000 45.8000 135.2000 ;
	    RECT 43.8000 127.8000 44.2000 128.2000 ;
	    RECT 43.8000 127.2000 44.1000 127.8000 ;
	    RECT 43.8000 126.8000 44.2000 127.2000 ;
	    RECT 44.6000 125.1000 45.0000 127.9000 ;
	    RECT 45.4000 127.2000 45.7000 134.8000 ;
	    RECT 46.2000 132.1000 46.6000 137.9000 ;
	    RECT 50.2000 136.8000 50.6000 137.2000 ;
	    RECT 50.2000 136.2000 50.5000 136.8000 ;
	    RECT 50.2000 135.8000 50.6000 136.2000 ;
	    RECT 55.8000 135.8000 56.2000 136.2000 ;
	    RECT 55.8000 135.2000 56.1000 135.8000 ;
	    RECT 51.0000 134.8000 51.4000 135.2000 ;
	    RECT 51.8000 134.8000 52.2000 135.2000 ;
	    RECT 55.8000 134.8000 56.2000 135.2000 ;
	    RECT 57.4000 134.8000 57.8000 135.2000 ;
	    RECT 51.0000 133.2000 51.3000 134.8000 ;
	    RECT 51.8000 134.2000 52.1000 134.8000 ;
	    RECT 51.8000 133.8000 52.2000 134.2000 ;
	    RECT 52.6000 134.0000 53.0000 134.4000 ;
	    RECT 52.6000 133.2000 52.9000 134.0000 ;
	    RECT 48.6000 132.8000 49.0000 133.2000 ;
	    RECT 51.0000 132.8000 51.4000 133.2000 ;
	    RECT 52.6000 132.8000 53.0000 133.2000 ;
	    RECT 48.6000 132.2000 48.9000 132.8000 ;
	    RECT 48.6000 131.8000 49.0000 132.2000 ;
	    RECT 45.4000 126.8000 45.8000 127.2000 ;
	    RECT 46.2000 123.1000 46.6000 128.9000 ;
	    RECT 49.4000 128.8000 49.8000 129.2000 ;
	    RECT 47.0000 125.9000 47.4000 126.3000 ;
	    RECT 47.0000 125.2000 47.3000 125.9000 ;
	    RECT 47.0000 124.8000 47.4000 125.2000 ;
	    RECT 48.6000 123.8000 49.0000 124.2000 ;
	    RECT 43.0000 121.8000 43.4000 122.2000 ;
	    RECT 46.2000 121.8000 46.6000 122.2000 ;
	    RECT 35.0000 116.8000 35.4000 117.2000 ;
	    RECT 31.8000 116.1000 32.2000 116.2000 ;
	    RECT 31.0000 115.8000 32.2000 116.1000 ;
	    RECT 33.4000 115.8000 33.8000 116.2000 ;
	    RECT 30.2000 115.1000 30.6000 115.2000 ;
	    RECT 31.0000 115.1000 31.4000 115.2000 ;
	    RECT 30.2000 114.8000 31.4000 115.1000 ;
	    RECT 31.8000 114.8000 32.2000 115.2000 ;
	    RECT 28.6000 114.1000 29.0000 114.2000 ;
	    RECT 29.4000 114.1000 29.8000 114.2000 ;
	    RECT 28.6000 113.8000 29.8000 114.1000 ;
	    RECT 25.4000 111.8000 25.8000 112.2000 ;
	    RECT 27.8000 111.8000 28.2000 112.2000 ;
	    RECT 10.2000 108.8000 10.6000 109.2000 ;
	    RECT 11.0000 108.8000 11.4000 109.2000 ;
	    RECT 13.4000 108.8000 13.8000 109.2000 ;
	    RECT 18.2000 108.8000 18.6000 109.2000 ;
	    RECT 11.0000 108.2000 11.3000 108.8000 ;
	    RECT 7.8000 107.8000 8.2000 108.2000 ;
	    RECT 11.0000 107.8000 11.4000 108.2000 ;
	    RECT 1.4000 106.1000 1.8000 106.2000 ;
	    RECT 1.4000 105.8000 2.5000 106.1000 ;
	    RECT 6.2000 105.8000 6.6000 106.2000 ;
	    RECT 0.6000 96.1000 1.0000 96.2000 ;
	    RECT 1.4000 96.1000 1.8000 96.2000 ;
	    RECT 0.6000 95.8000 1.8000 96.1000 ;
	    RECT 2.2000 85.2000 2.5000 105.8000 ;
	    RECT 3.0000 105.1000 3.4000 105.2000 ;
	    RECT 3.8000 105.1000 4.2000 105.2000 ;
	    RECT 3.0000 104.8000 4.2000 105.1000 ;
	    RECT 5.4000 105.1000 5.8000 105.2000 ;
	    RECT 6.2000 105.1000 6.6000 105.2000 ;
	    RECT 5.4000 104.8000 6.6000 105.1000 ;
	    RECT 7.8000 104.2000 8.1000 107.8000 ;
	    RECT 15.0000 107.5000 15.4000 107.9000 ;
	    RECT 18.3000 107.5000 18.7000 107.9000 ;
	    RECT 8.6000 106.8000 9.0000 107.2000 ;
	    RECT 9.4000 106.8000 9.8000 107.2000 ;
	    RECT 11.0000 107.1000 11.4000 107.2000 ;
	    RECT 11.8000 107.1000 12.2000 107.2000 ;
	    RECT 11.0000 106.8000 12.2000 107.1000 ;
	    RECT 15.0000 107.1000 15.3000 107.5000 ;
	    RECT 15.0000 106.8000 17.4000 107.1000 ;
	    RECT 8.6000 106.2000 8.9000 106.8000 ;
	    RECT 9.4000 106.2000 9.7000 106.8000 ;
	    RECT 8.6000 105.8000 9.0000 106.2000 ;
	    RECT 9.4000 105.8000 9.8000 106.2000 ;
	    RECT 13.4000 104.8000 13.8000 105.2000 ;
	    RECT 15.0000 105.1000 15.3000 106.8000 ;
	    RECT 17.0000 106.7000 17.4000 106.8000 ;
	    RECT 15.8000 105.8000 16.2000 106.2000 ;
	    RECT 15.8000 105.2000 16.1000 105.8000 ;
	    RECT 13.4000 104.2000 13.7000 104.8000 ;
	    RECT 15.0000 104.7000 15.4000 105.1000 ;
	    RECT 15.8000 104.8000 16.2000 105.2000 ;
	    RECT 18.4000 105.1000 18.7000 107.5000 ;
	    RECT 21.4000 106.8000 21.8000 107.2000 ;
	    RECT 21.4000 106.2000 21.7000 106.8000 ;
	    RECT 21.4000 105.8000 21.8000 106.2000 ;
	    RECT 22.2000 106.1000 22.6000 106.2000 ;
	    RECT 23.0000 106.1000 23.4000 106.2000 ;
	    RECT 22.2000 105.8000 23.4000 106.1000 ;
	    RECT 18.3000 104.7000 18.7000 105.1000 ;
	    RECT 7.8000 103.8000 8.2000 104.2000 ;
	    RECT 12.6000 103.8000 13.0000 104.2000 ;
	    RECT 13.4000 103.8000 13.8000 104.2000 ;
	    RECT 23.8000 104.1000 24.2000 104.2000 ;
	    RECT 24.6000 104.1000 25.0000 104.2000 ;
	    RECT 23.8000 103.8000 25.0000 104.1000 ;
	    RECT 12.6000 99.2000 12.9000 103.8000 ;
	    RECT 23.8000 102.8000 24.2000 103.2000 ;
	    RECT 23.0000 101.8000 23.4000 102.2000 ;
	    RECT 12.6000 98.8000 13.0000 99.2000 ;
	    RECT 11.0000 95.8000 11.4000 96.2000 ;
	    RECT 11.8000 95.8000 12.2000 96.2000 ;
	    RECT 18.2000 95.9000 18.6000 96.3000 ;
	    RECT 21.3000 95.9000 21.7000 96.3000 ;
	    RECT 11.0000 95.2000 11.3000 95.8000 ;
	    RECT 11.8000 95.2000 12.1000 95.8000 ;
	    RECT 9.4000 94.8000 9.8000 95.2000 ;
	    RECT 11.0000 94.8000 11.4000 95.2000 ;
	    RECT 11.8000 94.8000 12.2000 95.2000 ;
	    RECT 14.2000 95.1000 14.6000 95.2000 ;
	    RECT 15.0000 95.1000 15.4000 95.2000 ;
	    RECT 14.2000 94.8000 15.4000 95.1000 ;
	    RECT 9.4000 94.2000 9.7000 94.8000 ;
	    RECT 18.2000 94.2000 18.5000 95.9000 ;
	    RECT 20.7000 94.9000 21.1000 95.3000 ;
	    RECT 20.7000 94.2000 21.0000 94.9000 ;
	    RECT 9.4000 93.8000 9.8000 94.2000 ;
	    RECT 13.4000 93.8000 13.8000 94.2000 ;
	    RECT 18.2000 93.9000 21.0000 94.2000 ;
	    RECT 13.4000 93.2000 13.7000 93.8000 ;
	    RECT 18.2000 93.5000 18.5000 93.9000 ;
	    RECT 18.9000 93.5000 19.3000 93.6000 ;
	    RECT 20.6000 93.5000 21.0000 93.6000 ;
	    RECT 21.4000 93.5000 21.7000 95.9000 ;
	    RECT 23.0000 96.2000 23.3000 101.8000 ;
	    RECT 23.8000 99.2000 24.1000 102.8000 ;
	    RECT 23.8000 98.8000 24.2000 99.2000 ;
	    RECT 25.4000 96.2000 25.7000 111.8000 ;
	    RECT 26.2000 103.1000 26.6000 108.9000 ;
	    RECT 30.2000 108.8000 30.6000 109.2000 ;
	    RECT 30.2000 108.2000 30.5000 108.8000 ;
	    RECT 30.2000 107.8000 30.6000 108.2000 ;
	    RECT 30.2000 106.8000 30.6000 107.2000 ;
	    RECT 30.2000 106.3000 30.5000 106.8000 ;
	    RECT 30.2000 105.9000 30.6000 106.3000 ;
	    RECT 31.0000 103.1000 31.4000 108.9000 ;
	    RECT 31.8000 103.2000 32.1000 114.8000 ;
	    RECT 33.4000 114.2000 33.7000 115.8000 ;
	    RECT 34.2000 114.8000 34.6000 115.2000 ;
	    RECT 34.2000 114.2000 34.5000 114.8000 ;
	    RECT 35.0000 114.2000 35.3000 116.8000 ;
	    RECT 35.8000 114.8000 36.2000 115.2000 ;
	    RECT 35.8000 114.2000 36.1000 114.8000 ;
	    RECT 33.4000 113.8000 33.8000 114.2000 ;
	    RECT 34.2000 113.8000 34.6000 114.2000 ;
	    RECT 35.0000 113.8000 35.4000 114.2000 ;
	    RECT 35.8000 113.8000 36.2000 114.2000 ;
	    RECT 36.6000 113.1000 37.0000 115.9000 ;
	    RECT 37.4000 113.8000 37.8000 114.2000 ;
	    RECT 36.6000 110.8000 37.0000 111.2000 ;
	    RECT 32.6000 105.1000 33.0000 107.9000 ;
	    RECT 33.4000 107.8000 33.8000 108.2000 ;
	    RECT 33.4000 104.2000 33.7000 107.8000 ;
	    RECT 35.0000 106.8000 35.4000 107.2000 ;
	    RECT 35.0000 106.2000 35.3000 106.8000 ;
	    RECT 36.6000 106.2000 36.9000 110.8000 ;
	    RECT 37.4000 108.2000 37.7000 113.8000 ;
	    RECT 38.2000 112.1000 38.6000 117.9000 ;
	    RECT 42.2000 116.8000 42.6000 117.2000 ;
	    RECT 39.0000 115.8000 39.4000 116.2000 ;
	    RECT 39.0000 115.1000 39.3000 115.8000 ;
	    RECT 42.2000 115.2000 42.5000 116.8000 ;
	    RECT 39.0000 114.7000 39.4000 115.1000 ;
	    RECT 42.2000 114.8000 42.6000 115.2000 ;
	    RECT 43.0000 112.1000 43.4000 117.9000 ;
	    RECT 46.2000 117.2000 46.5000 121.8000 ;
	    RECT 46.2000 116.8000 46.6000 117.2000 ;
	    RECT 46.2000 114.2000 46.5000 116.8000 ;
	    RECT 46.2000 113.8000 46.6000 114.2000 ;
	    RECT 47.0000 114.1000 47.4000 114.2000 ;
	    RECT 47.8000 114.1000 48.2000 114.2000 ;
	    RECT 47.0000 113.8000 48.2000 114.1000 ;
	    RECT 41.4000 109.1000 41.8000 109.2000 ;
	    RECT 42.2000 109.1000 42.6000 109.2000 ;
	    RECT 41.4000 108.8000 42.6000 109.1000 ;
	    RECT 48.6000 108.2000 48.9000 123.8000 ;
	    RECT 49.4000 113.2000 49.7000 128.8000 ;
	    RECT 50.2000 125.8000 50.6000 126.2000 ;
	    RECT 50.2000 117.2000 50.5000 125.8000 ;
	    RECT 51.0000 123.1000 51.4000 128.9000 ;
	    RECT 52.6000 128.2000 52.9000 132.8000 ;
	    RECT 57.4000 129.2000 57.7000 134.8000 ;
	    RECT 58.2000 133.8000 58.6000 134.2000 ;
	    RECT 58.2000 132.2000 58.5000 133.8000 ;
	    RECT 60.6000 132.8000 61.0000 133.2000 ;
	    RECT 58.2000 131.8000 58.6000 132.2000 ;
	    RECT 53.4000 128.8000 53.8000 129.2000 ;
	    RECT 57.4000 128.8000 57.8000 129.2000 ;
	    RECT 53.4000 128.2000 53.7000 128.8000 ;
	    RECT 52.6000 127.8000 53.0000 128.2000 ;
	    RECT 53.4000 127.8000 53.8000 128.2000 ;
	    RECT 54.2000 126.8000 54.6000 127.2000 ;
	    RECT 54.2000 126.2000 54.5000 126.8000 ;
	    RECT 54.2000 125.8000 54.6000 126.2000 ;
	    RECT 55.0000 126.1000 55.4000 126.2000 ;
	    RECT 55.8000 126.1000 56.2000 126.2000 ;
	    RECT 55.0000 125.8000 56.2000 126.1000 ;
	    RECT 57.4000 126.1000 57.8000 126.2000 ;
	    RECT 58.2000 126.1000 58.6000 126.2000 ;
	    RECT 57.4000 125.8000 58.6000 126.1000 ;
	    RECT 60.6000 122.2000 60.9000 132.8000 ;
	    RECT 62.2000 132.1000 62.6000 132.2000 ;
	    RECT 61.4000 131.8000 62.6000 132.1000 ;
	    RECT 61.4000 127.2000 61.7000 131.8000 ;
	    RECT 62.2000 128.8000 62.6000 129.2000 ;
	    RECT 62.2000 128.2000 62.5000 128.8000 ;
	    RECT 63.0000 128.2000 63.3000 146.8000 ;
	    RECT 64.6000 145.1000 65.0000 147.9000 ;
	    RECT 65.4000 147.2000 65.7000 153.8000 ;
	    RECT 65.4000 146.8000 65.8000 147.2000 ;
	    RECT 66.2000 143.1000 66.6000 148.9000 ;
	    RECT 67.0000 148.2000 67.3000 167.8000 ;
	    RECT 68.6000 166.8000 69.0000 167.2000 ;
	    RECT 73.4000 166.8000 73.8000 167.2000 ;
	    RECT 68.6000 164.2000 68.9000 166.8000 ;
	    RECT 71.8000 166.1000 72.2000 166.2000 ;
	    RECT 72.6000 166.1000 73.0000 166.2000 ;
	    RECT 71.8000 165.8000 73.0000 166.1000 ;
	    RECT 72.6000 164.8000 73.0000 165.2000 ;
	    RECT 68.6000 163.8000 69.0000 164.2000 ;
	    RECT 71.0000 161.8000 71.4000 162.2000 ;
	    RECT 71.0000 159.2000 71.3000 161.8000 ;
	    RECT 72.6000 159.2000 72.9000 164.8000 ;
	    RECT 73.4000 164.2000 73.7000 166.8000 ;
	    RECT 73.4000 163.8000 73.8000 164.2000 ;
	    RECT 75.0000 162.2000 75.3000 174.8000 ;
	    RECT 77.4000 167.2000 77.7000 174.8000 ;
	    RECT 79.8000 173.1000 80.2000 175.9000 ;
	    RECT 81.4000 172.1000 81.8000 177.9000 ;
	    RECT 83.0000 175.1000 83.4000 175.2000 ;
	    RECT 83.8000 175.1000 84.2000 175.2000 ;
	    RECT 83.0000 174.8000 84.2000 175.1000 ;
	    RECT 82.2000 172.8000 82.6000 173.2000 ;
	    RECT 77.4000 166.8000 77.8000 167.2000 ;
	    RECT 79.0000 163.1000 79.4000 168.9000 ;
	    RECT 82.2000 167.2000 82.5000 172.8000 ;
	    RECT 86.2000 172.1000 86.6000 177.9000 ;
	    RECT 89.4000 176.8000 89.8000 177.2000 ;
	    RECT 89.4000 176.2000 89.7000 176.8000 ;
	    RECT 89.4000 175.8000 89.8000 176.2000 ;
	    RECT 93.4000 175.8000 93.8000 176.2000 ;
	    RECT 93.4000 175.2000 93.7000 175.8000 ;
	    RECT 91.0000 174.8000 91.4000 175.2000 ;
	    RECT 91.8000 175.1000 92.2000 175.2000 ;
	    RECT 92.6000 175.1000 93.0000 175.2000 ;
	    RECT 91.8000 174.8000 93.0000 175.1000 ;
	    RECT 93.4000 174.8000 93.8000 175.2000 ;
	    RECT 95.8000 174.8000 96.2000 175.2000 ;
	    RECT 91.0000 174.2000 91.3000 174.8000 ;
	    RECT 91.0000 173.8000 91.4000 174.2000 ;
	    RECT 91.8000 173.8000 92.2000 174.2000 ;
	    RECT 82.2000 166.8000 82.6000 167.2000 ;
	    RECT 80.6000 166.1000 81.0000 166.2000 ;
	    RECT 81.4000 166.1000 81.8000 166.2000 ;
	    RECT 80.6000 165.8000 81.8000 166.1000 ;
	    RECT 82.2000 165.8000 82.6000 166.2000 ;
	    RECT 75.0000 161.8000 75.4000 162.2000 ;
	    RECT 82.2000 159.2000 82.5000 165.8000 ;
	    RECT 83.8000 163.1000 84.2000 168.9000 ;
	    RECT 85.4000 165.1000 85.8000 167.9000 ;
	    RECT 86.2000 165.1000 86.6000 167.9000 ;
	    RECT 84.6000 163.8000 85.0000 164.2000 ;
	    RECT 71.0000 158.8000 71.4000 159.2000 ;
	    RECT 72.6000 158.8000 73.0000 159.2000 ;
	    RECT 82.2000 158.8000 82.6000 159.2000 ;
	    RECT 68.6000 152.1000 69.0000 157.9000 ;
	    RECT 84.6000 156.2000 84.9000 163.8000 ;
	    RECT 87.8000 163.1000 88.2000 168.9000 ;
	    RECT 88.6000 167.8000 89.0000 168.2000 ;
	    RECT 88.6000 162.2000 88.9000 167.8000 ;
	    RECT 89.4000 166.8000 89.8000 167.2000 ;
	    RECT 89.4000 166.2000 89.7000 166.8000 ;
	    RECT 91.8000 166.2000 92.1000 173.8000 ;
	    RECT 89.4000 165.8000 89.8000 166.2000 ;
	    RECT 91.8000 165.8000 92.2000 166.2000 ;
	    RECT 91.0000 164.8000 91.4000 165.2000 ;
	    RECT 88.6000 161.8000 89.0000 162.2000 ;
	    RECT 88.6000 159.2000 88.9000 161.8000 ;
	    RECT 91.0000 159.2000 91.3000 164.8000 ;
	    RECT 88.6000 158.8000 89.0000 159.2000 ;
	    RECT 91.0000 158.8000 91.4000 159.2000 ;
	    RECT 84.6000 155.8000 85.0000 156.2000 ;
	    RECT 75.0000 154.8000 75.4000 155.2000 ;
	    RECT 83.8000 154.8000 84.2000 155.2000 ;
	    RECT 75.0000 153.2000 75.3000 154.8000 ;
	    RECT 77.4000 153.8000 77.8000 154.2000 ;
	    RECT 78.2000 153.8000 78.6000 154.2000 ;
	    RECT 77.4000 153.2000 77.7000 153.8000 ;
	    RECT 75.0000 153.1000 75.4000 153.2000 ;
	    RECT 74.2000 152.8000 75.4000 153.1000 ;
	    RECT 77.4000 152.8000 77.8000 153.2000 ;
	    RECT 70.2000 152.1000 70.6000 152.2000 ;
	    RECT 71.0000 152.1000 71.4000 152.2000 ;
	    RECT 70.2000 151.8000 71.4000 152.1000 ;
	    RECT 72.6000 151.8000 73.0000 152.2000 ;
	    RECT 72.6000 149.2000 72.9000 151.8000 ;
	    RECT 74.2000 149.2000 74.5000 152.8000 ;
	    RECT 67.8000 148.8000 68.2000 149.2000 ;
	    RECT 67.0000 147.8000 67.4000 148.2000 ;
	    RECT 67.8000 146.2000 68.1000 148.8000 ;
	    RECT 67.8000 145.8000 68.2000 146.2000 ;
	    RECT 69.4000 146.1000 69.8000 146.2000 ;
	    RECT 70.2000 146.1000 70.6000 146.2000 ;
	    RECT 69.4000 145.8000 70.6000 146.1000 ;
	    RECT 71.0000 143.1000 71.4000 148.9000 ;
	    RECT 72.6000 148.8000 73.0000 149.2000 ;
	    RECT 74.2000 148.8000 74.6000 149.2000 ;
	    RECT 72.6000 145.2000 72.9000 148.8000 ;
	    RECT 72.6000 144.8000 73.0000 145.2000 ;
	    RECT 73.4000 144.1000 73.8000 144.2000 ;
	    RECT 74.2000 144.1000 74.6000 144.2000 ;
	    RECT 73.4000 143.8000 74.6000 144.1000 ;
	    RECT 76.6000 143.1000 77.0000 148.9000 ;
	    RECT 77.4000 146.8000 77.8000 147.2000 ;
	    RECT 77.4000 146.2000 77.7000 146.8000 ;
	    RECT 77.4000 145.8000 77.8000 146.2000 ;
	    RECT 64.6000 132.1000 65.0000 137.9000 ;
	    RECT 66.2000 135.1000 66.6000 135.2000 ;
	    RECT 67.0000 135.1000 67.4000 135.2000 ;
	    RECT 66.2000 134.8000 67.4000 135.1000 ;
	    RECT 67.8000 134.8000 68.2000 135.2000 ;
	    RECT 67.8000 129.2000 68.1000 134.8000 ;
	    RECT 69.4000 132.1000 69.8000 137.9000 ;
	    RECT 76.6000 136.8000 77.0000 137.2000 ;
	    RECT 70.2000 133.8000 70.6000 134.2000 ;
	    RECT 67.8000 128.8000 68.2000 129.2000 ;
	    RECT 62.2000 127.8000 62.6000 128.2000 ;
	    RECT 63.0000 127.8000 63.4000 128.2000 ;
	    RECT 63.0000 127.2000 63.3000 127.8000 ;
	    RECT 61.4000 126.8000 61.8000 127.2000 ;
	    RECT 63.0000 126.8000 63.4000 127.2000 ;
	    RECT 64.6000 126.8000 65.0000 127.2000 ;
	    RECT 65.4000 126.8000 65.8000 127.2000 ;
	    RECT 66.2000 126.8000 66.6000 127.2000 ;
	    RECT 64.6000 126.2000 64.9000 126.8000 ;
	    RECT 64.6000 125.8000 65.0000 126.2000 ;
	    RECT 65.4000 123.2000 65.7000 126.8000 ;
	    RECT 66.2000 126.2000 66.5000 126.8000 ;
	    RECT 66.2000 125.8000 66.6000 126.2000 ;
	    RECT 70.2000 124.2000 70.5000 133.8000 ;
	    RECT 71.0000 133.1000 71.4000 135.9000 ;
	    RECT 72.6000 131.8000 73.0000 132.2000 ;
	    RECT 75.0000 131.8000 75.4000 132.2000 ;
	    RECT 72.6000 129.2000 72.9000 131.8000 ;
	    RECT 68.6000 124.1000 69.0000 124.2000 ;
	    RECT 69.4000 124.1000 69.8000 124.2000 ;
	    RECT 68.6000 123.8000 69.8000 124.1000 ;
	    RECT 70.2000 123.8000 70.6000 124.2000 ;
	    RECT 65.4000 122.8000 65.8000 123.2000 ;
	    RECT 60.6000 121.8000 61.0000 122.2000 ;
	    RECT 50.2000 116.8000 50.6000 117.2000 ;
	    RECT 49.4000 112.8000 49.8000 113.2000 ;
	    RECT 50.2000 113.1000 50.6000 115.9000 ;
	    RECT 51.8000 112.1000 52.2000 117.9000 ;
	    RECT 55.8000 116.8000 56.2000 117.2000 ;
	    RECT 55.8000 115.2000 56.1000 116.8000 ;
	    RECT 53.4000 115.1000 53.8000 115.2000 ;
	    RECT 54.2000 115.1000 54.6000 115.2000 ;
	    RECT 53.4000 114.8000 54.6000 115.1000 ;
	    RECT 55.8000 114.8000 56.2000 115.2000 ;
	    RECT 56.6000 112.1000 57.0000 117.9000 ;
	    RECT 59.8000 115.1000 60.2000 115.2000 ;
	    RECT 60.6000 115.1000 61.0000 115.2000 ;
	    RECT 59.8000 114.8000 61.0000 115.1000 ;
	    RECT 63.0000 113.8000 63.4000 114.2000 ;
	    RECT 63.0000 112.2000 63.3000 113.8000 ;
	    RECT 63.8000 112.8000 64.2000 113.2000 ;
	    RECT 64.6000 113.1000 65.0000 115.9000 ;
	    RECT 59.0000 112.1000 59.4000 112.2000 ;
	    RECT 59.8000 112.1000 60.2000 112.2000 ;
	    RECT 59.0000 111.8000 60.2000 112.1000 ;
	    RECT 63.0000 111.8000 63.4000 112.2000 ;
	    RECT 63.8000 111.2000 64.1000 112.8000 ;
	    RECT 66.2000 112.1000 66.6000 117.9000 ;
	    RECT 70.2000 117.2000 70.5000 123.8000 ;
	    RECT 71.0000 123.1000 71.4000 128.9000 ;
	    RECT 72.6000 128.8000 73.0000 129.2000 ;
	    RECT 75.0000 128.2000 75.3000 131.8000 ;
	    RECT 75.0000 127.8000 75.4000 128.2000 ;
	    RECT 75.0000 126.8000 75.4000 127.2000 ;
	    RECT 75.0000 126.3000 75.3000 126.8000 ;
	    RECT 75.0000 125.9000 75.4000 126.3000 ;
	    RECT 75.8000 123.1000 76.2000 128.9000 ;
	    RECT 76.6000 127.2000 76.9000 136.8000 ;
	    RECT 77.4000 132.1000 77.8000 137.9000 ;
	    RECT 78.2000 128.2000 78.5000 153.8000 ;
	    RECT 79.8000 151.8000 80.2000 152.2000 ;
	    RECT 79.8000 146.2000 80.1000 151.8000 ;
	    RECT 79.8000 145.8000 80.2000 146.2000 ;
	    RECT 81.4000 143.1000 81.8000 148.9000 ;
	    RECT 82.2000 147.8000 82.6000 148.2000 ;
	    RECT 82.2000 147.2000 82.5000 147.8000 ;
	    RECT 82.2000 146.8000 82.6000 147.2000 ;
	    RECT 83.0000 145.1000 83.4000 147.9000 ;
	    RECT 83.8000 146.2000 84.1000 154.8000 ;
	    RECT 84.6000 149.2000 84.9000 155.8000 ;
	    RECT 91.0000 154.8000 91.4000 155.2000 ;
	    RECT 91.0000 154.2000 91.3000 154.8000 ;
	    RECT 86.2000 154.1000 86.6000 154.2000 ;
	    RECT 87.0000 154.1000 87.4000 154.2000 ;
	    RECT 86.2000 153.8000 87.4000 154.1000 ;
	    RECT 90.2000 153.8000 90.6000 154.2000 ;
	    RECT 91.0000 153.8000 91.4000 154.2000 ;
	    RECT 84.6000 148.8000 85.0000 149.2000 ;
	    RECT 85.4000 148.8000 85.8000 149.2000 ;
	    RECT 85.4000 147.2000 85.7000 148.8000 ;
	    RECT 85.4000 146.8000 85.8000 147.2000 ;
	    RECT 83.8000 145.8000 84.2000 146.2000 ;
	    RECT 85.4000 145.2000 85.7000 146.8000 ;
	    RECT 83.8000 144.8000 84.2000 145.2000 ;
	    RECT 85.4000 144.8000 85.8000 145.2000 ;
	    RECT 86.2000 145.1000 86.6000 147.9000 ;
	    RECT 87.0000 147.8000 87.4000 148.2000 ;
	    RECT 87.0000 147.2000 87.3000 147.8000 ;
	    RECT 87.0000 146.8000 87.4000 147.2000 ;
	    RECT 87.0000 145.8000 87.4000 146.2000 ;
	    RECT 83.8000 144.2000 84.1000 144.8000 ;
	    RECT 83.8000 143.8000 84.2000 144.2000 ;
	    RECT 83.8000 138.2000 84.1000 143.8000 ;
	    RECT 87.0000 142.2000 87.3000 145.8000 ;
	    RECT 87.8000 143.1000 88.2000 148.9000 ;
	    RECT 88.6000 146.1000 89.0000 146.2000 ;
	    RECT 89.4000 146.1000 89.8000 146.2000 ;
	    RECT 88.6000 145.8000 89.8000 146.1000 ;
	    RECT 90.2000 144.2000 90.5000 153.8000 ;
	    RECT 91.8000 146.2000 92.1000 165.8000 ;
	    RECT 92.6000 163.1000 93.0000 168.9000 ;
	    RECT 95.8000 168.2000 96.1000 174.8000 ;
	    RECT 98.2000 173.1000 98.6000 175.9000 ;
	    RECT 99.0000 173.8000 99.4000 174.2000 ;
	    RECT 99.0000 173.2000 99.3000 173.8000 ;
	    RECT 99.0000 172.8000 99.4000 173.2000 ;
	    RECT 99.8000 172.1000 100.2000 177.9000 ;
	    RECT 101.4000 174.8000 101.8000 175.2000 ;
	    RECT 101.4000 174.2000 101.7000 174.8000 ;
	    RECT 101.4000 173.8000 101.8000 174.2000 ;
	    RECT 103.8000 173.8000 104.2000 174.2000 ;
	    RECT 95.8000 167.8000 96.2000 168.2000 ;
	    RECT 103.8000 167.2000 104.1000 173.8000 ;
	    RECT 104.6000 172.1000 105.0000 177.9000 ;
	    RECT 114.2000 176.8000 114.6000 177.2000 ;
	    RECT 114.2000 175.2000 114.5000 176.8000 ;
	    RECT 106.2000 174.8000 106.6000 175.2000 ;
	    RECT 107.0000 175.1000 107.4000 175.2000 ;
	    RECT 107.8000 175.1000 108.2000 175.2000 ;
	    RECT 107.0000 174.8000 108.2000 175.1000 ;
	    RECT 111.8000 174.8000 112.2000 175.2000 ;
	    RECT 114.2000 174.8000 114.6000 175.2000 ;
	    RECT 106.2000 169.2000 106.5000 174.8000 ;
	    RECT 111.8000 172.2000 112.1000 174.8000 ;
	    RECT 107.0000 172.1000 107.4000 172.2000 ;
	    RECT 107.8000 172.1000 108.2000 172.2000 ;
	    RECT 107.0000 171.8000 108.2000 172.1000 ;
	    RECT 111.8000 171.8000 112.2000 172.2000 ;
	    RECT 116.6000 172.1000 117.0000 177.9000 ;
	    RECT 120.6000 174.7000 121.0000 175.1000 ;
	    RECT 120.6000 174.2000 120.9000 174.7000 ;
	    RECT 119.8000 173.8000 120.2000 174.2000 ;
	    RECT 120.6000 173.8000 121.0000 174.2000 ;
	    RECT 111.8000 171.2000 112.1000 171.8000 ;
	    RECT 111.8000 170.8000 112.2000 171.2000 ;
	    RECT 116.6000 170.8000 117.0000 171.2000 ;
	    RECT 106.2000 168.8000 106.6000 169.2000 ;
	    RECT 115.0000 169.1000 115.4000 169.2000 ;
	    RECT 115.8000 169.1000 116.2000 169.2000 ;
	    RECT 106.2000 168.2000 106.5000 168.8000 ;
	    RECT 106.2000 167.8000 106.6000 168.2000 ;
	    RECT 97.4000 166.8000 97.8000 167.2000 ;
	    RECT 100.6000 166.8000 101.0000 167.2000 ;
	    RECT 101.4000 166.8000 101.8000 167.2000 ;
	    RECT 102.2000 166.8000 102.6000 167.2000 ;
	    RECT 103.8000 166.8000 104.2000 167.2000 ;
	    RECT 97.4000 166.2000 97.7000 166.8000 ;
	    RECT 97.4000 165.8000 97.8000 166.2000 ;
	    RECT 98.2000 166.1000 98.6000 166.2000 ;
	    RECT 99.0000 166.1000 99.4000 166.2000 ;
	    RECT 98.2000 165.8000 99.4000 166.1000 ;
	    RECT 99.8000 165.8000 100.2000 166.2000 ;
	    RECT 99.0000 163.2000 99.3000 165.8000 ;
	    RECT 99.8000 165.2000 100.1000 165.8000 ;
	    RECT 99.8000 164.8000 100.2000 165.2000 ;
	    RECT 99.0000 162.8000 99.4000 163.2000 ;
	    RECT 99.8000 156.8000 100.2000 157.2000 ;
	    RECT 99.8000 156.2000 100.1000 156.8000 ;
	    RECT 95.0000 155.8000 95.4000 156.2000 ;
	    RECT 99.8000 155.8000 100.2000 156.2000 ;
	    RECT 93.4000 153.8000 93.8000 154.2000 ;
	    RECT 93.4000 149.2000 93.7000 153.8000 ;
	    RECT 95.0000 153.2000 95.3000 155.8000 ;
	    RECT 99.8000 153.8000 100.2000 154.2000 ;
	    RECT 99.8000 153.2000 100.1000 153.8000 ;
	    RECT 100.6000 153.2000 100.9000 166.8000 ;
	    RECT 101.4000 166.2000 101.7000 166.8000 ;
	    RECT 101.4000 165.8000 101.8000 166.2000 ;
	    RECT 102.2000 164.2000 102.5000 166.8000 ;
	    RECT 107.0000 165.1000 107.4000 167.9000 ;
	    RECT 107.8000 167.8000 108.2000 168.2000 ;
	    RECT 107.8000 167.2000 108.1000 167.8000 ;
	    RECT 107.8000 166.8000 108.2000 167.2000 ;
	    RECT 102.2000 163.8000 102.6000 164.2000 ;
	    RECT 108.6000 163.1000 109.0000 168.9000 ;
	    RECT 109.4000 166.2000 109.8000 166.3000 ;
	    RECT 110.2000 166.2000 110.6000 166.3000 ;
	    RECT 109.4000 165.9000 110.6000 166.2000 ;
	    RECT 113.4000 163.1000 113.8000 168.9000 ;
	    RECT 115.0000 168.8000 116.2000 169.1000 ;
	    RECT 116.6000 168.2000 116.9000 170.8000 ;
	    RECT 119.8000 169.2000 120.1000 173.8000 ;
	    RECT 120.6000 172.8000 121.0000 173.2000 ;
	    RECT 120.6000 172.2000 120.9000 172.8000 ;
	    RECT 120.6000 171.8000 121.0000 172.2000 ;
	    RECT 121.4000 172.1000 121.8000 177.9000 ;
	    RECT 123.0000 173.1000 123.4000 175.9000 ;
	    RECT 125.4000 174.8000 125.8000 175.2000 ;
	    RECT 126.2000 174.8000 126.6000 175.2000 ;
	    RECT 129.4000 174.8000 129.8000 175.2000 ;
	    RECT 121.4000 169.8000 121.8000 170.2000 ;
	    RECT 121.4000 169.2000 121.7000 169.8000 ;
	    RECT 125.4000 169.2000 125.7000 174.8000 ;
	    RECT 119.8000 168.8000 120.2000 169.2000 ;
	    RECT 121.4000 168.8000 121.8000 169.2000 ;
	    RECT 116.6000 167.8000 117.0000 168.2000 ;
	    RECT 120.6000 167.8000 121.0000 168.2000 ;
	    RECT 119.0000 166.8000 119.4000 167.2000 ;
	    RECT 119.0000 164.2000 119.3000 166.8000 ;
	    RECT 119.0000 163.8000 119.4000 164.2000 ;
	    RECT 120.6000 162.2000 120.9000 167.8000 ;
	    RECT 123.8000 163.1000 124.2000 168.9000 ;
	    RECT 125.4000 168.8000 125.8000 169.2000 ;
	    RECT 126.2000 163.2000 126.5000 174.8000 ;
	    RECT 127.0000 174.1000 127.4000 174.2000 ;
	    RECT 127.8000 174.1000 128.2000 174.2000 ;
	    RECT 127.0000 173.8000 128.2000 174.1000 ;
	    RECT 129.4000 173.2000 129.7000 174.8000 ;
	    RECT 129.4000 172.8000 129.8000 173.2000 ;
	    RECT 132.6000 173.1000 133.0000 175.9000 ;
	    RECT 133.4000 173.8000 133.8000 174.2000 ;
	    RECT 133.4000 172.2000 133.7000 173.8000 ;
	    RECT 129.4000 171.8000 129.8000 172.2000 ;
	    RECT 133.4000 171.8000 133.8000 172.2000 ;
	    RECT 134.2000 172.1000 134.6000 177.9000 ;
	    RECT 135.8000 174.8000 136.2000 175.2000 ;
	    RECT 127.8000 166.8000 128.2000 167.2000 ;
	    RECT 127.8000 166.3000 128.1000 166.8000 ;
	    RECT 127.8000 165.9000 128.2000 166.3000 ;
	    RECT 126.2000 162.8000 126.6000 163.2000 ;
	    RECT 128.6000 163.1000 129.0000 168.9000 ;
	    RECT 129.4000 167.2000 129.7000 171.8000 ;
	    RECT 135.8000 169.2000 136.1000 174.8000 ;
	    RECT 139.0000 172.1000 139.4000 177.9000 ;
	    RECT 154.2000 176.8000 154.6000 177.2000 ;
	    RECT 154.2000 175.2000 154.5000 176.8000 ;
	    RECT 142.2000 174.8000 142.6000 175.2000 ;
	    RECT 144.6000 174.8000 145.0000 175.2000 ;
	    RECT 147.0000 174.8000 147.4000 175.2000 ;
	    RECT 149.4000 174.8000 149.8000 175.2000 ;
	    RECT 153.4000 174.8000 153.8000 175.2000 ;
	    RECT 154.2000 174.8000 154.6000 175.2000 ;
	    RECT 139.8000 171.8000 140.2000 172.2000 ;
	    RECT 140.6000 172.1000 141.0000 172.2000 ;
	    RECT 141.4000 172.1000 141.8000 172.2000 ;
	    RECT 140.6000 171.8000 141.8000 172.1000 ;
	    RECT 131.0000 168.8000 131.4000 169.2000 ;
	    RECT 135.8000 168.8000 136.2000 169.2000 ;
	    RECT 131.0000 168.2000 131.3000 168.8000 ;
	    RECT 139.8000 168.2000 140.1000 171.8000 ;
	    RECT 129.4000 166.8000 129.8000 167.2000 ;
	    RECT 120.6000 161.8000 121.0000 162.2000 ;
	    RECT 101.4000 156.8000 101.8000 157.2000 ;
	    RECT 101.4000 156.2000 101.7000 156.8000 ;
	    RECT 101.4000 155.8000 101.8000 156.2000 ;
	    RECT 103.0000 156.1000 103.4000 156.2000 ;
	    RECT 103.8000 156.1000 104.2000 156.2000 ;
	    RECT 103.0000 155.8000 104.2000 156.1000 ;
	    RECT 104.6000 155.8000 105.0000 156.2000 ;
	    RECT 107.8000 155.8000 108.2000 156.2000 ;
	    RECT 104.6000 153.2000 104.9000 155.8000 ;
	    RECT 107.8000 155.2000 108.1000 155.8000 ;
	    RECT 107.8000 154.8000 108.2000 155.2000 ;
	    RECT 107.8000 153.2000 108.1000 154.8000 ;
	    RECT 95.0000 152.8000 95.4000 153.2000 ;
	    RECT 95.8000 152.8000 96.2000 153.2000 ;
	    RECT 98.2000 152.8000 98.6000 153.2000 ;
	    RECT 99.8000 152.8000 100.2000 153.2000 ;
	    RECT 100.6000 152.8000 101.0000 153.2000 ;
	    RECT 102.2000 152.8000 102.6000 153.2000 ;
	    RECT 103.0000 152.8000 103.4000 153.2000 ;
	    RECT 104.6000 152.8000 105.0000 153.2000 ;
	    RECT 107.8000 152.8000 108.2000 153.2000 ;
	    RECT 111.8000 152.8000 112.2000 153.2000 ;
	    RECT 91.8000 145.8000 92.2000 146.2000 ;
	    RECT 88.6000 143.8000 89.0000 144.2000 ;
	    RECT 90.2000 143.8000 90.6000 144.2000 ;
	    RECT 87.0000 141.8000 87.4000 142.2000 ;
	    RECT 85.4000 139.1000 85.8000 139.2000 ;
	    RECT 86.2000 139.1000 86.6000 139.2000 ;
	    RECT 85.4000 138.8000 86.6000 139.1000 ;
	    RECT 79.0000 134.8000 79.4000 135.2000 ;
	    RECT 79.0000 134.2000 79.3000 134.8000 ;
	    RECT 79.0000 133.8000 79.4000 134.2000 ;
	    RECT 82.2000 132.1000 82.6000 137.9000 ;
	    RECT 83.8000 137.8000 84.2000 138.2000 ;
	    RECT 83.0000 133.8000 83.4000 134.2000 ;
	    RECT 76.6000 126.8000 77.0000 127.2000 ;
	    RECT 76.6000 125.8000 77.0000 126.2000 ;
	    RECT 76.6000 119.2000 76.9000 125.8000 ;
	    RECT 77.4000 125.1000 77.8000 127.9000 ;
	    RECT 78.2000 127.8000 78.6000 128.2000 ;
	    RECT 79.0000 127.8000 79.4000 128.2000 ;
	    RECT 76.6000 118.8000 77.0000 119.2000 ;
	    RECT 70.2000 116.8000 70.6000 117.2000 ;
	    RECT 70.2000 115.2000 70.5000 116.8000 ;
	    RECT 67.8000 114.8000 68.2000 115.2000 ;
	    RECT 70.2000 114.8000 70.6000 115.2000 ;
	    RECT 63.8000 110.8000 64.2000 111.2000 ;
	    RECT 63.8000 109.8000 64.2000 110.2000 ;
	    RECT 66.2000 109.8000 66.6000 110.2000 ;
	    RECT 52.6000 108.8000 53.0000 109.2000 ;
	    RECT 55.8000 108.8000 56.2000 109.2000 ;
	    RECT 59.8000 108.8000 60.2000 109.2000 ;
	    RECT 52.6000 108.2000 52.9000 108.8000 ;
	    RECT 37.4000 107.8000 37.8000 108.2000 ;
	    RECT 42.2000 107.8000 42.6000 108.2000 ;
	    RECT 44.6000 108.1000 45.0000 108.2000 ;
	    RECT 45.4000 108.1000 45.8000 108.2000 ;
	    RECT 44.6000 107.8000 45.8000 108.1000 ;
	    RECT 48.6000 107.8000 49.0000 108.2000 ;
	    RECT 51.0000 108.1000 51.4000 108.2000 ;
	    RECT 51.8000 108.1000 52.2000 108.2000 ;
	    RECT 51.0000 107.8000 52.2000 108.1000 ;
	    RECT 52.6000 107.8000 53.0000 108.2000 ;
	    RECT 42.2000 107.2000 42.5000 107.8000 ;
	    RECT 42.2000 106.8000 42.6000 107.2000 ;
	    RECT 45.4000 106.8000 45.8000 107.2000 ;
	    RECT 35.0000 105.8000 35.4000 106.2000 ;
	    RECT 36.6000 105.8000 37.0000 106.2000 ;
	    RECT 40.6000 106.1000 41.0000 106.2000 ;
	    RECT 41.4000 106.1000 41.8000 106.2000 ;
	    RECT 40.6000 105.8000 41.8000 106.1000 ;
	    RECT 33.4000 103.8000 33.8000 104.2000 ;
	    RECT 35.8000 103.8000 36.2000 104.2000 ;
	    RECT 31.8000 102.8000 32.2000 103.2000 ;
	    RECT 23.0000 95.8000 23.4000 96.2000 ;
	    RECT 25.4000 95.8000 25.8000 96.2000 ;
	    RECT 26.2000 95.8000 26.6000 96.2000 ;
	    RECT 28.6000 95.8000 29.0000 96.2000 ;
	    RECT 23.8000 95.1000 24.2000 95.2000 ;
	    RECT 24.6000 95.1000 25.0000 95.2000 ;
	    RECT 23.8000 94.8000 25.0000 95.1000 ;
	    RECT 26.2000 94.2000 26.5000 95.8000 ;
	    RECT 28.6000 95.2000 28.9000 95.8000 ;
	    RECT 28.6000 94.8000 29.0000 95.2000 ;
	    RECT 35.8000 94.2000 36.1000 103.8000 ;
	    RECT 45.4000 99.2000 45.7000 106.8000 ;
	    RECT 48.6000 106.2000 48.9000 107.8000 ;
	    RECT 55.8000 107.2000 56.1000 108.8000 ;
	    RECT 58.2000 107.8000 58.6000 108.2000 ;
	    RECT 58.2000 107.2000 58.5000 107.8000 ;
	    RECT 59.8000 107.2000 60.1000 108.8000 ;
	    RECT 63.8000 108.2000 64.1000 109.8000 ;
	    RECT 65.4000 108.8000 65.8000 109.2000 ;
	    RECT 63.8000 107.8000 64.2000 108.2000 ;
	    RECT 54.2000 107.1000 54.6000 107.2000 ;
	    RECT 55.0000 107.1000 55.4000 107.2000 ;
	    RECT 54.2000 106.8000 55.4000 107.1000 ;
	    RECT 55.8000 106.8000 56.2000 107.2000 ;
	    RECT 58.2000 106.8000 58.6000 107.2000 ;
	    RECT 59.8000 106.8000 60.2000 107.2000 ;
	    RECT 47.8000 105.8000 48.2000 106.2000 ;
	    RECT 48.6000 105.8000 49.0000 106.2000 ;
	    RECT 55.0000 105.8000 55.4000 106.2000 ;
	    RECT 61.4000 105.8000 61.8000 106.2000 ;
	    RECT 47.0000 101.8000 47.4000 102.2000 ;
	    RECT 45.4000 98.8000 45.8000 99.2000 ;
	    RECT 36.6000 96.8000 37.0000 97.2000 ;
	    RECT 40.6000 96.8000 41.0000 97.2000 ;
	    RECT 36.6000 96.2000 36.9000 96.8000 ;
	    RECT 36.6000 95.8000 37.0000 96.2000 ;
	    RECT 38.2000 95.9000 38.6000 96.3000 ;
	    RECT 38.2000 94.2000 38.5000 95.9000 ;
	    RECT 40.6000 95.2000 40.9000 96.8000 ;
	    RECT 41.5000 95.9000 41.9000 96.3000 ;
	    RECT 47.0000 96.2000 47.3000 101.8000 ;
	    RECT 40.6000 94.8000 41.0000 95.2000 ;
	    RECT 40.2000 94.2000 40.6000 94.3000 ;
	    RECT 7.8000 92.8000 8.2000 93.2000 ;
	    RECT 13.4000 92.8000 13.8000 93.2000 ;
	    RECT 18.2000 93.1000 18.6000 93.5000 ;
	    RECT 18.9000 93.2000 21.7000 93.5000 ;
	    RECT 21.3000 93.1000 21.7000 93.2000 ;
	    RECT 23.0000 93.8000 23.4000 94.2000 ;
	    RECT 24.6000 93.8000 25.0000 94.2000 ;
	    RECT 26.2000 93.8000 26.6000 94.2000 ;
	    RECT 29.4000 93.8000 29.8000 94.2000 ;
	    RECT 35.8000 93.8000 36.2000 94.2000 ;
	    RECT 36.6000 94.1000 37.0000 94.2000 ;
	    RECT 37.4000 94.1000 37.8000 94.2000 ;
	    RECT 36.6000 93.8000 37.8000 94.1000 ;
	    RECT 38.2000 93.9000 40.6000 94.2000 ;
	    RECT 23.0000 93.2000 23.3000 93.8000 ;
	    RECT 23.0000 92.8000 23.4000 93.2000 ;
	    RECT 4.6000 91.8000 5.0000 92.2000 ;
	    RECT 4.6000 85.2000 4.9000 91.8000 ;
	    RECT 7.8000 89.2000 8.1000 92.8000 ;
	    RECT 16.6000 91.8000 17.0000 92.2000 ;
	    RECT 20.6000 91.8000 21.0000 92.2000 ;
	    RECT 7.8000 88.8000 8.2000 89.2000 ;
	    RECT 13.4000 89.1000 13.8000 89.2000 ;
	    RECT 14.2000 89.1000 14.6000 89.2000 ;
	    RECT 13.4000 88.8000 14.6000 89.1000 ;
	    RECT 11.9000 87.8000 12.3000 87.9000 ;
	    RECT 11.9000 87.5000 14.7000 87.8000 ;
	    RECT 15.0000 87.5000 15.4000 87.9000 ;
	    RECT 0.6000 85.1000 1.0000 85.2000 ;
	    RECT 1.4000 85.1000 1.8000 85.2000 ;
	    RECT 0.6000 84.8000 1.8000 85.1000 ;
	    RECT 2.2000 84.8000 2.6000 85.2000 ;
	    RECT 4.6000 84.8000 5.0000 85.2000 ;
	    RECT 11.9000 85.1000 12.2000 87.5000 ;
	    RECT 12.6000 87.4000 13.0000 87.5000 ;
	    RECT 14.3000 87.4000 14.7000 87.5000 ;
	    RECT 15.1000 87.1000 15.4000 87.5000 ;
	    RECT 12.6000 86.8000 15.4000 87.1000 ;
	    RECT 12.6000 86.1000 12.9000 86.8000 ;
	    RECT 12.5000 85.7000 12.9000 86.1000 ;
	    RECT 15.1000 85.1000 15.4000 86.8000 ;
	    RECT 11.9000 84.7000 12.3000 85.1000 ;
	    RECT 15.0000 84.7000 15.4000 85.1000 ;
	    RECT 16.6000 85.2000 16.9000 91.8000 ;
	    RECT 19.0000 88.8000 19.4000 89.2000 ;
	    RECT 19.0000 88.2000 19.3000 88.8000 ;
	    RECT 19.0000 87.8000 19.4000 88.2000 ;
	    RECT 20.6000 86.2000 20.9000 91.8000 ;
	    RECT 24.6000 89.2000 24.9000 93.8000 ;
	    RECT 27.0000 91.8000 27.4000 92.2000 ;
	    RECT 27.0000 89.2000 27.3000 91.8000 ;
	    RECT 29.4000 89.2000 29.7000 93.8000 ;
	    RECT 35.8000 93.2000 36.1000 93.8000 ;
	    RECT 38.2000 93.5000 38.5000 93.9000 ;
	    RECT 38.9000 93.5000 39.3000 93.6000 ;
	    RECT 40.6000 93.5000 41.0000 93.6000 ;
	    RECT 41.6000 93.5000 41.9000 95.9000 ;
	    RECT 43.0000 95.8000 43.4000 96.2000 ;
	    RECT 47.0000 95.8000 47.4000 96.2000 ;
	    RECT 43.0000 95.2000 43.3000 95.8000 ;
	    RECT 43.0000 94.8000 43.4000 95.2000 ;
	    RECT 35.8000 92.8000 36.2000 93.2000 ;
	    RECT 38.2000 93.1000 38.6000 93.5000 ;
	    RECT 38.9000 93.2000 41.0000 93.5000 ;
	    RECT 41.5000 93.1000 41.9000 93.5000 ;
	    RECT 42.2000 93.8000 42.6000 94.2000 ;
	    RECT 47.0000 93.8000 47.4000 94.2000 ;
	    RECT 42.2000 92.2000 42.5000 93.8000 ;
	    RECT 47.0000 93.2000 47.3000 93.8000 ;
	    RECT 47.8000 93.2000 48.1000 105.8000 ;
	    RECT 50.2000 105.1000 50.6000 105.2000 ;
	    RECT 51.0000 105.1000 51.4000 105.2000 ;
	    RECT 50.2000 104.8000 51.4000 105.1000 ;
	    RECT 53.4000 104.8000 53.8000 105.2000 ;
	    RECT 52.6000 95.8000 53.0000 96.2000 ;
	    RECT 48.6000 94.8000 49.0000 95.2000 ;
	    RECT 49.4000 94.8000 49.8000 95.2000 ;
	    RECT 50.2000 95.1000 50.6000 95.2000 ;
	    RECT 51.0000 95.1000 51.4000 95.2000 ;
	    RECT 50.2000 94.8000 51.4000 95.1000 ;
	    RECT 48.6000 94.2000 48.9000 94.8000 ;
	    RECT 48.6000 93.8000 49.0000 94.2000 ;
	    RECT 43.0000 93.1000 43.4000 93.2000 ;
	    RECT 43.8000 93.1000 44.2000 93.2000 ;
	    RECT 43.0000 92.8000 44.2000 93.1000 ;
	    RECT 44.6000 92.8000 45.0000 93.2000 ;
	    RECT 46.2000 92.8000 46.6000 93.2000 ;
	    RECT 47.0000 92.8000 47.4000 93.2000 ;
	    RECT 47.8000 92.8000 48.2000 93.2000 ;
	    RECT 49.4000 93.1000 49.7000 94.8000 ;
	    RECT 52.6000 94.2000 52.9000 95.8000 ;
	    RECT 53.4000 94.2000 53.7000 104.8000 ;
	    RECT 55.0000 104.2000 55.3000 105.8000 ;
	    RECT 61.4000 104.2000 61.7000 105.8000 ;
	    RECT 65.4000 104.2000 65.7000 108.8000 ;
	    RECT 66.2000 106.2000 66.5000 109.8000 ;
	    RECT 67.8000 108.2000 68.1000 114.8000 ;
	    RECT 71.0000 112.1000 71.4000 117.9000 ;
	    RECT 73.4000 116.8000 73.8000 117.2000 ;
	    RECT 75.0000 117.1000 75.4000 117.2000 ;
	    RECT 75.8000 117.1000 76.2000 117.2000 ;
	    RECT 75.0000 116.8000 76.2000 117.1000 ;
	    RECT 67.8000 107.8000 68.2000 108.2000 ;
	    RECT 66.2000 105.8000 66.6000 106.2000 ;
	    RECT 55.0000 103.8000 55.4000 104.2000 ;
	    RECT 61.4000 103.8000 61.8000 104.2000 ;
	    RECT 65.4000 103.8000 65.8000 104.2000 ;
	    RECT 67.8000 104.1000 68.2000 104.2000 ;
	    RECT 68.6000 104.1000 69.0000 104.2000 ;
	    RECT 67.8000 103.8000 69.0000 104.1000 ;
	    RECT 70.2000 103.1000 70.6000 108.9000 ;
	    RECT 71.0000 105.8000 71.4000 106.2000 ;
	    RECT 57.4000 102.1000 57.8000 102.2000 ;
	    RECT 58.2000 102.1000 58.6000 102.2000 ;
	    RECT 57.4000 101.8000 58.6000 102.1000 ;
	    RECT 63.8000 101.8000 64.2000 102.2000 ;
	    RECT 66.2000 101.8000 66.6000 102.2000 ;
	    RECT 63.8000 99.2000 64.1000 101.8000 ;
	    RECT 63.8000 98.8000 64.2000 99.2000 ;
	    RECT 66.2000 98.2000 66.5000 101.8000 ;
	    RECT 61.4000 95.8000 61.8000 96.2000 ;
	    RECT 61.4000 95.2000 61.7000 95.8000 ;
	    RECT 54.2000 94.8000 54.6000 95.2000 ;
	    RECT 61.4000 94.8000 61.8000 95.2000 ;
	    RECT 48.6000 92.8000 49.7000 93.1000 ;
	    RECT 50.2000 93.8000 50.6000 94.2000 ;
	    RECT 52.6000 93.8000 53.0000 94.2000 ;
	    RECT 53.4000 93.8000 53.8000 94.2000 ;
	    RECT 50.2000 93.2000 50.5000 93.8000 ;
	    RECT 50.2000 92.8000 50.6000 93.2000 ;
	    RECT 44.6000 92.2000 44.9000 92.8000 ;
	    RECT 46.2000 92.2000 46.5000 92.8000 ;
	    RECT 30.2000 91.8000 30.6000 92.2000 ;
	    RECT 38.2000 91.8000 38.6000 92.2000 ;
	    RECT 42.2000 91.8000 42.6000 92.2000 ;
	    RECT 44.6000 91.8000 45.0000 92.2000 ;
	    RECT 46.2000 91.8000 46.6000 92.2000 ;
	    RECT 47.8000 91.8000 48.2000 92.2000 ;
	    RECT 30.2000 90.2000 30.5000 91.8000 ;
	    RECT 30.2000 89.8000 30.6000 90.2000 ;
	    RECT 38.2000 89.2000 38.5000 91.8000 ;
	    RECT 47.8000 89.2000 48.1000 91.8000 ;
	    RECT 48.6000 89.2000 48.9000 92.8000 ;
	    RECT 54.2000 92.2000 54.5000 94.8000 ;
	    RECT 60.6000 93.8000 61.0000 94.2000 ;
	    RECT 55.0000 93.1000 55.4000 93.2000 ;
	    RECT 55.8000 93.1000 56.2000 93.2000 ;
	    RECT 55.0000 92.8000 56.2000 93.1000 ;
	    RECT 59.0000 93.1000 59.4000 93.2000 ;
	    RECT 59.8000 93.1000 60.2000 93.2000 ;
	    RECT 59.0000 92.8000 60.2000 93.1000 ;
	    RECT 54.2000 91.8000 54.6000 92.2000 ;
	    RECT 57.4000 91.8000 57.8000 92.2000 ;
	    RECT 59.8000 91.8000 60.2000 92.2000 ;
	    RECT 24.6000 88.8000 25.0000 89.2000 ;
	    RECT 27.0000 88.8000 27.4000 89.2000 ;
	    RECT 29.4000 88.8000 29.8000 89.2000 ;
	    RECT 38.2000 88.8000 38.6000 89.2000 ;
	    RECT 22.1000 87.5000 22.5000 87.9000 ;
	    RECT 25.4000 87.5000 25.8000 87.9000 ;
	    RECT 20.6000 85.8000 21.0000 86.2000 ;
	    RECT 16.6000 84.8000 17.0000 85.2000 ;
	    RECT 22.1000 85.1000 22.4000 87.5000 ;
	    RECT 25.5000 87.1000 25.8000 87.5000 ;
	    RECT 23.4000 86.8000 25.8000 87.1000 ;
	    RECT 23.4000 86.7000 23.8000 86.8000 ;
	    RECT 25.5000 85.1000 25.8000 86.8000 ;
	    RECT 22.1000 84.7000 22.5000 85.1000 ;
	    RECT 25.4000 84.7000 25.8000 85.1000 ;
	    RECT 27.8000 87.5000 28.2000 87.9000 ;
	    RECT 31.1000 87.5000 31.5000 87.9000 ;
	    RECT 27.8000 87.1000 28.1000 87.5000 ;
	    RECT 27.8000 86.8000 30.2000 87.1000 ;
	    RECT 27.8000 85.1000 28.1000 86.8000 ;
	    RECT 29.8000 86.7000 30.2000 86.8000 ;
	    RECT 31.2000 85.1000 31.5000 87.5000 ;
	    RECT 27.8000 84.7000 28.2000 85.1000 ;
	    RECT 31.1000 84.7000 31.5000 85.1000 ;
	    RECT 33.5000 87.8000 33.9000 87.9000 ;
	    RECT 33.5000 87.5000 36.3000 87.8000 ;
	    RECT 36.6000 87.5000 37.0000 87.9000 ;
	    RECT 33.5000 85.1000 33.8000 87.5000 ;
	    RECT 34.2000 87.4000 34.6000 87.5000 ;
	    RECT 35.9000 87.4000 36.3000 87.5000 ;
	    RECT 36.7000 87.1000 37.0000 87.5000 ;
	    RECT 34.2000 86.8000 37.0000 87.1000 ;
	    RECT 34.2000 86.1000 34.5000 86.8000 ;
	    RECT 34.1000 85.7000 34.5000 86.1000 ;
	    RECT 36.7000 85.1000 37.0000 86.8000 ;
	    RECT 33.5000 84.7000 33.9000 85.1000 ;
	    RECT 36.6000 84.7000 37.0000 85.1000 ;
	    RECT 40.6000 83.1000 41.0000 88.9000 ;
	    RECT 44.6000 86.8000 45.0000 87.2000 ;
	    RECT 44.6000 86.3000 44.9000 86.8000 ;
	    RECT 44.6000 85.9000 45.0000 86.3000 ;
	    RECT 45.4000 83.1000 45.8000 88.9000 ;
	    RECT 47.8000 88.8000 48.2000 89.2000 ;
	    RECT 48.6000 88.8000 49.0000 89.2000 ;
	    RECT 53.4000 88.8000 53.8000 89.2000 ;
	    RECT 46.2000 86.8000 46.6000 87.2000 ;
	    RECT 17.4000 81.8000 17.8000 82.2000 ;
	    RECT 35.0000 81.8000 35.4000 82.2000 ;
	    RECT 17.4000 78.2000 17.7000 81.8000 ;
	    RECT 7.8000 78.1000 8.2000 78.2000 ;
	    RECT 8.6000 78.1000 9.0000 78.2000 ;
	    RECT 7.8000 77.8000 9.0000 78.1000 ;
	    RECT 10.2000 77.8000 10.6000 78.2000 ;
	    RECT 17.4000 77.8000 17.8000 78.2000 ;
	    RECT 10.2000 77.2000 10.5000 77.8000 ;
	    RECT 5.4000 76.8000 5.8000 77.2000 ;
	    RECT 10.2000 76.8000 10.6000 77.2000 ;
	    RECT 17.4000 76.8000 17.8000 77.2000 ;
	    RECT 27.0000 76.8000 27.4000 77.2000 ;
	    RECT 30.2000 76.8000 30.6000 77.2000 ;
	    RECT 31.0000 76.8000 31.4000 77.2000 ;
	    RECT 5.4000 75.2000 5.7000 76.8000 ;
	    RECT 17.4000 76.2000 17.7000 76.8000 ;
	    RECT 27.0000 76.2000 27.3000 76.8000 ;
	    RECT 30.2000 76.2000 30.5000 76.8000 ;
	    RECT 31.0000 76.2000 31.3000 76.8000 ;
	    RECT 16.6000 75.8000 17.0000 76.2000 ;
	    RECT 17.4000 75.8000 17.8000 76.2000 ;
	    RECT 20.6000 76.1000 21.0000 76.2000 ;
	    RECT 21.4000 76.1000 21.8000 76.2000 ;
	    RECT 20.6000 75.8000 21.8000 76.1000 ;
	    RECT 23.0000 76.1000 23.4000 76.2000 ;
	    RECT 23.8000 76.1000 24.2000 76.2000 ;
	    RECT 23.0000 75.8000 24.2000 76.1000 ;
	    RECT 25.4000 75.8000 25.8000 76.2000 ;
	    RECT 27.0000 75.8000 27.4000 76.2000 ;
	    RECT 30.2000 75.8000 30.6000 76.2000 ;
	    RECT 31.0000 75.8000 31.4000 76.2000 ;
	    RECT 16.6000 75.2000 16.9000 75.8000 ;
	    RECT 25.4000 75.2000 25.7000 75.8000 ;
	    RECT 35.0000 75.2000 35.3000 81.8000 ;
	    RECT 46.2000 79.2000 46.5000 86.8000 ;
	    RECT 47.0000 85.1000 47.4000 87.9000 ;
	    RECT 49.4000 87.8000 49.8000 88.2000 ;
	    RECT 51.8000 87.8000 52.2000 88.2000 ;
	    RECT 49.4000 87.2000 49.7000 87.8000 ;
	    RECT 49.4000 86.8000 49.8000 87.2000 ;
	    RECT 51.8000 86.2000 52.1000 87.8000 ;
	    RECT 47.8000 85.8000 48.2000 86.2000 ;
	    RECT 51.8000 85.8000 52.2000 86.2000 ;
	    RECT 47.8000 83.2000 48.1000 85.8000 ;
	    RECT 50.2000 84.1000 50.6000 84.2000 ;
	    RECT 51.0000 84.1000 51.4000 84.2000 ;
	    RECT 50.2000 83.8000 51.4000 84.1000 ;
	    RECT 47.8000 82.8000 48.2000 83.2000 ;
	    RECT 46.2000 78.8000 46.6000 79.2000 ;
	    RECT 44.6000 76.8000 45.0000 77.2000 ;
	    RECT 36.6000 75.9000 37.0000 76.3000 ;
	    RECT 39.7000 75.9000 40.1000 76.3000 ;
	    RECT 44.6000 76.2000 44.9000 76.8000 ;
	    RECT 2.2000 74.8000 2.6000 75.2000 ;
	    RECT 3.8000 75.1000 4.2000 75.2000 ;
	    RECT 4.6000 75.1000 5.0000 75.2000 ;
	    RECT 3.8000 74.8000 5.0000 75.1000 ;
	    RECT 5.4000 74.8000 5.8000 75.2000 ;
	    RECT 6.2000 74.8000 6.6000 75.2000 ;
	    RECT 10.2000 74.8000 10.6000 75.2000 ;
	    RECT 16.6000 74.8000 17.0000 75.2000 ;
	    RECT 25.4000 74.8000 25.8000 75.2000 ;
	    RECT 27.8000 75.1000 28.2000 75.2000 ;
	    RECT 28.6000 75.1000 29.0000 75.2000 ;
	    RECT 27.8000 74.8000 29.0000 75.1000 ;
	    RECT 35.0000 74.8000 35.4000 75.2000 ;
	    RECT 2.2000 74.2000 2.5000 74.8000 ;
	    RECT 6.2000 74.2000 6.5000 74.8000 ;
	    RECT 2.2000 73.8000 2.6000 74.2000 ;
	    RECT 6.2000 73.8000 6.6000 74.2000 ;
	    RECT 10.2000 69.2000 10.5000 74.8000 ;
	    RECT 36.6000 74.2000 36.9000 75.9000 ;
	    RECT 39.1000 74.9000 39.5000 75.3000 ;
	    RECT 39.1000 74.2000 39.4000 74.9000 ;
	    RECT 17.4000 74.1000 17.8000 74.2000 ;
	    RECT 18.2000 74.1000 18.6000 74.2000 ;
	    RECT 17.4000 73.8000 18.6000 74.1000 ;
	    RECT 22.2000 73.8000 22.6000 74.2000 ;
	    RECT 24.6000 73.8000 25.0000 74.2000 ;
	    RECT 27.0000 74.1000 27.4000 74.2000 ;
	    RECT 27.8000 74.1000 28.2000 74.2000 ;
	    RECT 26.2000 73.8000 28.2000 74.1000 ;
	    RECT 29.4000 73.8000 29.8000 74.2000 ;
	    RECT 36.6000 73.9000 39.4000 74.2000 ;
	    RECT 22.2000 73.2000 22.5000 73.8000 ;
	    RECT 24.6000 73.2000 24.9000 73.8000 ;
	    RECT 14.2000 73.1000 14.6000 73.2000 ;
	    RECT 15.0000 73.1000 15.4000 73.2000 ;
	    RECT 14.2000 72.8000 15.4000 73.1000 ;
	    RECT 22.2000 72.8000 22.6000 73.2000 ;
	    RECT 24.6000 72.8000 25.0000 73.2000 ;
	    RECT 14.2000 71.8000 14.6000 72.2000 ;
	    RECT 22.2000 72.1000 22.6000 72.2000 ;
	    RECT 23.0000 72.1000 23.4000 72.2000 ;
	    RECT 22.2000 71.8000 23.4000 72.1000 ;
	    RECT 23.8000 71.8000 24.2000 72.2000 ;
	    RECT 14.2000 69.2000 14.5000 71.8000 ;
	    RECT 17.4000 70.8000 17.8000 71.2000 ;
	    RECT 23.0000 70.8000 23.4000 71.2000 ;
	    RECT 17.4000 69.2000 17.7000 70.8000 ;
	    RECT 23.0000 69.2000 23.3000 70.8000 ;
	    RECT 10.2000 68.8000 10.6000 69.2000 ;
	    RECT 14.2000 68.8000 14.6000 69.2000 ;
	    RECT 17.4000 68.8000 17.8000 69.2000 ;
	    RECT 18.2000 68.8000 18.6000 69.2000 ;
	    RECT 23.0000 68.8000 23.4000 69.2000 ;
	    RECT 18.2000 68.2000 18.5000 68.8000 ;
	    RECT 23.8000 68.2000 24.1000 71.8000 ;
	    RECT 24.6000 68.8000 25.0000 69.2000 ;
	    RECT 24.6000 68.2000 24.9000 68.8000 ;
	    RECT 15.0000 67.8000 15.4000 68.2000 ;
	    RECT 18.2000 67.8000 18.6000 68.2000 ;
	    RECT 23.8000 67.8000 24.2000 68.2000 ;
	    RECT 24.6000 67.8000 25.0000 68.2000 ;
	    RECT 15.0000 67.2000 15.3000 67.8000 ;
	    RECT 4.6000 66.8000 5.0000 67.2000 ;
	    RECT 8.6000 67.1000 9.0000 67.2000 ;
	    RECT 9.4000 67.1000 9.8000 67.2000 ;
	    RECT 8.6000 66.8000 9.8000 67.1000 ;
	    RECT 12.6000 66.8000 13.0000 67.2000 ;
	    RECT 15.0000 66.8000 15.4000 67.2000 ;
	    RECT 16.6000 66.8000 17.0000 67.2000 ;
	    RECT 18.2000 67.1000 18.6000 67.2000 ;
	    RECT 19.0000 67.1000 19.4000 67.2000 ;
	    RECT 18.2000 66.8000 19.4000 67.1000 ;
	    RECT 21.4000 66.8000 21.8000 67.2000 ;
	    RECT 22.2000 66.8000 22.6000 67.2000 ;
	    RECT 4.6000 66.2000 4.9000 66.8000 ;
	    RECT 12.6000 66.2000 12.9000 66.8000 ;
	    RECT 2.2000 65.8000 2.6000 66.2000 ;
	    RECT 3.8000 65.8000 4.2000 66.2000 ;
	    RECT 4.6000 65.8000 5.0000 66.2000 ;
	    RECT 7.8000 65.8000 8.2000 66.2000 ;
	    RECT 8.6000 66.1000 9.0000 66.2000 ;
	    RECT 9.4000 66.1000 9.8000 66.2000 ;
	    RECT 8.6000 65.8000 9.8000 66.1000 ;
	    RECT 11.8000 65.8000 12.2000 66.2000 ;
	    RECT 12.6000 65.8000 13.0000 66.2000 ;
	    RECT 15.8000 65.8000 16.2000 66.2000 ;
	    RECT 2.2000 65.2000 2.5000 65.8000 ;
	    RECT 3.8000 65.2000 4.1000 65.8000 ;
	    RECT 7.8000 65.2000 8.1000 65.8000 ;
	    RECT 2.2000 64.8000 2.6000 65.2000 ;
	    RECT 3.8000 64.8000 4.2000 65.2000 ;
	    RECT 7.8000 64.8000 8.2000 65.2000 ;
	    RECT 9.4000 65.1000 9.8000 65.2000 ;
	    RECT 10.2000 65.1000 10.6000 65.2000 ;
	    RECT 9.4000 64.8000 10.6000 65.1000 ;
	    RECT 11.8000 64.2000 12.1000 65.8000 ;
	    RECT 11.8000 63.8000 12.2000 64.2000 ;
	    RECT 8.6000 62.8000 9.0000 63.2000 ;
	    RECT 8.6000 59.2000 8.9000 62.8000 ;
	    RECT 8.6000 58.8000 9.0000 59.2000 ;
	    RECT 3.8000 56.8000 4.2000 57.2000 ;
	    RECT 1.3000 55.9000 1.7000 56.3000 ;
	    RECT 3.8000 56.2000 4.1000 56.8000 ;
	    RECT 1.3000 53.5000 1.6000 55.9000 ;
	    RECT 3.8000 55.8000 4.2000 56.2000 ;
	    RECT 4.6000 55.9000 5.0000 56.3000 ;
	    RECT 2.6000 54.2000 3.0000 54.3000 ;
	    RECT 4.7000 54.2000 5.0000 55.9000 ;
	    RECT 11.0000 56.1000 11.4000 56.2000 ;
	    RECT 11.8000 56.1000 12.2000 56.2000 ;
	    RECT 11.0000 55.8000 12.2000 56.1000 ;
	    RECT 12.6000 55.2000 12.9000 65.8000 ;
	    RECT 15.8000 65.2000 16.1000 65.8000 ;
	    RECT 15.8000 64.8000 16.2000 65.2000 ;
	    RECT 16.6000 64.1000 16.9000 66.8000 ;
	    RECT 19.8000 66.1000 20.2000 66.2000 ;
	    RECT 20.6000 66.1000 21.0000 66.2000 ;
	    RECT 19.8000 65.8000 21.0000 66.1000 ;
	    RECT 19.0000 65.1000 19.4000 65.2000 ;
	    RECT 19.8000 65.1000 20.2000 65.2000 ;
	    RECT 19.0000 64.8000 20.2000 65.1000 ;
	    RECT 15.8000 63.8000 16.9000 64.1000 ;
	    RECT 19.0000 63.8000 19.4000 64.2000 ;
	    RECT 13.4000 55.8000 13.8000 56.2000 ;
	    RECT 13.4000 55.2000 13.7000 55.8000 ;
	    RECT 11.0000 55.1000 11.4000 55.2000 ;
	    RECT 11.8000 55.1000 12.2000 55.2000 ;
	    RECT 11.0000 54.8000 12.2000 55.1000 ;
	    RECT 12.6000 54.8000 13.0000 55.2000 ;
	    RECT 13.4000 54.8000 13.8000 55.2000 ;
	    RECT 2.6000 53.9000 5.0000 54.2000 ;
	    RECT 4.7000 53.5000 5.0000 53.9000 ;
	    RECT 1.3000 53.1000 1.7000 53.5000 ;
	    RECT 4.6000 53.1000 5.0000 53.5000 ;
	    RECT 14.2000 53.8000 14.6000 54.2000 ;
	    RECT 10.2000 52.8000 10.6000 53.2000 ;
	    RECT 3.0000 49.1000 3.4000 49.2000 ;
	    RECT 3.8000 49.1000 4.2000 49.2000 ;
	    RECT 3.0000 48.8000 4.2000 49.1000 ;
	    RECT 8.6000 48.8000 9.0000 49.2000 ;
	    RECT 8.6000 48.2000 8.9000 48.8000 ;
	    RECT 1.4000 47.5000 1.8000 47.9000 ;
	    RECT 4.5000 47.8000 4.9000 47.9000 ;
	    RECT 8.6000 47.8000 9.0000 48.2000 ;
	    RECT 2.1000 47.5000 4.9000 47.8000 ;
	    RECT 1.4000 47.1000 1.7000 47.5000 ;
	    RECT 2.1000 47.4000 2.5000 47.5000 ;
	    RECT 3.8000 47.4000 4.2000 47.5000 ;
	    RECT 1.4000 46.8000 4.2000 47.1000 ;
	    RECT 1.4000 45.1000 1.7000 46.8000 ;
	    RECT 3.9000 46.1000 4.2000 46.8000 ;
	    RECT 3.9000 45.7000 4.3000 46.1000 ;
	    RECT 4.6000 45.1000 4.9000 47.5000 ;
	    RECT 10.2000 47.2000 10.5000 52.8000 ;
	    RECT 14.2000 49.2000 14.5000 53.8000 ;
	    RECT 15.8000 49.2000 16.1000 63.8000 ;
	    RECT 19.0000 59.2000 19.3000 63.8000 ;
	    RECT 19.0000 58.8000 19.4000 59.2000 ;
	    RECT 16.6000 54.8000 17.0000 55.2000 ;
	    RECT 17.4000 55.1000 17.8000 55.2000 ;
	    RECT 18.2000 55.1000 18.6000 55.2000 ;
	    RECT 17.4000 54.8000 18.6000 55.1000 ;
	    RECT 16.6000 54.2000 16.9000 54.8000 ;
	    RECT 16.6000 53.8000 17.0000 54.2000 ;
	    RECT 20.6000 53.8000 21.0000 54.2000 ;
	    RECT 20.6000 52.2000 20.9000 53.8000 ;
	    RECT 20.6000 51.8000 21.0000 52.2000 ;
	    RECT 21.4000 49.2000 21.7000 66.8000 ;
	    RECT 22.2000 66.2000 22.5000 66.8000 ;
	    RECT 26.2000 66.2000 26.5000 73.8000 ;
	    RECT 27.8000 72.8000 28.2000 73.2000 ;
	    RECT 27.8000 69.2000 28.1000 72.8000 ;
	    RECT 29.4000 69.2000 29.7000 73.8000 ;
	    RECT 36.6000 73.5000 36.9000 73.9000 ;
	    RECT 37.3000 73.5000 37.7000 73.6000 ;
	    RECT 39.0000 73.5000 39.4000 73.6000 ;
	    RECT 39.8000 73.5000 40.1000 75.9000 ;
	    RECT 43.0000 75.8000 43.4000 76.2000 ;
	    RECT 44.6000 75.8000 45.0000 76.2000 ;
	    RECT 41.4000 74.1000 41.8000 74.2000 ;
	    RECT 42.2000 74.1000 42.6000 74.2000 ;
	    RECT 41.4000 73.8000 42.6000 74.1000 ;
	    RECT 33.4000 72.8000 33.8000 73.2000 ;
	    RECT 36.6000 73.1000 37.0000 73.5000 ;
	    RECT 37.3000 73.2000 40.1000 73.5000 ;
	    RECT 39.7000 73.1000 40.1000 73.2000 ;
	    RECT 41.4000 72.8000 41.8000 73.2000 ;
	    RECT 33.4000 72.2000 33.7000 72.8000 ;
	    RECT 31.0000 72.1000 31.4000 72.2000 ;
	    RECT 31.8000 72.1000 32.2000 72.2000 ;
	    RECT 31.0000 71.8000 32.2000 72.1000 ;
	    RECT 33.4000 71.8000 33.8000 72.2000 ;
	    RECT 37.4000 72.1000 37.8000 72.2000 ;
	    RECT 38.2000 72.1000 38.6000 72.2000 ;
	    RECT 37.4000 71.8000 38.6000 72.1000 ;
	    RECT 37.4000 70.8000 37.8000 71.2000 ;
	    RECT 31.0000 69.8000 31.4000 70.2000 ;
	    RECT 31.0000 69.2000 31.3000 69.8000 ;
	    RECT 37.4000 69.2000 37.7000 70.8000 ;
	    RECT 27.0000 68.8000 27.4000 69.2000 ;
	    RECT 27.8000 68.8000 28.2000 69.2000 ;
	    RECT 29.4000 68.8000 29.8000 69.2000 ;
	    RECT 31.0000 68.8000 31.4000 69.2000 ;
	    RECT 37.4000 68.8000 37.8000 69.2000 ;
	    RECT 27.0000 68.2000 27.3000 68.8000 ;
	    RECT 41.4000 68.2000 41.7000 72.8000 ;
	    RECT 43.0000 71.2000 43.3000 75.8000 ;
	    RECT 44.6000 75.1000 45.0000 75.2000 ;
	    RECT 45.4000 75.1000 45.8000 75.2000 ;
	    RECT 44.6000 74.8000 45.8000 75.1000 ;
	    RECT 47.0000 74.8000 47.4000 75.2000 ;
	    RECT 47.0000 74.2000 47.3000 74.8000 ;
	    RECT 44.6000 74.1000 45.0000 74.2000 ;
	    RECT 45.4000 74.1000 45.8000 74.2000 ;
	    RECT 44.6000 73.8000 45.8000 74.1000 ;
	    RECT 47.0000 73.8000 47.4000 74.2000 ;
	    RECT 46.2000 72.8000 46.6000 73.2000 ;
	    RECT 43.0000 70.8000 43.4000 71.2000 ;
	    RECT 43.0000 68.8000 43.4000 69.2000 ;
	    RECT 27.0000 67.8000 27.4000 68.2000 ;
	    RECT 28.6000 67.8000 29.0000 68.2000 ;
	    RECT 33.4000 67.8000 33.8000 68.2000 ;
	    RECT 36.6000 67.8000 37.0000 68.2000 ;
	    RECT 39.0000 67.8000 39.4000 68.2000 ;
	    RECT 41.4000 67.8000 41.8000 68.2000 ;
	    RECT 42.2000 67.8000 42.6000 68.2000 ;
	    RECT 28.6000 67.2000 28.9000 67.8000 ;
	    RECT 28.6000 66.8000 29.0000 67.2000 ;
	    RECT 31.0000 66.8000 31.4000 67.2000 ;
	    RECT 22.2000 65.8000 22.6000 66.2000 ;
	    RECT 24.6000 66.1000 25.0000 66.2000 ;
	    RECT 25.4000 66.1000 25.8000 66.2000 ;
	    RECT 24.6000 65.8000 25.8000 66.1000 ;
	    RECT 26.2000 65.8000 26.6000 66.2000 ;
	    RECT 28.6000 66.1000 29.0000 66.2000 ;
	    RECT 29.4000 66.1000 29.8000 66.2000 ;
	    RECT 28.6000 65.8000 29.8000 66.1000 ;
	    RECT 26.2000 64.8000 26.6000 65.2000 ;
	    RECT 26.2000 59.2000 26.5000 64.8000 ;
	    RECT 26.2000 58.8000 26.6000 59.2000 ;
	    RECT 29.4000 57.8000 29.8000 58.2000 ;
	    RECT 22.2000 55.8000 22.6000 56.2000 ;
	    RECT 25.3000 55.9000 25.7000 56.3000 ;
	    RECT 28.6000 55.9000 29.0000 56.3000 ;
	    RECT 22.2000 55.2000 22.5000 55.8000 ;
	    RECT 22.2000 54.8000 22.6000 55.2000 ;
	    RECT 25.3000 53.5000 25.6000 55.9000 ;
	    RECT 26.6000 54.2000 27.0000 54.3000 ;
	    RECT 28.7000 54.2000 29.0000 55.9000 ;
	    RECT 26.6000 53.9000 29.0000 54.2000 ;
	    RECT 28.7000 53.5000 29.0000 53.9000 ;
	    RECT 25.3000 53.1000 25.7000 53.5000 ;
	    RECT 28.6000 53.1000 29.0000 53.5000 ;
	    RECT 29.4000 54.2000 29.7000 57.8000 ;
	    RECT 30.2000 56.8000 30.6000 57.2000 ;
	    RECT 30.2000 56.2000 30.5000 56.8000 ;
	    RECT 30.2000 55.8000 30.6000 56.2000 ;
	    RECT 31.0000 55.2000 31.3000 66.8000 ;
	    RECT 31.8000 64.8000 32.2000 65.2000 ;
	    RECT 31.8000 64.2000 32.1000 64.8000 ;
	    RECT 31.8000 63.8000 32.2000 64.2000 ;
	    RECT 33.4000 59.2000 33.7000 67.8000 ;
	    RECT 36.6000 67.2000 36.9000 67.8000 ;
	    RECT 34.2000 66.8000 34.6000 67.2000 ;
	    RECT 35.8000 66.8000 36.2000 67.2000 ;
	    RECT 36.6000 66.8000 37.0000 67.2000 ;
	    RECT 34.2000 66.2000 34.5000 66.8000 ;
	    RECT 35.8000 66.2000 36.1000 66.8000 ;
	    RECT 39.0000 66.2000 39.3000 67.8000 ;
	    RECT 42.2000 67.2000 42.5000 67.8000 ;
	    RECT 39.8000 66.8000 40.2000 67.2000 ;
	    RECT 42.2000 66.8000 42.6000 67.2000 ;
	    RECT 34.2000 65.8000 34.6000 66.2000 ;
	    RECT 35.8000 65.8000 36.2000 66.2000 ;
	    RECT 37.4000 66.1000 37.8000 66.2000 ;
	    RECT 38.2000 66.1000 38.6000 66.2000 ;
	    RECT 37.4000 65.8000 38.6000 66.1000 ;
	    RECT 39.0000 65.8000 39.4000 66.2000 ;
	    RECT 35.8000 64.8000 36.2000 65.2000 ;
	    RECT 35.8000 64.2000 36.1000 64.8000 ;
	    RECT 39.8000 64.2000 40.1000 66.8000 ;
	    RECT 42.2000 65.8000 42.6000 66.2000 ;
	    RECT 42.2000 65.2000 42.5000 65.8000 ;
	    RECT 42.2000 64.8000 42.6000 65.2000 ;
	    RECT 43.0000 64.2000 43.3000 68.8000 ;
	    RECT 45.4000 67.8000 45.8000 68.2000 ;
	    RECT 45.4000 67.2000 45.7000 67.8000 ;
	    RECT 45.4000 66.8000 45.8000 67.2000 ;
	    RECT 45.4000 65.8000 45.8000 66.2000 ;
	    RECT 45.4000 65.2000 45.7000 65.8000 ;
	    RECT 43.8000 65.1000 44.2000 65.2000 ;
	    RECT 44.6000 65.1000 45.0000 65.2000 ;
	    RECT 43.8000 64.8000 45.0000 65.1000 ;
	    RECT 45.4000 64.8000 45.8000 65.2000 ;
	    RECT 43.8000 64.2000 44.1000 64.8000 ;
	    RECT 35.8000 63.8000 36.2000 64.2000 ;
	    RECT 39.8000 63.8000 40.2000 64.2000 ;
	    RECT 43.0000 63.8000 43.4000 64.2000 ;
	    RECT 43.8000 63.8000 44.2000 64.2000 ;
	    RECT 33.4000 58.8000 33.8000 59.2000 ;
	    RECT 43.0000 59.1000 43.4000 59.2000 ;
	    RECT 43.8000 59.1000 44.2000 59.2000 ;
	    RECT 43.0000 58.8000 44.2000 59.1000 ;
	    RECT 31.0000 54.8000 31.4000 55.2000 ;
	    RECT 31.8000 54.8000 32.2000 55.2000 ;
	    RECT 32.6000 54.8000 33.0000 55.2000 ;
	    RECT 37.4000 55.1000 37.8000 55.2000 ;
	    RECT 38.2000 55.1000 38.6000 55.2000 ;
	    RECT 37.4000 54.8000 38.6000 55.1000 ;
	    RECT 39.8000 54.8000 40.2000 55.2000 ;
	    RECT 40.6000 54.8000 41.0000 55.2000 ;
	    RECT 29.4000 53.8000 29.8000 54.2000 ;
	    RECT 25.4000 51.8000 25.8000 52.2000 ;
	    RECT 25.4000 49.2000 25.7000 51.8000 ;
	    RECT 14.2000 48.8000 14.6000 49.2000 ;
	    RECT 15.8000 48.8000 16.2000 49.2000 ;
	    RECT 21.4000 48.8000 21.8000 49.2000 ;
	    RECT 25.4000 48.8000 25.8000 49.2000 ;
	    RECT 29.4000 48.2000 29.7000 53.8000 ;
	    RECT 31.8000 52.2000 32.1000 54.8000 ;
	    RECT 32.6000 54.2000 32.9000 54.8000 ;
	    RECT 32.6000 53.8000 33.0000 54.2000 ;
	    RECT 36.6000 54.1000 37.0000 54.2000 ;
	    RECT 37.4000 54.1000 37.8000 54.2000 ;
	    RECT 36.6000 53.8000 37.8000 54.1000 ;
	    RECT 38.2000 53.8000 38.6000 54.2000 ;
	    RECT 35.0000 53.1000 35.4000 53.2000 ;
	    RECT 35.8000 53.1000 36.2000 53.2000 ;
	    RECT 35.0000 52.8000 36.2000 53.1000 ;
	    RECT 31.8000 51.8000 32.2000 52.2000 ;
	    RECT 36.6000 48.2000 36.9000 53.8000 ;
	    RECT 38.2000 53.2000 38.5000 53.8000 ;
	    RECT 38.2000 52.8000 38.6000 53.2000 ;
	    RECT 39.0000 52.8000 39.4000 53.2000 ;
	    RECT 39.0000 52.2000 39.3000 52.8000 ;
	    RECT 39.0000 51.8000 39.4000 52.2000 ;
	    RECT 39.8000 49.2000 40.1000 54.8000 ;
	    RECT 40.6000 50.2000 40.9000 54.8000 ;
	    RECT 45.4000 52.1000 45.8000 57.9000 ;
	    RECT 40.6000 49.8000 41.0000 50.2000 ;
	    RECT 42.2000 49.8000 42.6000 50.2000 ;
	    RECT 42.2000 49.2000 42.5000 49.8000 ;
	    RECT 39.8000 48.8000 40.2000 49.2000 ;
	    RECT 42.2000 48.8000 42.6000 49.2000 ;
	    RECT 43.0000 49.1000 43.4000 49.2000 ;
	    RECT 43.8000 49.1000 44.2000 49.2000 ;
	    RECT 43.0000 48.8000 44.2000 49.1000 ;
	    RECT 18.9000 47.5000 19.3000 47.9000 ;
	    RECT 22.2000 47.5000 22.6000 47.9000 ;
	    RECT 29.4000 47.8000 29.8000 48.2000 ;
	    RECT 30.2000 48.1000 30.6000 48.2000 ;
	    RECT 31.0000 48.1000 31.4000 48.2000 ;
	    RECT 30.2000 47.8000 31.4000 48.1000 ;
	    RECT 10.2000 46.8000 10.6000 47.2000 ;
	    RECT 17.4000 46.8000 17.8000 47.2000 ;
	    RECT 10.2000 46.2000 10.5000 46.8000 ;
	    RECT 17.4000 46.2000 17.7000 46.8000 ;
	    RECT 6.2000 46.1000 6.6000 46.2000 ;
	    RECT 7.0000 46.1000 7.4000 46.2000 ;
	    RECT 6.2000 45.8000 7.4000 46.1000 ;
	    RECT 9.4000 45.8000 9.8000 46.2000 ;
	    RECT 10.2000 45.8000 10.6000 46.2000 ;
	    RECT 17.4000 45.8000 17.8000 46.2000 ;
	    RECT 1.4000 44.7000 1.8000 45.1000 ;
	    RECT 4.5000 44.7000 4.9000 45.1000 ;
	    RECT 9.4000 45.2000 9.7000 45.8000 ;
	    RECT 9.4000 44.8000 9.8000 45.2000 ;
	    RECT 15.0000 45.1000 15.4000 45.2000 ;
	    RECT 15.8000 45.1000 16.2000 45.2000 ;
	    RECT 15.0000 44.8000 16.2000 45.1000 ;
	    RECT 18.9000 45.1000 19.2000 47.5000 ;
	    RECT 22.3000 47.1000 22.6000 47.5000 ;
	    RECT 32.5000 47.5000 32.9000 47.9000 ;
	    RECT 35.8000 47.5000 36.2000 47.9000 ;
	    RECT 20.2000 46.8000 22.6000 47.1000 ;
	    RECT 27.0000 47.1000 27.4000 47.2000 ;
	    RECT 27.8000 47.1000 28.2000 47.2000 ;
	    RECT 27.0000 46.8000 28.2000 47.1000 ;
	    RECT 20.2000 46.7000 20.6000 46.8000 ;
	    RECT 19.8000 45.8000 20.2000 46.2000 ;
	    RECT 18.9000 44.7000 19.3000 45.1000 ;
	    RECT 19.8000 39.2000 20.1000 45.8000 ;
	    RECT 22.3000 45.1000 22.6000 46.8000 ;
	    RECT 22.2000 44.7000 22.6000 45.1000 ;
	    RECT 27.0000 45.8000 27.4000 46.2000 ;
	    RECT 19.8000 38.8000 20.2000 39.2000 ;
	    RECT 3.0000 37.1000 3.4000 37.2000 ;
	    RECT 3.8000 37.1000 4.2000 37.2000 ;
	    RECT 3.0000 36.8000 4.2000 37.1000 ;
	    RECT 1.3000 35.9000 1.7000 36.3000 ;
	    RECT 4.6000 35.9000 5.0000 36.3000 ;
	    RECT 1.3000 33.5000 1.6000 35.9000 ;
	    RECT 2.6000 34.2000 3.0000 34.3000 ;
	    RECT 4.7000 34.2000 5.0000 35.9000 ;
	    RECT 2.6000 33.9000 5.0000 34.2000 ;
	    RECT 4.7000 33.5000 5.0000 33.9000 ;
	    RECT 1.3000 33.1000 1.7000 33.5000 ;
	    RECT 4.6000 33.1000 5.0000 33.5000 ;
	    RECT 7.1000 35.9000 7.5000 36.3000 ;
	    RECT 10.2000 35.9000 10.6000 36.3000 ;
	    RECT 27.0000 36.2000 27.3000 45.8000 ;
	    RECT 32.5000 45.1000 32.8000 47.5000 ;
	    RECT 35.9000 47.1000 36.2000 47.5000 ;
	    RECT 33.8000 46.8000 36.2000 47.1000 ;
	    RECT 36.6000 47.8000 37.0000 48.2000 ;
	    RECT 37.4000 48.1000 37.8000 48.2000 ;
	    RECT 38.2000 48.1000 38.6000 48.2000 ;
	    RECT 37.4000 47.8000 38.6000 48.1000 ;
	    RECT 36.6000 47.2000 36.9000 47.8000 ;
	    RECT 36.6000 46.8000 37.0000 47.2000 ;
	    RECT 33.8000 46.7000 34.2000 46.8000 ;
	    RECT 35.9000 45.1000 36.2000 46.8000 ;
	    RECT 32.5000 44.7000 32.9000 45.1000 ;
	    RECT 35.8000 44.7000 36.2000 45.1000 ;
	    RECT 31.8000 43.8000 32.2000 44.2000 ;
	    RECT 31.8000 39.2000 32.1000 43.8000 ;
	    RECT 45.4000 43.1000 45.8000 48.9000 ;
	    RECT 33.4000 41.8000 33.8000 42.2000 ;
	    RECT 37.4000 41.8000 37.8000 42.2000 ;
	    RECT 31.8000 38.8000 32.2000 39.2000 ;
	    RECT 27.8000 36.8000 28.2000 37.2000 ;
	    RECT 27.8000 36.2000 28.1000 36.8000 ;
	    RECT 33.4000 36.2000 33.7000 41.8000 ;
	    RECT 7.1000 33.5000 7.4000 35.9000 ;
	    RECT 7.7000 34.9000 8.1000 35.3000 ;
	    RECT 7.8000 34.2000 8.1000 34.9000 ;
	    RECT 10.3000 34.2000 10.6000 35.9000 ;
	    RECT 15.0000 35.8000 15.4000 36.2000 ;
	    RECT 18.2000 35.8000 18.6000 36.2000 ;
	    RECT 19.8000 35.8000 20.2000 36.2000 ;
	    RECT 27.0000 35.8000 27.4000 36.2000 ;
	    RECT 27.8000 35.8000 28.2000 36.2000 ;
	    RECT 30.2000 35.8000 30.6000 36.2000 ;
	    RECT 33.4000 35.8000 33.8000 36.2000 ;
	    RECT 36.6000 35.9000 37.0000 36.3000 ;
	    RECT 37.4000 36.2000 37.7000 41.8000 ;
	    RECT 46.2000 39.2000 46.5000 72.8000 ;
	    RECT 47.0000 68.2000 47.3000 73.8000 ;
	    RECT 47.8000 73.2000 48.1000 82.8000 ;
	    RECT 51.8000 81.8000 52.2000 82.2000 ;
	    RECT 51.0000 75.8000 51.4000 76.2000 ;
	    RECT 51.0000 75.2000 51.3000 75.8000 ;
	    RECT 49.4000 74.8000 49.8000 75.2000 ;
	    RECT 51.0000 74.8000 51.4000 75.2000 ;
	    RECT 49.4000 74.2000 49.7000 74.8000 ;
	    RECT 51.8000 74.2000 52.1000 81.8000 ;
	    RECT 52.6000 78.8000 53.0000 79.2000 ;
	    RECT 49.4000 73.8000 49.8000 74.2000 ;
	    RECT 51.8000 73.8000 52.2000 74.2000 ;
	    RECT 47.8000 72.8000 48.2000 73.2000 ;
	    RECT 51.0000 72.8000 51.4000 73.2000 ;
	    RECT 47.8000 71.8000 48.2000 72.2000 ;
	    RECT 49.4000 71.8000 49.8000 72.2000 ;
	    RECT 47.8000 69.2000 48.1000 71.8000 ;
	    RECT 47.8000 68.8000 48.2000 69.2000 ;
	    RECT 47.0000 67.8000 47.4000 68.2000 ;
	    RECT 47.8000 67.8000 48.2000 68.2000 ;
	    RECT 47.0000 49.2000 47.3000 67.8000 ;
	    RECT 47.8000 67.2000 48.1000 67.8000 ;
	    RECT 47.8000 66.8000 48.2000 67.2000 ;
	    RECT 49.4000 66.2000 49.7000 71.8000 ;
	    RECT 49.4000 65.8000 49.8000 66.2000 ;
	    RECT 50.2000 65.1000 50.6000 67.9000 ;
	    RECT 51.0000 66.2000 51.3000 72.8000 ;
	    RECT 51.8000 72.2000 52.1000 73.8000 ;
	    RECT 51.8000 71.8000 52.2000 72.2000 ;
	    RECT 51.0000 65.8000 51.4000 66.2000 ;
	    RECT 51.8000 63.1000 52.2000 68.9000 ;
	    RECT 52.6000 68.2000 52.9000 78.8000 ;
	    RECT 53.4000 76.1000 53.7000 88.8000 ;
	    RECT 54.2000 85.2000 54.5000 91.8000 ;
	    RECT 57.4000 90.2000 57.7000 91.8000 ;
	    RECT 57.4000 89.8000 57.8000 90.2000 ;
	    RECT 57.4000 88.8000 57.8000 89.2000 ;
	    RECT 57.4000 88.2000 57.7000 88.8000 ;
	    RECT 55.8000 88.1000 56.2000 88.2000 ;
	    RECT 55.8000 87.8000 56.9000 88.1000 ;
	    RECT 57.4000 87.8000 57.8000 88.2000 ;
	    RECT 55.8000 86.8000 56.2000 87.2000 ;
	    RECT 54.2000 84.8000 54.6000 85.2000 ;
	    RECT 55.8000 77.2000 56.1000 86.8000 ;
	    RECT 56.6000 85.2000 56.9000 87.8000 ;
	    RECT 57.4000 87.1000 57.8000 87.2000 ;
	    RECT 58.2000 87.1000 58.6000 87.2000 ;
	    RECT 57.4000 86.8000 58.6000 87.1000 ;
	    RECT 59.8000 86.2000 60.1000 91.8000 ;
	    RECT 60.6000 89.2000 60.9000 93.8000 ;
	    RECT 62.2000 93.1000 62.6000 95.9000 ;
	    RECT 63.8000 92.1000 64.2000 97.9000 ;
	    RECT 66.2000 97.8000 66.6000 98.2000 ;
	    RECT 64.6000 95.0000 65.0000 95.1000 ;
	    RECT 65.4000 95.0000 65.8000 95.1000 ;
	    RECT 64.6000 94.7000 65.8000 95.0000 ;
	    RECT 67.8000 94.8000 68.2000 95.2000 ;
	    RECT 60.6000 88.8000 61.0000 89.2000 ;
	    RECT 67.8000 88.2000 68.1000 94.8000 ;
	    RECT 68.6000 92.1000 69.0000 97.9000 ;
	    RECT 67.8000 87.8000 68.2000 88.2000 ;
	    RECT 63.0000 86.8000 63.4000 87.2000 ;
	    RECT 59.8000 85.8000 60.2000 86.2000 ;
	    RECT 62.2000 85.8000 62.6000 86.2000 ;
	    RECT 56.6000 84.8000 57.0000 85.2000 ;
	    RECT 58.2000 85.1000 58.6000 85.2000 ;
	    RECT 59.0000 85.1000 59.4000 85.2000 ;
	    RECT 58.2000 84.8000 59.4000 85.1000 ;
	    RECT 56.6000 83.2000 56.9000 84.8000 ;
	    RECT 56.6000 82.8000 57.0000 83.2000 ;
	    RECT 62.2000 82.2000 62.5000 85.8000 ;
	    RECT 63.0000 85.2000 63.3000 86.8000 ;
	    RECT 65.4000 85.8000 65.8000 86.2000 ;
	    RECT 63.0000 84.8000 63.4000 85.2000 ;
	    RECT 65.4000 84.2000 65.7000 85.8000 ;
	    RECT 64.6000 83.8000 65.0000 84.2000 ;
	    RECT 65.4000 83.8000 65.8000 84.2000 ;
	    RECT 62.2000 81.8000 62.6000 82.2000 ;
	    RECT 57.4000 79.1000 57.8000 79.2000 ;
	    RECT 58.2000 79.1000 58.6000 79.2000 ;
	    RECT 57.4000 78.8000 58.6000 79.1000 ;
	    RECT 55.8000 76.8000 56.2000 77.2000 ;
	    RECT 56.6000 76.8000 57.0000 77.2000 ;
	    RECT 59.8000 77.1000 60.2000 77.2000 ;
	    RECT 60.6000 77.1000 61.0000 77.2000 ;
	    RECT 59.8000 76.8000 61.0000 77.1000 ;
	    RECT 54.2000 76.1000 54.6000 76.2000 ;
	    RECT 53.4000 75.8000 54.6000 76.1000 ;
	    RECT 55.0000 75.8000 55.4000 76.2000 ;
	    RECT 54.2000 74.8000 54.6000 75.2000 ;
	    RECT 54.2000 74.2000 54.5000 74.8000 ;
	    RECT 54.2000 73.8000 54.6000 74.2000 ;
	    RECT 55.0000 68.2000 55.3000 75.8000 ;
	    RECT 55.8000 75.2000 56.1000 76.8000 ;
	    RECT 55.8000 74.8000 56.2000 75.2000 ;
	    RECT 55.8000 70.8000 56.2000 71.2000 ;
	    RECT 52.6000 67.8000 53.0000 68.2000 ;
	    RECT 55.0000 67.8000 55.4000 68.2000 ;
	    RECT 53.4000 66.8000 53.8000 67.2000 ;
	    RECT 53.4000 66.2000 53.7000 66.8000 ;
	    RECT 55.8000 66.2000 56.1000 70.8000 ;
	    RECT 56.6000 70.2000 56.9000 76.8000 ;
	    RECT 62.2000 72.1000 62.6000 77.9000 ;
	    RECT 64.6000 74.1000 64.9000 83.8000 ;
	    RECT 69.4000 83.1000 69.8000 88.9000 ;
	    RECT 71.0000 88.2000 71.3000 105.8000 ;
	    RECT 72.6000 97.8000 73.0000 98.2000 ;
	    RECT 72.6000 96.2000 72.9000 97.8000 ;
	    RECT 73.4000 97.2000 73.7000 116.8000 ;
	    RECT 75.0000 115.1000 75.4000 115.2000 ;
	    RECT 75.8000 115.1000 76.2000 115.2000 ;
	    RECT 75.0000 114.8000 76.2000 115.1000 ;
	    RECT 77.4000 111.8000 77.8000 112.2000 ;
	    RECT 77.4000 110.2000 77.7000 111.8000 ;
	    RECT 77.4000 109.8000 77.8000 110.2000 ;
	    RECT 74.2000 105.9000 74.6000 106.3000 ;
	    RECT 74.2000 105.2000 74.5000 105.9000 ;
	    RECT 74.2000 104.8000 74.6000 105.2000 ;
	    RECT 75.0000 103.1000 75.4000 108.9000 ;
	    RECT 78.2000 108.2000 78.5000 127.8000 ;
	    RECT 79.0000 127.2000 79.3000 127.8000 ;
	    RECT 79.0000 126.8000 79.4000 127.2000 ;
	    RECT 79.8000 126.1000 80.2000 126.2000 ;
	    RECT 80.6000 126.1000 81.0000 126.2000 ;
	    RECT 79.8000 125.8000 81.0000 126.1000 ;
	    RECT 81.4000 124.8000 81.8000 125.2000 ;
	    RECT 81.4000 124.2000 81.7000 124.8000 ;
	    RECT 81.4000 123.8000 81.8000 124.2000 ;
	    RECT 79.8000 112.1000 80.2000 117.9000 ;
	    RECT 81.4000 112.2000 81.7000 123.8000 ;
	    RECT 82.2000 121.8000 82.6000 122.2000 ;
	    RECT 81.4000 111.8000 81.8000 112.2000 ;
	    RECT 77.4000 108.1000 77.8000 108.2000 ;
	    RECT 78.2000 108.1000 78.6000 108.2000 ;
	    RECT 76.6000 105.1000 77.0000 107.9000 ;
	    RECT 77.4000 107.8000 78.6000 108.1000 ;
	    RECT 77.4000 106.8000 77.8000 107.2000 ;
	    RECT 77.4000 106.2000 77.7000 106.8000 ;
	    RECT 82.2000 106.2000 82.5000 121.8000 ;
	    RECT 83.0000 116.2000 83.3000 133.8000 ;
	    RECT 83.8000 133.1000 84.2000 135.9000 ;
	    RECT 87.0000 135.2000 87.3000 141.8000 ;
	    RECT 88.6000 139.2000 88.9000 143.8000 ;
	    RECT 91.8000 142.1000 92.1000 145.8000 ;
	    RECT 92.6000 143.1000 93.0000 148.9000 ;
	    RECT 93.4000 148.8000 93.8000 149.2000 ;
	    RECT 94.2000 149.1000 94.6000 149.2000 ;
	    RECT 95.0000 149.1000 95.4000 149.2000 ;
	    RECT 94.2000 148.8000 95.4000 149.1000 ;
	    RECT 95.0000 147.2000 95.3000 148.8000 ;
	    RECT 95.8000 148.2000 96.1000 152.8000 ;
	    RECT 98.2000 152.2000 98.5000 152.8000 ;
	    RECT 96.6000 151.8000 97.0000 152.2000 ;
	    RECT 98.2000 151.8000 98.6000 152.2000 ;
	    RECT 95.8000 147.8000 96.2000 148.2000 ;
	    RECT 95.0000 146.8000 95.4000 147.2000 ;
	    RECT 95.8000 146.8000 96.2000 147.2000 ;
	    RECT 95.8000 146.2000 96.1000 146.8000 ;
	    RECT 95.8000 145.8000 96.2000 146.2000 ;
	    RECT 91.8000 141.8000 92.9000 142.1000 ;
	    RECT 92.6000 139.2000 92.9000 141.8000 ;
	    RECT 95.0000 141.8000 95.4000 142.2000 ;
	    RECT 88.6000 138.8000 89.0000 139.2000 ;
	    RECT 92.6000 138.8000 93.0000 139.2000 ;
	    RECT 87.8000 137.8000 88.2000 138.2000 ;
	    RECT 87.0000 134.8000 87.4000 135.2000 ;
	    RECT 87.8000 133.2000 88.1000 137.8000 ;
	    RECT 92.6000 134.8000 93.0000 135.2000 ;
	    RECT 87.8000 132.8000 88.2000 133.2000 ;
	    RECT 92.6000 129.2000 92.9000 134.8000 ;
	    RECT 95.0000 133.2000 95.3000 141.8000 ;
	    RECT 95.0000 132.8000 95.4000 133.2000 ;
	    RECT 92.6000 128.8000 93.0000 129.2000 ;
	    RECT 91.8000 127.8000 92.2000 128.2000 ;
	    RECT 93.4000 127.8000 93.8000 128.2000 ;
	    RECT 83.8000 126.8000 84.2000 127.2000 ;
	    RECT 83.8000 126.2000 84.1000 126.8000 ;
	    RECT 83.8000 125.8000 84.2000 126.2000 ;
	    RECT 84.6000 125.8000 85.0000 126.2000 ;
	    RECT 83.0000 115.8000 83.4000 116.2000 ;
	    RECT 83.0000 114.8000 83.4000 115.2000 ;
	    RECT 83.0000 111.2000 83.3000 114.8000 ;
	    RECT 83.0000 110.8000 83.4000 111.2000 ;
	    RECT 83.8000 110.1000 84.1000 125.8000 ;
	    RECT 84.6000 122.2000 84.9000 125.8000 ;
	    RECT 91.8000 122.2000 92.1000 127.8000 ;
	    RECT 93.4000 127.2000 93.7000 127.8000 ;
	    RECT 93.4000 126.8000 93.8000 127.2000 ;
	    RECT 96.6000 127.1000 96.9000 151.8000 ;
	    RECT 99.8000 149.2000 100.1000 152.8000 ;
	    RECT 99.8000 148.8000 100.2000 149.2000 ;
	    RECT 102.2000 148.2000 102.5000 152.8000 ;
	    RECT 102.2000 147.8000 102.6000 148.2000 ;
	    RECT 99.8000 146.8000 100.2000 147.2000 ;
	    RECT 99.8000 146.2000 100.1000 146.8000 ;
	    RECT 99.8000 145.8000 100.2000 146.2000 ;
	    RECT 97.4000 145.1000 97.8000 145.2000 ;
	    RECT 98.2000 145.1000 98.6000 145.2000 ;
	    RECT 97.4000 144.8000 98.6000 145.1000 ;
	    RECT 102.2000 144.2000 102.5000 147.8000 ;
	    RECT 103.0000 145.2000 103.3000 152.8000 ;
	    RECT 111.8000 152.2000 112.1000 152.8000 ;
	    RECT 106.2000 151.8000 106.6000 152.2000 ;
	    RECT 107.8000 152.1000 108.2000 152.2000 ;
	    RECT 108.6000 152.1000 109.0000 152.2000 ;
	    RECT 107.8000 151.8000 109.0000 152.1000 ;
	    RECT 111.8000 151.8000 112.2000 152.2000 ;
	    RECT 114.2000 152.1000 114.6000 157.9000 ;
	    RECT 117.4000 155.8000 117.8000 156.2000 ;
	    RECT 117.4000 155.2000 117.7000 155.8000 ;
	    RECT 117.4000 154.8000 117.8000 155.2000 ;
	    RECT 119.0000 152.1000 119.4000 157.9000 ;
	    RECT 119.8000 153.8000 120.2000 154.2000 ;
	    RECT 119.8000 153.2000 120.1000 153.8000 ;
	    RECT 119.8000 152.8000 120.2000 153.2000 ;
	    RECT 120.6000 153.1000 121.0000 155.9000 ;
	    RECT 123.0000 154.8000 123.4000 155.2000 ;
	    RECT 104.6000 148.1000 105.0000 148.2000 ;
	    RECT 105.4000 148.1000 105.8000 148.2000 ;
	    RECT 104.6000 147.8000 105.8000 148.1000 ;
	    RECT 103.8000 146.1000 104.2000 146.2000 ;
	    RECT 104.6000 146.1000 105.0000 146.2000 ;
	    RECT 103.8000 145.8000 105.0000 146.1000 ;
	    RECT 106.2000 145.2000 106.5000 151.8000 ;
	    RECT 111.8000 150.2000 112.1000 151.8000 ;
	    RECT 111.8000 149.8000 112.2000 150.2000 ;
	    RECT 115.0000 149.8000 115.4000 150.2000 ;
	    RECT 111.8000 148.8000 112.2000 149.2000 ;
	    RECT 111.8000 148.2000 112.1000 148.8000 ;
	    RECT 109.4000 148.1000 109.8000 148.2000 ;
	    RECT 110.2000 148.1000 110.6000 148.2000 ;
	    RECT 109.4000 147.8000 110.6000 148.1000 ;
	    RECT 111.8000 148.1000 112.2000 148.2000 ;
	    RECT 112.6000 148.1000 113.0000 148.2000 ;
	    RECT 111.8000 147.8000 113.0000 148.1000 ;
	    RECT 115.0000 147.2000 115.3000 149.8000 ;
	    RECT 122.2000 148.8000 122.6000 149.2000 ;
	    RECT 122.2000 148.2000 122.5000 148.8000 ;
	    RECT 120.6000 148.1000 121.0000 148.2000 ;
	    RECT 121.4000 148.1000 121.8000 148.2000 ;
	    RECT 120.6000 147.8000 121.8000 148.1000 ;
	    RECT 122.2000 147.8000 122.6000 148.2000 ;
	    RECT 109.4000 147.1000 109.8000 147.2000 ;
	    RECT 110.2000 147.1000 110.6000 147.2000 ;
	    RECT 109.4000 146.8000 110.6000 147.1000 ;
	    RECT 112.6000 146.8000 113.0000 147.2000 ;
	    RECT 115.0000 146.8000 115.4000 147.2000 ;
	    RECT 119.0000 146.8000 119.4000 147.2000 ;
	    RECT 119.8000 147.1000 120.2000 147.2000 ;
	    RECT 120.6000 147.1000 121.0000 147.2000 ;
	    RECT 119.8000 146.8000 121.0000 147.1000 ;
	    RECT 107.0000 146.1000 107.4000 146.2000 ;
	    RECT 107.8000 146.1000 108.2000 146.2000 ;
	    RECT 107.0000 145.8000 108.2000 146.1000 ;
	    RECT 111.8000 145.8000 112.2000 146.2000 ;
	    RECT 103.0000 145.1000 103.4000 145.2000 ;
	    RECT 103.8000 145.1000 104.2000 145.2000 ;
	    RECT 103.0000 144.8000 104.2000 145.1000 ;
	    RECT 106.2000 144.8000 106.6000 145.2000 ;
	    RECT 102.2000 143.8000 102.6000 144.2000 ;
	    RECT 107.8000 137.8000 108.2000 138.2000 ;
	    RECT 99.8000 136.1000 100.2000 136.2000 ;
	    RECT 100.6000 136.1000 101.0000 136.2000 ;
	    RECT 99.8000 135.8000 101.0000 136.1000 ;
	    RECT 102.2000 136.1000 102.6000 136.2000 ;
	    RECT 103.0000 136.1000 103.4000 136.2000 ;
	    RECT 102.2000 135.8000 103.4000 136.1000 ;
	    RECT 106.2000 134.8000 106.6000 135.2000 ;
	    RECT 100.6000 133.8000 101.0000 134.2000 ;
	    RECT 98.2000 133.1000 98.6000 133.2000 ;
	    RECT 99.0000 133.1000 99.4000 133.2000 ;
	    RECT 98.2000 132.8000 99.4000 133.1000 ;
	    RECT 100.6000 132.2000 100.9000 133.8000 ;
	    RECT 103.0000 133.1000 103.4000 133.2000 ;
	    RECT 103.8000 133.1000 104.2000 133.2000 ;
	    RECT 103.0000 132.8000 104.2000 133.1000 ;
	    RECT 100.6000 131.8000 101.0000 132.2000 ;
	    RECT 103.8000 131.8000 104.2000 132.2000 ;
	    RECT 105.4000 131.8000 105.8000 132.2000 ;
	    RECT 99.8000 127.8000 100.2000 128.2000 ;
	    RECT 97.4000 127.1000 97.8000 127.2000 ;
	    RECT 96.6000 126.8000 97.8000 127.1000 ;
	    RECT 98.2000 126.9000 98.6000 127.0000 ;
	    RECT 99.0000 126.9000 99.4000 127.0000 ;
	    RECT 96.6000 125.8000 97.0000 126.2000 ;
	    RECT 96.6000 123.2000 96.9000 125.8000 ;
	    RECT 97.4000 125.2000 97.7000 126.8000 ;
	    RECT 98.2000 126.6000 99.4000 126.9000 ;
	    RECT 99.8000 126.2000 100.1000 127.8000 ;
	    RECT 100.6000 127.2000 100.9000 131.8000 ;
	    RECT 100.6000 126.8000 101.0000 127.2000 ;
	    RECT 102.2000 126.8000 102.6000 127.2000 ;
	    RECT 99.8000 125.8000 100.2000 126.2000 ;
	    RECT 102.2000 125.2000 102.5000 126.8000 ;
	    RECT 103.8000 126.2000 104.1000 131.8000 ;
	    RECT 105.4000 131.2000 105.7000 131.8000 ;
	    RECT 105.4000 130.8000 105.8000 131.2000 ;
	    RECT 106.2000 129.2000 106.5000 134.8000 ;
	    RECT 107.0000 133.8000 107.4000 134.2000 ;
	    RECT 107.0000 133.2000 107.3000 133.8000 ;
	    RECT 107.8000 133.2000 108.1000 137.8000 ;
	    RECT 111.8000 135.2000 112.1000 145.8000 ;
	    RECT 112.6000 145.2000 112.9000 146.8000 ;
	    RECT 115.0000 146.2000 115.3000 146.8000 ;
	    RECT 115.0000 145.8000 115.4000 146.2000 ;
	    RECT 117.4000 145.8000 117.8000 146.2000 ;
	    RECT 118.2000 145.8000 118.6000 146.2000 ;
	    RECT 117.4000 145.2000 117.7000 145.8000 ;
	    RECT 112.6000 144.8000 113.0000 145.2000 ;
	    RECT 117.4000 144.8000 117.8000 145.2000 ;
	    RECT 118.2000 144.2000 118.5000 145.8000 ;
	    RECT 119.0000 144.2000 119.3000 146.8000 ;
	    RECT 116.6000 143.8000 117.0000 144.2000 ;
	    RECT 118.2000 143.8000 118.6000 144.2000 ;
	    RECT 119.0000 143.8000 119.4000 144.2000 ;
	    RECT 113.4000 141.8000 113.8000 142.2000 ;
	    RECT 112.6000 135.8000 113.0000 136.2000 ;
	    RECT 112.6000 135.2000 112.9000 135.8000 ;
	    RECT 110.2000 134.8000 110.6000 135.2000 ;
	    RECT 111.8000 134.8000 112.2000 135.2000 ;
	    RECT 112.6000 134.8000 113.0000 135.2000 ;
	    RECT 107.0000 132.8000 107.4000 133.2000 ;
	    RECT 107.8000 132.8000 108.2000 133.2000 ;
	    RECT 110.2000 129.2000 110.5000 134.8000 ;
	    RECT 111.8000 134.1000 112.1000 134.8000 ;
	    RECT 111.8000 133.8000 112.9000 134.1000 ;
	    RECT 112.6000 133.2000 112.9000 133.8000 ;
	    RECT 111.0000 133.1000 111.4000 133.2000 ;
	    RECT 111.8000 133.1000 112.2000 133.2000 ;
	    RECT 111.0000 132.8000 112.2000 133.1000 ;
	    RECT 112.6000 132.8000 113.0000 133.2000 ;
	    RECT 113.4000 129.2000 113.7000 141.8000 ;
	    RECT 116.6000 135.2000 116.9000 143.8000 ;
	    RECT 118.2000 143.2000 118.5000 143.8000 ;
	    RECT 118.2000 142.8000 118.6000 143.2000 ;
	    RECT 118.2000 141.8000 118.6000 142.2000 ;
	    RECT 118.2000 138.2000 118.5000 141.8000 ;
	    RECT 123.0000 139.2000 123.3000 154.8000 ;
	    RECT 123.8000 153.1000 124.2000 155.9000 ;
	    RECT 125.4000 152.1000 125.8000 157.9000 ;
	    RECT 129.4000 155.2000 129.7000 166.8000 ;
	    RECT 130.2000 165.1000 130.6000 167.9000 ;
	    RECT 131.0000 167.8000 131.4000 168.2000 ;
	    RECT 133.4000 167.8000 133.8000 168.2000 ;
	    RECT 134.2000 168.1000 134.6000 168.2000 ;
	    RECT 135.0000 168.1000 135.4000 168.2000 ;
	    RECT 134.2000 167.8000 135.4000 168.1000 ;
	    RECT 139.8000 167.8000 140.2000 168.2000 ;
	    RECT 132.6000 166.8000 133.0000 167.2000 ;
	    RECT 132.6000 166.2000 132.9000 166.8000 ;
	    RECT 132.6000 165.8000 133.0000 166.2000 ;
	    RECT 132.6000 161.8000 133.0000 162.2000 ;
	    RECT 132.6000 159.2000 132.9000 161.8000 ;
	    RECT 132.6000 158.8000 133.0000 159.2000 ;
	    RECT 127.0000 154.8000 127.4000 155.2000 ;
	    RECT 129.4000 154.8000 129.8000 155.2000 ;
	    RECT 127.0000 151.2000 127.3000 154.8000 ;
	    RECT 129.4000 153.2000 129.7000 154.8000 ;
	    RECT 129.4000 153.1000 129.8000 153.2000 ;
	    RECT 128.6000 152.8000 129.8000 153.1000 ;
	    RECT 127.0000 150.8000 127.4000 151.2000 ;
	    RECT 124.6000 143.1000 125.0000 148.9000 ;
	    RECT 128.6000 148.2000 128.9000 152.8000 ;
	    RECT 130.2000 152.1000 130.6000 157.9000 ;
	    RECT 133.4000 155.2000 133.7000 167.8000 ;
	    RECT 136.6000 166.8000 137.0000 167.2000 ;
	    RECT 141.4000 166.8000 141.8000 167.2000 ;
	    RECT 134.2000 165.8000 134.6000 166.2000 ;
	    RECT 134.2000 163.2000 134.5000 165.8000 ;
	    RECT 136.6000 164.2000 136.9000 166.8000 ;
	    RECT 141.4000 166.2000 141.7000 166.8000 ;
	    RECT 139.8000 165.8000 140.2000 166.2000 ;
	    RECT 141.4000 165.8000 141.8000 166.2000 ;
	    RECT 136.6000 163.8000 137.0000 164.2000 ;
	    RECT 138.2000 163.8000 138.6000 164.2000 ;
	    RECT 134.2000 162.8000 134.6000 163.2000 ;
	    RECT 135.8000 156.8000 136.2000 157.2000 ;
	    RECT 135.8000 156.2000 136.1000 156.8000 ;
	    RECT 135.8000 155.8000 136.2000 156.2000 ;
	    RECT 133.4000 154.8000 133.8000 155.2000 ;
	    RECT 135.8000 154.8000 136.2000 155.2000 ;
	    RECT 136.6000 154.8000 137.0000 155.2000 ;
	    RECT 137.4000 154.8000 137.8000 155.2000 ;
	    RECT 133.4000 153.2000 133.7000 154.8000 ;
	    RECT 134.2000 154.1000 134.6000 154.2000 ;
	    RECT 135.0000 154.1000 135.4000 154.2000 ;
	    RECT 134.2000 153.8000 135.4000 154.1000 ;
	    RECT 133.4000 152.8000 133.8000 153.2000 ;
	    RECT 132.6000 152.1000 133.0000 152.2000 ;
	    RECT 133.4000 152.1000 133.8000 152.2000 ;
	    RECT 132.6000 151.8000 133.8000 152.1000 ;
	    RECT 128.6000 147.8000 129.0000 148.2000 ;
	    RECT 127.8000 145.8000 128.2000 146.2000 ;
	    RECT 127.8000 145.2000 128.1000 145.8000 ;
	    RECT 127.8000 144.8000 128.2000 145.2000 ;
	    RECT 128.6000 142.8000 129.0000 143.2000 ;
	    RECT 129.4000 143.1000 129.8000 148.9000 ;
	    RECT 135.8000 148.2000 136.1000 154.8000 ;
	    RECT 136.6000 153.2000 136.9000 154.8000 ;
	    RECT 137.4000 154.2000 137.7000 154.8000 ;
	    RECT 138.2000 154.2000 138.5000 163.8000 ;
	    RECT 139.8000 163.2000 140.1000 165.8000 ;
	    RECT 139.8000 162.8000 140.2000 163.2000 ;
	    RECT 142.2000 162.2000 142.5000 174.8000 ;
	    RECT 144.6000 167.2000 144.9000 174.8000 ;
	    RECT 147.0000 172.2000 147.3000 174.8000 ;
	    RECT 147.0000 171.8000 147.4000 172.2000 ;
	    RECT 144.6000 166.8000 145.0000 167.2000 ;
	    RECT 146.2000 163.1000 146.6000 168.9000 ;
	    RECT 147.0000 165.8000 147.4000 166.2000 ;
	    RECT 147.8000 166.1000 148.2000 166.2000 ;
	    RECT 148.6000 166.1000 149.0000 166.2000 ;
	    RECT 147.8000 165.8000 149.0000 166.1000 ;
	    RECT 142.2000 161.8000 142.6000 162.2000 ;
	    RECT 140.6000 155.8000 141.0000 156.2000 ;
	    RECT 137.4000 153.8000 137.8000 154.2000 ;
	    RECT 138.2000 153.8000 138.6000 154.2000 ;
	    RECT 136.6000 152.8000 137.0000 153.2000 ;
	    RECT 136.6000 151.8000 137.0000 152.2000 ;
	    RECT 136.6000 148.2000 136.9000 151.8000 ;
	    RECT 131.0000 145.1000 131.4000 147.9000 ;
	    RECT 135.8000 147.8000 136.2000 148.2000 ;
	    RECT 136.6000 147.8000 137.0000 148.2000 ;
	    RECT 138.2000 147.2000 138.5000 153.8000 ;
	    RECT 140.6000 153.2000 140.9000 155.8000 ;
	    RECT 140.6000 152.8000 141.0000 153.2000 ;
	    RECT 141.4000 153.1000 141.8000 155.9000 ;
	    RECT 142.2000 153.8000 142.6000 154.2000 ;
	    RECT 139.8000 150.8000 140.2000 151.2000 ;
	    RECT 139.8000 149.2000 140.1000 150.8000 ;
	    RECT 139.8000 148.8000 140.2000 149.2000 ;
	    RECT 131.8000 146.8000 132.2000 147.2000 ;
	    RECT 134.2000 147.1000 134.6000 147.2000 ;
	    RECT 135.0000 147.1000 135.4000 147.2000 ;
	    RECT 134.2000 146.8000 135.4000 147.1000 ;
	    RECT 138.2000 146.8000 138.6000 147.2000 ;
	    RECT 140.6000 146.8000 141.0000 147.2000 ;
	    RECT 128.6000 139.2000 128.9000 142.8000 ;
	    RECT 131.8000 139.2000 132.1000 146.8000 ;
	    RECT 140.6000 146.2000 140.9000 146.8000 ;
	    RECT 142.2000 146.2000 142.5000 153.8000 ;
	    RECT 143.0000 152.1000 143.4000 157.9000 ;
	    RECT 147.0000 155.2000 147.3000 165.8000 ;
	    RECT 143.8000 155.0000 144.2000 155.1000 ;
	    RECT 144.6000 155.0000 145.0000 155.1000 ;
	    RECT 143.8000 154.7000 145.0000 155.0000 ;
	    RECT 147.0000 154.8000 147.4000 155.2000 ;
	    RECT 147.0000 153.2000 147.3000 154.8000 ;
	    RECT 147.0000 152.8000 147.4000 153.2000 ;
	    RECT 147.8000 152.1000 148.2000 157.9000 ;
	    RECT 149.4000 148.2000 149.7000 174.8000 ;
	    RECT 153.4000 169.2000 153.7000 174.8000 ;
	    RECT 156.6000 172.1000 157.0000 177.9000 ;
	    RECT 160.6000 174.7000 161.0000 175.1000 ;
	    RECT 160.6000 174.2000 160.9000 174.7000 ;
	    RECT 160.6000 173.8000 161.0000 174.2000 ;
	    RECT 161.4000 172.1000 161.8000 177.9000 ;
	    RECT 163.0000 173.1000 163.4000 175.9000 ;
	    RECT 165.4000 174.8000 165.8000 175.2000 ;
	    RECT 166.2000 175.1000 166.6000 175.2000 ;
	    RECT 167.0000 175.1000 167.4000 175.2000 ;
	    RECT 166.2000 174.8000 167.4000 175.1000 ;
	    RECT 171.0000 174.8000 171.4000 175.2000 ;
	    RECT 171.8000 174.8000 172.2000 175.2000 ;
	    RECT 164.6000 173.8000 165.0000 174.2000 ;
	    RECT 164.6000 173.2000 164.9000 173.8000 ;
	    RECT 165.4000 173.2000 165.7000 174.8000 ;
	    RECT 167.0000 173.8000 167.4000 174.2000 ;
	    RECT 164.6000 172.8000 165.0000 173.2000 ;
	    RECT 165.4000 172.8000 165.8000 173.2000 ;
	    RECT 151.0000 163.1000 151.4000 168.9000 ;
	    RECT 153.4000 168.8000 153.8000 169.2000 ;
	    RECT 154.2000 169.1000 154.6000 169.2000 ;
	    RECT 155.0000 169.1000 155.4000 169.2000 ;
	    RECT 154.2000 168.8000 155.4000 169.1000 ;
	    RECT 153.4000 168.2000 153.7000 168.8000 ;
	    RECT 151.8000 165.8000 152.2000 166.2000 ;
	    RECT 151.8000 159.2000 152.1000 165.8000 ;
	    RECT 152.6000 165.1000 153.0000 167.9000 ;
	    RECT 153.4000 167.8000 153.8000 168.2000 ;
	    RECT 153.4000 166.8000 153.8000 167.2000 ;
	    RECT 153.4000 166.2000 153.7000 166.8000 ;
	    RECT 153.4000 165.8000 153.8000 166.2000 ;
	    RECT 157.4000 163.1000 157.8000 168.9000 ;
	    RECT 158.2000 166.8000 158.6000 167.2000 ;
	    RECT 158.2000 166.2000 158.5000 166.8000 ;
	    RECT 158.2000 165.8000 158.6000 166.2000 ;
	    RECT 159.8000 166.1000 160.2000 166.2000 ;
	    RECT 160.6000 166.1000 161.0000 166.2000 ;
	    RECT 159.8000 165.8000 161.0000 166.1000 ;
	    RECT 158.2000 164.8000 158.6000 165.2000 ;
	    RECT 154.2000 161.8000 154.6000 162.2000 ;
	    RECT 151.8000 158.8000 152.2000 159.2000 ;
	    RECT 150.2000 156.8000 150.6000 157.2000 ;
	    RECT 151.0000 156.8000 151.4000 157.2000 ;
	    RECT 150.2000 156.2000 150.5000 156.8000 ;
	    RECT 150.2000 155.8000 150.6000 156.2000 ;
	    RECT 151.0000 155.2000 151.3000 156.8000 ;
	    RECT 154.2000 155.2000 154.5000 161.8000 ;
	    RECT 155.0000 155.8000 155.4000 156.2000 ;
	    RECT 155.0000 155.2000 155.3000 155.8000 ;
	    RECT 151.0000 154.8000 151.4000 155.2000 ;
	    RECT 154.2000 154.8000 154.6000 155.2000 ;
	    RECT 155.0000 154.8000 155.4000 155.2000 ;
	    RECT 158.2000 154.2000 158.5000 164.8000 ;
	    RECT 162.2000 163.1000 162.6000 168.9000 ;
	    RECT 163.8000 165.1000 164.2000 167.9000 ;
	    RECT 159.0000 157.1000 159.4000 157.2000 ;
	    RECT 159.8000 157.1000 160.2000 157.2000 ;
	    RECT 159.0000 156.8000 160.2000 157.1000 ;
	    RECT 151.8000 154.1000 152.2000 154.2000 ;
	    RECT 152.6000 154.1000 153.0000 154.2000 ;
	    RECT 151.8000 153.8000 153.0000 154.1000 ;
	    RECT 153.4000 153.8000 153.8000 154.2000 ;
	    RECT 158.2000 153.8000 158.6000 154.2000 ;
	    RECT 151.8000 152.8000 152.2000 153.2000 ;
	    RECT 149.4000 147.8000 149.8000 148.2000 ;
	    RECT 143.0000 146.8000 143.4000 147.2000 ;
	    RECT 143.8000 147.1000 144.2000 147.2000 ;
	    RECT 144.6000 147.1000 145.0000 147.2000 ;
	    RECT 143.8000 146.8000 145.0000 147.1000 ;
	    RECT 143.0000 146.2000 143.3000 146.8000 ;
	    RECT 140.6000 145.8000 141.0000 146.2000 ;
	    RECT 142.2000 145.8000 142.6000 146.2000 ;
	    RECT 143.0000 145.8000 143.4000 146.2000 ;
	    RECT 143.8000 146.1000 144.2000 146.2000 ;
	    RECT 144.6000 146.1000 145.0000 146.2000 ;
	    RECT 143.8000 145.8000 145.0000 146.1000 ;
	    RECT 150.2000 143.1000 150.6000 148.9000 ;
	    RECT 151.8000 146.2000 152.1000 152.8000 ;
	    RECT 153.4000 147.2000 153.7000 153.8000 ;
	    RECT 158.2000 149.2000 158.5000 153.8000 ;
	    RECT 161.4000 152.1000 161.8000 157.9000 ;
	    RECT 164.6000 154.2000 164.9000 172.8000 ;
	    RECT 166.2000 171.8000 166.6000 172.2000 ;
	    RECT 166.2000 168.2000 166.5000 171.8000 ;
	    RECT 167.0000 169.2000 167.3000 173.8000 ;
	    RECT 171.0000 173.1000 171.3000 174.8000 ;
	    RECT 171.8000 174.2000 172.1000 174.8000 ;
	    RECT 171.8000 173.8000 172.2000 174.2000 ;
	    RECT 174.2000 173.1000 174.6000 175.9000 ;
	    RECT 175.0000 173.8000 175.4000 174.2000 ;
	    RECT 175.0000 173.2000 175.3000 173.8000 ;
	    RECT 171.0000 172.8000 172.1000 173.1000 ;
	    RECT 175.0000 172.8000 175.4000 173.2000 ;
	    RECT 171.8000 169.2000 172.1000 172.8000 ;
	    RECT 175.8000 172.1000 176.2000 177.9000 ;
	    RECT 177.4000 174.8000 177.8000 175.2000 ;
	    RECT 177.4000 173.2000 177.7000 174.8000 ;
	    RECT 177.4000 172.8000 177.8000 173.2000 ;
	    RECT 180.6000 172.1000 181.0000 177.9000 ;
	    RECT 183.0000 177.1000 183.4000 177.2000 ;
	    RECT 183.8000 177.1000 184.2000 177.2000 ;
	    RECT 183.0000 176.8000 184.2000 177.1000 ;
	    RECT 187.0000 176.8000 187.4000 177.2000 ;
	    RECT 187.0000 175.2000 187.3000 176.8000 ;
	    RECT 183.8000 175.1000 184.2000 175.2000 ;
	    RECT 183.0000 174.8000 184.2000 175.1000 ;
	    RECT 187.0000 174.8000 187.4000 175.2000 ;
	    RECT 167.0000 168.8000 167.4000 169.2000 ;
	    RECT 171.8000 168.8000 172.2000 169.2000 ;
	    RECT 180.6000 169.1000 181.0000 169.2000 ;
	    RECT 181.4000 169.1000 181.8000 169.2000 ;
	    RECT 171.8000 168.2000 172.1000 168.8000 ;
	    RECT 166.2000 167.8000 166.6000 168.2000 ;
	    RECT 171.8000 167.8000 172.2000 168.2000 ;
	    RECT 170.2000 166.8000 170.6000 167.2000 ;
	    RECT 170.2000 166.2000 170.5000 166.8000 ;
	    RECT 167.8000 165.8000 168.2000 166.2000 ;
	    RECT 170.2000 165.8000 170.6000 166.2000 ;
	    RECT 167.8000 165.2000 168.1000 165.8000 ;
	    RECT 167.8000 164.8000 168.2000 165.2000 ;
	    RECT 172.6000 165.1000 173.0000 167.9000 ;
	    RECT 173.4000 167.8000 173.8000 168.2000 ;
	    RECT 173.4000 167.2000 173.7000 167.8000 ;
	    RECT 173.4000 166.8000 173.8000 167.2000 ;
	    RECT 174.2000 163.1000 174.6000 168.9000 ;
	    RECT 175.0000 166.8000 175.4000 167.2000 ;
	    RECT 175.0000 166.3000 175.3000 166.8000 ;
	    RECT 175.0000 165.9000 175.4000 166.3000 ;
	    RECT 179.0000 163.1000 179.4000 168.9000 ;
	    RECT 180.6000 168.8000 181.8000 169.1000 ;
	    RECT 182.2000 165.8000 182.6000 166.2000 ;
	    RECT 182.2000 165.2000 182.5000 165.8000 ;
	    RECT 182.2000 164.8000 182.6000 165.2000 ;
	    RECT 165.4000 155.8000 165.8000 156.2000 ;
	    RECT 165.4000 155.1000 165.7000 155.8000 ;
	    RECT 165.4000 154.7000 165.8000 155.1000 ;
	    RECT 164.6000 153.8000 165.0000 154.2000 ;
	    RECT 166.2000 152.1000 166.6000 157.9000 ;
	    RECT 171.8000 156.8000 172.2000 157.2000 ;
	    RECT 171.8000 156.2000 172.1000 156.8000 ;
	    RECT 171.8000 156.1000 172.2000 156.2000 ;
	    RECT 172.6000 156.1000 173.0000 156.2000 ;
	    RECT 167.0000 153.8000 167.4000 154.2000 ;
	    RECT 153.4000 146.8000 153.8000 147.2000 ;
	    RECT 151.8000 145.8000 152.2000 146.2000 ;
	    RECT 152.6000 146.1000 153.0000 146.2000 ;
	    RECT 153.4000 146.1000 153.8000 146.2000 ;
	    RECT 152.6000 145.8000 153.8000 146.1000 ;
	    RECT 132.6000 141.8000 133.0000 142.2000 ;
	    RECT 135.8000 141.8000 136.2000 142.2000 ;
	    RECT 123.0000 138.8000 123.4000 139.2000 ;
	    RECT 128.6000 138.8000 129.0000 139.2000 ;
	    RECT 131.8000 138.8000 132.2000 139.2000 ;
	    RECT 118.2000 137.8000 118.6000 138.2000 ;
	    RECT 116.6000 134.8000 117.0000 135.2000 ;
	    RECT 114.2000 134.0000 114.6000 134.4000 ;
	    RECT 114.2000 132.2000 114.5000 134.0000 ;
	    RECT 118.2000 133.8000 118.6000 134.2000 ;
	    RECT 118.2000 133.2000 118.5000 133.8000 ;
	    RECT 118.2000 132.8000 118.6000 133.2000 ;
	    RECT 119.8000 132.8000 120.2000 133.2000 ;
	    RECT 114.2000 131.8000 114.6000 132.2000 ;
	    RECT 115.8000 131.8000 116.2000 132.2000 ;
	    RECT 117.4000 131.8000 117.8000 132.2000 ;
	    RECT 118.2000 132.1000 118.6000 132.2000 ;
	    RECT 119.0000 132.1000 119.4000 132.2000 ;
	    RECT 118.2000 131.8000 119.4000 132.1000 ;
	    RECT 106.2000 128.8000 106.6000 129.2000 ;
	    RECT 110.2000 128.8000 110.6000 129.2000 ;
	    RECT 111.0000 129.1000 111.4000 129.2000 ;
	    RECT 111.8000 129.1000 112.2000 129.2000 ;
	    RECT 111.0000 128.8000 112.2000 129.1000 ;
	    RECT 113.4000 128.8000 113.8000 129.2000 ;
	    RECT 115.8000 128.2000 116.1000 131.8000 ;
	    RECT 105.4000 128.1000 105.8000 128.2000 ;
	    RECT 106.2000 128.1000 106.6000 128.2000 ;
	    RECT 105.4000 127.8000 106.6000 128.1000 ;
	    RECT 114.2000 127.8000 114.6000 128.2000 ;
	    RECT 115.8000 127.8000 116.2000 128.2000 ;
	    RECT 103.8000 125.8000 104.2000 126.2000 ;
	    RECT 97.4000 124.8000 97.8000 125.2000 ;
	    RECT 101.4000 125.1000 101.8000 125.2000 ;
	    RECT 102.2000 125.1000 102.6000 125.2000 ;
	    RECT 101.4000 124.8000 102.6000 125.1000 ;
	    RECT 105.4000 124.8000 105.8000 125.2000 ;
	    RECT 96.6000 122.8000 97.0000 123.2000 ;
	    RECT 84.6000 121.8000 85.0000 122.2000 ;
	    RECT 90.2000 121.8000 90.6000 122.2000 ;
	    RECT 91.8000 121.8000 92.2000 122.2000 ;
	    RECT 101.4000 121.8000 101.8000 122.2000 ;
	    RECT 84.6000 112.1000 85.0000 117.9000 ;
	    RECT 90.2000 116.2000 90.5000 121.8000 ;
	    RECT 101.4000 118.2000 101.7000 121.8000 ;
	    RECT 105.4000 121.2000 105.7000 124.8000 ;
	    RECT 105.4000 120.8000 105.8000 121.2000 ;
	    RECT 85.4000 115.8000 85.8000 116.2000 ;
	    RECT 85.4000 114.2000 85.7000 115.8000 ;
	    RECT 85.4000 113.8000 85.8000 114.2000 ;
	    RECT 86.2000 113.1000 86.6000 115.9000 ;
	    RECT 87.0000 114.8000 87.4000 115.2000 ;
	    RECT 88.6000 114.8000 89.0000 115.2000 ;
	    RECT 87.0000 113.2000 87.3000 114.8000 ;
	    RECT 88.6000 114.2000 88.9000 114.8000 ;
	    RECT 88.6000 113.8000 89.0000 114.2000 ;
	    RECT 87.0000 112.8000 87.4000 113.2000 ;
	    RECT 87.8000 113.1000 88.2000 113.2000 ;
	    RECT 88.6000 113.1000 89.0000 113.2000 ;
	    RECT 89.4000 113.1000 89.8000 115.9000 ;
	    RECT 90.2000 115.8000 90.6000 116.2000 ;
	    RECT 90.2000 114.2000 90.5000 115.8000 ;
	    RECT 90.2000 113.8000 90.6000 114.2000 ;
	    RECT 87.8000 112.8000 89.0000 113.1000 ;
	    RECT 90.2000 111.8000 90.6000 112.2000 ;
	    RECT 91.0000 112.1000 91.4000 117.9000 ;
	    RECT 91.8000 115.0000 92.2000 115.1000 ;
	    RECT 92.6000 115.0000 93.0000 115.1000 ;
	    RECT 91.8000 114.7000 93.0000 115.0000 ;
	    RECT 93.4000 113.8000 93.8000 114.2000 ;
	    RECT 90.2000 111.2000 90.5000 111.8000 ;
	    RECT 83.0000 109.8000 84.1000 110.1000 ;
	    RECT 84.6000 110.8000 85.0000 111.2000 ;
	    RECT 90.2000 110.8000 90.6000 111.2000 ;
	    RECT 83.0000 107.2000 83.3000 109.8000 ;
	    RECT 84.6000 109.2000 84.9000 110.8000 ;
	    RECT 87.0000 109.8000 87.4000 110.2000 ;
	    RECT 87.0000 109.2000 87.3000 109.8000 ;
	    RECT 84.6000 108.8000 85.0000 109.2000 ;
	    RECT 87.0000 108.8000 87.4000 109.2000 ;
	    RECT 83.8000 107.8000 84.2000 108.2000 ;
	    RECT 83.0000 106.8000 83.4000 107.2000 ;
	    RECT 77.4000 105.8000 77.8000 106.2000 ;
	    RECT 79.8000 105.8000 80.2000 106.2000 ;
	    RECT 82.2000 105.8000 82.6000 106.2000 ;
	    RECT 79.8000 99.2000 80.1000 105.8000 ;
	    RECT 82.2000 105.2000 82.5000 105.8000 ;
	    RECT 80.6000 104.8000 81.0000 105.2000 ;
	    RECT 82.2000 104.8000 82.6000 105.2000 ;
	    RECT 80.6000 104.2000 80.9000 104.8000 ;
	    RECT 80.6000 103.8000 81.0000 104.2000 ;
	    RECT 83.8000 101.2000 84.1000 107.8000 ;
	    RECT 86.2000 105.8000 86.6000 106.2000 ;
	    RECT 86.2000 104.2000 86.5000 105.8000 ;
	    RECT 87.0000 105.2000 87.3000 108.8000 ;
	    RECT 90.2000 107.2000 90.5000 110.8000 ;
	    RECT 93.4000 108.2000 93.7000 113.8000 ;
	    RECT 95.8000 112.1000 96.2000 117.9000 ;
	    RECT 101.4000 117.8000 101.8000 118.2000 ;
	    RECT 106.2000 117.2000 106.5000 127.8000 ;
	    RECT 112.6000 127.1000 113.0000 127.2000 ;
	    RECT 113.4000 127.1000 113.8000 127.2000 ;
	    RECT 112.6000 126.8000 113.8000 127.1000 ;
	    RECT 114.2000 126.2000 114.5000 127.8000 ;
	    RECT 111.0000 125.8000 111.4000 126.2000 ;
	    RECT 114.2000 125.8000 114.6000 126.2000 ;
	    RECT 111.0000 125.2000 111.3000 125.8000 ;
	    RECT 117.4000 125.2000 117.7000 131.8000 ;
	    RECT 119.8000 129.2000 120.1000 132.8000 ;
	    RECT 121.4000 132.1000 121.8000 137.9000 ;
	    RECT 119.8000 128.8000 120.2000 129.2000 ;
	    RECT 123.0000 128.2000 123.3000 138.8000 ;
	    RECT 123.8000 135.1000 124.2000 135.2000 ;
	    RECT 124.6000 135.1000 125.0000 135.2000 ;
	    RECT 123.8000 134.8000 125.0000 135.1000 ;
	    RECT 126.2000 132.1000 126.6000 137.9000 ;
	    RECT 127.0000 133.8000 127.4000 134.2000 ;
	    RECT 124.6000 128.8000 125.0000 129.2000 ;
	    RECT 123.0000 127.8000 123.4000 128.2000 ;
	    RECT 119.0000 127.1000 119.4000 127.2000 ;
	    RECT 119.8000 127.1000 120.2000 127.2000 ;
	    RECT 119.0000 126.8000 120.2000 127.1000 ;
	    RECT 124.6000 126.2000 124.9000 128.8000 ;
	    RECT 127.0000 127.2000 127.3000 133.8000 ;
	    RECT 127.8000 133.1000 128.2000 135.9000 ;
	    RECT 127.8000 131.8000 128.2000 132.2000 ;
	    RECT 128.6000 131.8000 129.0000 132.2000 ;
	    RECT 131.0000 132.1000 131.4000 137.9000 ;
	    RECT 127.8000 129.2000 128.1000 131.8000 ;
	    RECT 128.6000 129.2000 128.9000 131.8000 ;
	    RECT 127.8000 128.8000 128.2000 129.2000 ;
	    RECT 128.6000 128.8000 129.0000 129.2000 ;
	    RECT 127.0000 126.8000 127.4000 127.2000 ;
	    RECT 118.2000 126.1000 118.6000 126.2000 ;
	    RECT 119.0000 126.1000 119.4000 126.2000 ;
	    RECT 118.2000 125.8000 119.4000 126.1000 ;
	    RECT 124.6000 125.8000 125.0000 126.2000 ;
	    RECT 125.4000 125.8000 125.8000 126.2000 ;
	    RECT 111.0000 124.8000 111.4000 125.2000 ;
	    RECT 113.4000 125.1000 113.8000 125.2000 ;
	    RECT 114.2000 125.1000 114.6000 125.2000 ;
	    RECT 113.4000 124.8000 114.6000 125.1000 ;
	    RECT 117.4000 124.8000 117.8000 125.2000 ;
	    RECT 115.0000 124.1000 115.4000 124.2000 ;
	    RECT 115.8000 124.1000 116.2000 124.2000 ;
	    RECT 115.0000 123.8000 116.2000 124.1000 ;
	    RECT 116.6000 123.8000 117.0000 124.2000 ;
	    RECT 116.6000 123.2000 116.9000 123.8000 ;
	    RECT 113.4000 123.1000 113.8000 123.2000 ;
	    RECT 114.2000 123.1000 114.6000 123.2000 ;
	    RECT 113.4000 122.8000 114.6000 123.1000 ;
	    RECT 116.6000 122.8000 117.0000 123.2000 ;
	    RECT 121.4000 121.8000 121.8000 122.2000 ;
	    RECT 121.4000 120.2000 121.7000 121.8000 ;
	    RECT 121.4000 119.8000 121.8000 120.2000 ;
	    RECT 125.4000 119.2000 125.7000 125.8000 ;
	    RECT 126.2000 124.8000 126.6000 125.2000 ;
	    RECT 126.2000 124.2000 126.5000 124.8000 ;
	    RECT 126.2000 123.8000 126.6000 124.2000 ;
	    RECT 125.4000 118.8000 125.8000 119.2000 ;
	    RECT 106.2000 116.8000 106.6000 117.2000 ;
	    RECT 106.2000 115.8000 106.6000 116.2000 ;
	    RECT 108.6000 116.1000 109.0000 116.2000 ;
	    RECT 109.4000 116.1000 109.8000 116.2000 ;
	    RECT 108.6000 115.8000 109.8000 116.1000 ;
	    RECT 106.2000 115.2000 106.5000 115.8000 ;
	    RECT 99.8000 114.8000 100.2000 115.2000 ;
	    RECT 102.2000 114.8000 102.6000 115.2000 ;
	    RECT 106.2000 114.8000 106.6000 115.2000 ;
	    RECT 112.6000 114.8000 113.0000 115.2000 ;
	    RECT 117.4000 114.8000 117.8000 115.2000 ;
	    RECT 125.4000 114.8000 125.8000 115.2000 ;
	    RECT 99.8000 113.2000 100.1000 114.8000 ;
	    RECT 102.2000 114.2000 102.5000 114.8000 ;
	    RECT 102.2000 113.8000 102.6000 114.2000 ;
	    RECT 104.6000 114.1000 105.0000 114.2000 ;
	    RECT 105.4000 114.1000 105.8000 114.2000 ;
	    RECT 104.6000 113.8000 105.8000 114.1000 ;
	    RECT 107.8000 113.8000 108.2000 114.2000 ;
	    RECT 107.8000 113.2000 108.1000 113.8000 ;
	    RECT 112.6000 113.2000 112.9000 114.8000 ;
	    RECT 117.4000 114.2000 117.7000 114.8000 ;
	    RECT 113.4000 113.8000 113.8000 114.2000 ;
	    RECT 116.6000 113.8000 117.0000 114.2000 ;
	    RECT 117.4000 113.8000 117.8000 114.2000 ;
	    RECT 113.4000 113.2000 113.7000 113.8000 ;
	    RECT 116.6000 113.2000 116.9000 113.8000 ;
	    RECT 98.2000 113.1000 98.6000 113.2000 ;
	    RECT 99.0000 113.1000 99.4000 113.2000 ;
	    RECT 98.2000 112.8000 99.4000 113.1000 ;
	    RECT 99.8000 112.8000 100.2000 113.2000 ;
	    RECT 100.6000 112.8000 101.0000 113.2000 ;
	    RECT 107.8000 112.8000 108.2000 113.2000 ;
	    RECT 110.2000 113.1000 110.6000 113.2000 ;
	    RECT 111.0000 113.1000 111.4000 113.2000 ;
	    RECT 110.2000 112.8000 111.4000 113.1000 ;
	    RECT 112.6000 112.8000 113.0000 113.2000 ;
	    RECT 113.4000 112.8000 113.8000 113.2000 ;
	    RECT 116.6000 112.8000 117.0000 113.2000 ;
	    RECT 120.6000 112.8000 121.0000 113.2000 ;
	    RECT 123.8000 113.1000 124.2000 113.2000 ;
	    RECT 124.6000 113.1000 125.0000 113.2000 ;
	    RECT 123.8000 112.8000 125.0000 113.1000 ;
	    RECT 99.8000 112.2000 100.1000 112.8000 ;
	    RECT 98.2000 112.1000 98.6000 112.2000 ;
	    RECT 99.0000 112.1000 99.4000 112.2000 ;
	    RECT 98.2000 111.8000 99.4000 112.1000 ;
	    RECT 99.8000 111.8000 100.2000 112.2000 ;
	    RECT 100.6000 111.2000 100.9000 112.8000 ;
	    RECT 103.0000 111.8000 103.4000 112.2000 ;
	    RECT 107.0000 111.8000 107.4000 112.2000 ;
	    RECT 111.8000 111.8000 112.2000 112.2000 ;
	    RECT 100.6000 110.8000 101.0000 111.2000 ;
	    RECT 101.4000 109.8000 101.8000 110.2000 ;
	    RECT 93.4000 107.8000 93.8000 108.2000 ;
	    RECT 95.0000 107.8000 95.4000 108.2000 ;
	    RECT 95.8000 107.8000 96.2000 108.2000 ;
	    RECT 99.0000 107.8000 99.4000 108.2000 ;
	    RECT 99.8000 108.1000 100.2000 108.2000 ;
	    RECT 100.6000 108.1000 101.0000 108.2000 ;
	    RECT 99.8000 107.8000 101.0000 108.1000 ;
	    RECT 88.6000 107.1000 89.0000 107.2000 ;
	    RECT 89.4000 107.1000 89.8000 107.2000 ;
	    RECT 88.6000 106.8000 89.8000 107.1000 ;
	    RECT 90.2000 106.8000 90.6000 107.2000 ;
	    RECT 89.4000 105.8000 89.8000 106.2000 ;
	    RECT 89.4000 105.2000 89.7000 105.8000 ;
	    RECT 87.0000 104.8000 87.4000 105.2000 ;
	    RECT 89.4000 104.8000 89.8000 105.2000 ;
	    RECT 90.2000 105.1000 90.6000 105.2000 ;
	    RECT 91.0000 105.1000 91.4000 105.2000 ;
	    RECT 90.2000 104.8000 91.4000 105.1000 ;
	    RECT 84.6000 103.8000 85.0000 104.2000 ;
	    RECT 86.2000 103.8000 86.6000 104.2000 ;
	    RECT 83.8000 100.8000 84.2000 101.2000 ;
	    RECT 84.6000 99.2000 84.9000 103.8000 ;
	    RECT 75.0000 98.8000 75.4000 99.2000 ;
	    RECT 79.8000 98.8000 80.2000 99.2000 ;
	    RECT 84.6000 98.8000 85.0000 99.2000 ;
	    RECT 73.4000 97.1000 73.8000 97.2000 ;
	    RECT 74.2000 97.1000 74.6000 97.2000 ;
	    RECT 73.4000 96.8000 74.6000 97.1000 ;
	    RECT 72.6000 95.8000 73.0000 96.2000 ;
	    RECT 72.6000 94.8000 73.0000 95.2000 ;
	    RECT 71.0000 87.8000 71.4000 88.2000 ;
	    RECT 72.6000 84.2000 72.9000 94.8000 ;
	    RECT 75.0000 93.2000 75.3000 98.8000 ;
	    RECT 77.4000 97.8000 77.8000 98.2000 ;
	    RECT 77.4000 96.2000 77.7000 97.8000 ;
	    RECT 80.6000 97.1000 81.0000 97.2000 ;
	    RECT 81.4000 97.1000 81.8000 97.2000 ;
	    RECT 80.6000 96.8000 81.8000 97.1000 ;
	    RECT 83.8000 97.1000 84.2000 97.2000 ;
	    RECT 84.6000 97.1000 85.0000 97.2000 ;
	    RECT 83.8000 96.8000 85.0000 97.1000 ;
	    RECT 87.0000 96.8000 87.4000 97.2000 ;
	    RECT 87.0000 96.2000 87.3000 96.8000 ;
	    RECT 77.4000 95.8000 77.8000 96.2000 ;
	    RECT 87.0000 95.8000 87.4000 96.2000 ;
	    RECT 81.4000 94.8000 81.8000 95.2000 ;
	    RECT 82.2000 94.8000 82.6000 95.2000 ;
	    RECT 84.6000 94.8000 85.0000 95.2000 ;
	    RECT 86.2000 94.8000 86.6000 95.2000 ;
	    RECT 88.6000 94.8000 89.0000 95.2000 ;
	    RECT 79.0000 93.8000 79.4000 94.2000 ;
	    RECT 75.0000 92.8000 75.4000 93.2000 ;
	    RECT 75.8000 91.8000 76.2000 92.2000 ;
	    RECT 79.0000 92.1000 79.3000 93.8000 ;
	    RECT 81.4000 93.2000 81.7000 94.8000 ;
	    RECT 81.4000 92.8000 81.8000 93.2000 ;
	    RECT 79.0000 91.8000 80.1000 92.1000 ;
	    RECT 75.8000 89.2000 76.1000 91.8000 ;
	    RECT 76.6000 89.8000 77.0000 90.2000 ;
	    RECT 73.4000 86.8000 73.8000 87.2000 ;
	    RECT 73.4000 86.3000 73.7000 86.8000 ;
	    RECT 73.4000 85.9000 73.8000 86.3000 ;
	    RECT 72.6000 83.8000 73.0000 84.2000 ;
	    RECT 74.2000 83.1000 74.6000 88.9000 ;
	    RECT 75.8000 88.8000 76.2000 89.2000 ;
	    RECT 76.6000 88.2000 76.9000 89.8000 ;
	    RECT 75.0000 87.8000 75.4000 88.2000 ;
	    RECT 75.0000 87.2000 75.3000 87.8000 ;
	    RECT 75.0000 86.8000 75.4000 87.2000 ;
	    RECT 75.0000 84.8000 75.4000 85.2000 ;
	    RECT 75.8000 85.1000 76.2000 87.9000 ;
	    RECT 76.6000 87.8000 77.0000 88.2000 ;
	    RECT 76.6000 86.8000 77.0000 87.2000 ;
	    RECT 76.6000 86.2000 76.9000 86.8000 ;
	    RECT 76.6000 85.8000 77.0000 86.2000 ;
	    RECT 78.2000 86.1000 78.6000 86.2000 ;
	    RECT 77.4000 85.8000 78.6000 86.1000 ;
	    RECT 65.4000 81.8000 65.8000 82.2000 ;
	    RECT 74.2000 81.8000 74.6000 82.2000 ;
	    RECT 65.4000 76.2000 65.7000 81.8000 ;
	    RECT 65.4000 75.8000 65.8000 76.2000 ;
	    RECT 65.4000 75.0000 65.8000 75.1000 ;
	    RECT 66.2000 75.0000 66.6000 75.1000 ;
	    RECT 65.4000 74.7000 66.6000 75.0000 ;
	    RECT 64.6000 73.8000 65.7000 74.1000 ;
	    RECT 62.2000 70.8000 62.6000 71.2000 ;
	    RECT 56.6000 69.8000 57.0000 70.2000 ;
	    RECT 53.4000 65.8000 53.8000 66.2000 ;
	    RECT 55.8000 65.8000 56.2000 66.2000 ;
	    RECT 56.6000 63.1000 57.0000 68.9000 ;
	    RECT 61.4000 67.8000 61.8000 68.2000 ;
	    RECT 61.4000 67.2000 61.7000 67.8000 ;
	    RECT 59.8000 67.1000 60.2000 67.2000 ;
	    RECT 60.6000 67.1000 61.0000 67.2000 ;
	    RECT 59.8000 66.8000 61.0000 67.1000 ;
	    RECT 61.4000 66.8000 61.8000 67.2000 ;
	    RECT 60.6000 65.8000 61.0000 66.2000 ;
	    RECT 59.0000 64.1000 59.4000 64.2000 ;
	    RECT 59.8000 64.1000 60.2000 64.2000 ;
	    RECT 59.0000 63.8000 60.2000 64.1000 ;
	    RECT 48.6000 62.1000 49.0000 62.2000 ;
	    RECT 49.4000 62.1000 49.8000 62.2000 ;
	    RECT 48.6000 61.8000 49.8000 62.1000 ;
	    RECT 54.2000 58.8000 54.6000 59.2000 ;
	    RECT 49.4000 55.8000 49.8000 56.2000 ;
	    RECT 49.4000 55.1000 49.7000 55.8000 ;
	    RECT 49.4000 54.7000 49.8000 55.1000 ;
	    RECT 50.2000 52.1000 50.6000 57.9000 ;
	    RECT 52.6000 56.8000 53.0000 57.2000 ;
	    RECT 52.6000 56.2000 52.9000 56.8000 ;
	    RECT 51.0000 54.8000 51.4000 55.2000 ;
	    RECT 51.0000 54.2000 51.3000 54.8000 ;
	    RECT 51.0000 53.8000 51.4000 54.2000 ;
	    RECT 47.0000 48.8000 47.4000 49.2000 ;
	    RECT 49.4000 46.8000 49.8000 47.2000 ;
	    RECT 49.4000 46.3000 49.7000 46.8000 ;
	    RECT 49.4000 45.9000 49.8000 46.3000 ;
	    RECT 50.2000 43.1000 50.6000 48.9000 ;
	    RECT 51.0000 47.2000 51.3000 53.8000 ;
	    RECT 51.8000 53.1000 52.2000 55.9000 ;
	    RECT 52.6000 55.8000 53.0000 56.2000 ;
	    RECT 54.2000 54.2000 54.5000 58.8000 ;
	    RECT 53.4000 53.8000 53.8000 54.2000 ;
	    RECT 54.2000 53.8000 54.6000 54.2000 ;
	    RECT 51.0000 46.8000 51.4000 47.2000 ;
	    RECT 51.8000 45.1000 52.2000 47.9000 ;
	    RECT 52.6000 46.8000 53.0000 47.2000 ;
	    RECT 52.6000 46.2000 52.9000 46.8000 ;
	    RECT 52.6000 45.8000 53.0000 46.2000 ;
	    RECT 46.2000 38.8000 46.6000 39.2000 ;
	    RECT 50.2000 36.8000 50.6000 37.2000 ;
	    RECT 15.0000 35.2000 15.3000 35.8000 ;
	    RECT 18.2000 35.2000 18.5000 35.8000 ;
	    RECT 19.8000 35.2000 20.1000 35.8000 ;
	    RECT 30.2000 35.2000 30.5000 35.8000 ;
	    RECT 11.8000 35.1000 12.2000 35.2000 ;
	    RECT 12.6000 35.1000 13.0000 35.2000 ;
	    RECT 11.8000 34.8000 13.0000 35.1000 ;
	    RECT 15.0000 34.8000 15.4000 35.2000 ;
	    RECT 18.2000 34.8000 18.6000 35.2000 ;
	    RECT 19.8000 34.8000 20.2000 35.2000 ;
	    RECT 23.8000 34.8000 24.2000 35.2000 ;
	    RECT 27.0000 35.1000 27.4000 35.2000 ;
	    RECT 27.8000 35.1000 28.2000 35.2000 ;
	    RECT 27.0000 34.8000 28.2000 35.1000 ;
	    RECT 30.2000 34.8000 30.6000 35.2000 ;
	    RECT 31.0000 34.8000 31.4000 35.2000 ;
	    RECT 23.8000 34.2000 24.1000 34.8000 ;
	    RECT 31.0000 34.2000 31.3000 34.8000 ;
	    RECT 36.6000 34.2000 36.9000 35.9000 ;
	    RECT 37.4000 35.8000 37.8000 36.2000 ;
	    RECT 39.9000 35.9000 40.3000 36.3000 ;
	    RECT 38.6000 34.2000 39.0000 34.3000 ;
	    RECT 7.8000 33.9000 10.6000 34.2000 ;
	    RECT 7.8000 33.5000 8.2000 33.6000 ;
	    RECT 9.5000 33.5000 9.9000 33.6000 ;
	    RECT 10.3000 33.5000 10.6000 33.9000 ;
	    RECT 14.2000 34.1000 14.6000 34.2000 ;
	    RECT 15.0000 34.1000 15.4000 34.2000 ;
	    RECT 14.2000 33.8000 15.4000 34.1000 ;
	    RECT 15.8000 34.1000 16.2000 34.2000 ;
	    RECT 16.6000 34.1000 17.0000 34.2000 ;
	    RECT 15.8000 33.8000 17.0000 34.1000 ;
	    RECT 19.8000 34.1000 20.2000 34.2000 ;
	    RECT 20.6000 34.1000 21.0000 34.2000 ;
	    RECT 19.8000 33.8000 21.0000 34.1000 ;
	    RECT 23.8000 33.8000 24.2000 34.2000 ;
	    RECT 24.6000 34.1000 25.0000 34.2000 ;
	    RECT 25.4000 34.1000 25.8000 34.2000 ;
	    RECT 24.6000 33.8000 25.8000 34.1000 ;
	    RECT 31.0000 33.8000 31.4000 34.2000 ;
	    RECT 36.6000 33.9000 39.0000 34.2000 ;
	    RECT 7.1000 33.2000 9.9000 33.5000 ;
	    RECT 7.1000 33.1000 7.5000 33.2000 ;
	    RECT 10.2000 33.1000 10.6000 33.5000 ;
	    RECT 36.6000 33.5000 36.9000 33.9000 ;
	    RECT 40.0000 33.5000 40.3000 35.9000 ;
	    RECT 49.4000 35.8000 49.8000 36.2000 ;
	    RECT 49.4000 35.2000 49.7000 35.8000 ;
	    RECT 50.2000 35.2000 50.5000 36.8000 ;
	    RECT 44.6000 35.1000 45.0000 35.2000 ;
	    RECT 45.4000 35.1000 45.8000 35.2000 ;
	    RECT 44.6000 34.8000 45.8000 35.1000 ;
	    RECT 47.0000 34.8000 47.4000 35.2000 ;
	    RECT 49.4000 34.8000 49.8000 35.2000 ;
	    RECT 50.2000 34.8000 50.6000 35.2000 ;
	    RECT 47.0000 34.2000 47.3000 34.8000 ;
	    RECT 18.2000 32.8000 18.6000 33.2000 ;
	    RECT 23.8000 32.8000 24.2000 33.2000 ;
	    RECT 36.6000 33.1000 37.0000 33.5000 ;
	    RECT 39.9000 33.1000 40.3000 33.5000 ;
	    RECT 41.4000 33.8000 41.8000 34.2000 ;
	    RECT 44.6000 34.1000 45.0000 34.2000 ;
	    RECT 45.4000 34.1000 45.8000 34.2000 ;
	    RECT 44.6000 33.8000 45.8000 34.1000 ;
	    RECT 47.0000 33.8000 47.4000 34.2000 ;
	    RECT 41.4000 33.2000 41.7000 33.8000 ;
	    RECT 41.4000 32.8000 41.8000 33.2000 ;
	    RECT 9.4000 31.8000 9.8000 32.2000 ;
	    RECT 8.6000 29.8000 9.0000 30.2000 ;
	    RECT 8.6000 29.2000 8.9000 29.8000 ;
	    RECT 8.6000 28.8000 9.0000 29.2000 ;
	    RECT 9.4000 27.2000 9.7000 31.8000 ;
	    RECT 15.0000 28.8000 15.4000 29.2000 ;
	    RECT 15.0000 28.2000 15.3000 28.8000 ;
	    RECT 18.2000 28.2000 18.5000 32.8000 ;
	    RECT 23.8000 32.2000 24.1000 32.8000 ;
	    RECT 22.2000 31.8000 22.6000 32.2000 ;
	    RECT 23.8000 31.8000 24.2000 32.2000 ;
	    RECT 29.4000 31.8000 29.8000 32.2000 ;
	    RECT 22.2000 29.2000 22.5000 31.8000 ;
	    RECT 20.6000 28.8000 21.0000 29.2000 ;
	    RECT 22.2000 28.8000 22.6000 29.2000 ;
	    RECT 20.6000 28.2000 20.9000 28.8000 ;
	    RECT 15.0000 27.8000 15.4000 28.2000 ;
	    RECT 16.6000 27.8000 17.0000 28.2000 ;
	    RECT 18.2000 27.8000 18.6000 28.2000 ;
	    RECT 20.6000 27.8000 21.0000 28.2000 ;
	    RECT 21.4000 28.1000 21.8000 28.2000 ;
	    RECT 22.2000 28.1000 22.6000 28.2000 ;
	    RECT 21.4000 27.8000 22.6000 28.1000 ;
	    RECT 16.6000 27.2000 16.9000 27.8000 ;
	    RECT 18.2000 27.2000 18.5000 27.8000 ;
	    RECT 29.4000 27.2000 29.7000 31.8000 ;
	    RECT 41.4000 29.1000 41.7000 32.8000 ;
	    RECT 43.8000 31.8000 44.2000 32.2000 ;
	    RECT 42.2000 29.1000 42.6000 29.2000 ;
	    RECT 3.8000 26.8000 4.2000 27.2000 ;
	    RECT 7.0000 27.1000 7.4000 27.2000 ;
	    RECT 7.8000 27.1000 8.2000 27.2000 ;
	    RECT 7.0000 26.8000 8.2000 27.1000 ;
	    RECT 9.4000 26.8000 9.8000 27.2000 ;
	    RECT 11.8000 26.8000 12.2000 27.2000 ;
	    RECT 16.6000 26.8000 17.0000 27.2000 ;
	    RECT 18.2000 26.8000 18.6000 27.2000 ;
	    RECT 25.4000 26.8000 25.8000 27.2000 ;
	    RECT 29.4000 26.8000 29.8000 27.2000 ;
	    RECT 31.0000 26.8000 31.4000 27.2000 ;
	    RECT 3.8000 26.2000 4.1000 26.8000 ;
	    RECT 11.8000 26.2000 12.1000 26.8000 ;
	    RECT 25.4000 26.2000 25.7000 26.8000 ;
	    RECT 31.0000 26.2000 31.3000 26.8000 ;
	    RECT 3.8000 25.8000 4.2000 26.2000 ;
	    RECT 6.2000 25.8000 6.6000 26.2000 ;
	    RECT 10.2000 26.1000 10.6000 26.2000 ;
	    RECT 11.0000 26.1000 11.4000 26.2000 ;
	    RECT 10.2000 25.8000 11.4000 26.1000 ;
	    RECT 11.8000 25.8000 12.2000 26.2000 ;
	    RECT 17.4000 25.8000 17.8000 26.2000 ;
	    RECT 25.4000 25.8000 25.8000 26.2000 ;
	    RECT 27.0000 26.1000 27.4000 26.2000 ;
	    RECT 27.8000 26.1000 28.2000 26.2000 ;
	    RECT 27.0000 25.8000 28.2000 26.1000 ;
	    RECT 29.4000 25.8000 29.8000 26.2000 ;
	    RECT 31.0000 25.8000 31.4000 26.2000 ;
	    RECT 6.2000 25.2000 6.5000 25.8000 ;
	    RECT 17.4000 25.2000 17.7000 25.8000 ;
	    RECT 29.4000 25.2000 29.7000 25.8000 ;
	    RECT 6.2000 24.8000 6.6000 25.2000 ;
	    RECT 17.4000 24.8000 17.8000 25.2000 ;
	    RECT 19.8000 25.1000 20.2000 25.2000 ;
	    RECT 20.6000 25.1000 21.0000 25.2000 ;
	    RECT 19.8000 24.8000 21.0000 25.1000 ;
	    RECT 23.8000 25.1000 24.2000 25.2000 ;
	    RECT 24.6000 25.1000 25.0000 25.2000 ;
	    RECT 23.8000 24.8000 25.0000 25.1000 ;
	    RECT 29.4000 24.8000 29.8000 25.2000 ;
	    RECT 33.4000 25.1000 33.8000 27.9000 ;
	    RECT 35.0000 23.1000 35.4000 28.9000 ;
	    RECT 36.6000 26.8000 37.0000 27.2000 ;
	    RECT 36.6000 26.2000 36.9000 26.8000 ;
	    RECT 36.6000 25.8000 37.0000 26.2000 ;
	    RECT 39.0000 25.8000 39.4000 26.2000 ;
	    RECT 39.0000 23.2000 39.3000 25.8000 ;
	    RECT 35.8000 22.8000 36.2000 23.2000 ;
	    RECT 39.0000 22.8000 39.4000 23.2000 ;
	    RECT 39.8000 23.1000 40.2000 28.9000 ;
	    RECT 41.4000 28.8000 42.6000 29.1000 ;
	    RECT 43.0000 25.1000 43.4000 27.9000 ;
	    RECT 43.8000 27.2000 44.1000 31.8000 ;
	    RECT 43.8000 26.8000 44.2000 27.2000 ;
	    RECT 43.8000 25.8000 44.2000 26.2000 ;
	    RECT 2.2000 15.1000 2.6000 15.2000 ;
	    RECT 3.0000 15.1000 3.4000 15.2000 ;
	    RECT 2.2000 14.8000 3.4000 15.1000 ;
	    RECT 3.8000 14.8000 4.2000 15.2000 ;
	    RECT 1.4000 12.8000 1.8000 13.2000 ;
	    RECT 1.4000 12.2000 1.7000 12.8000 ;
	    RECT 1.4000 11.8000 1.8000 12.2000 ;
	    RECT 2.2000 11.8000 2.6000 12.2000 ;
	    RECT 2.2000 6.2000 2.5000 11.8000 ;
	    RECT 3.8000 6.2000 4.1000 14.8000 ;
	    RECT 4.6000 12.8000 5.0000 13.2000 ;
	    RECT 4.6000 12.2000 4.9000 12.8000 ;
	    RECT 4.6000 11.8000 5.0000 12.2000 ;
	    RECT 7.0000 12.1000 7.4000 17.9000 ;
	    RECT 9.4000 15.1000 9.8000 15.2000 ;
	    RECT 10.2000 15.1000 10.6000 15.2000 ;
	    RECT 9.4000 14.8000 10.6000 15.1000 ;
	    RECT 11.8000 12.1000 12.2000 17.9000 ;
	    RECT 12.6000 13.8000 13.0000 14.2000 ;
	    RECT 12.6000 9.2000 12.9000 13.8000 ;
	    RECT 13.4000 13.1000 13.8000 15.9000 ;
	    RECT 14.2000 14.8000 14.6000 15.2000 ;
	    RECT 15.8000 14.8000 16.2000 15.2000 ;
	    RECT 5.4000 8.8000 5.8000 9.2000 ;
	    RECT 8.6000 9.1000 9.0000 9.2000 ;
	    RECT 9.4000 9.1000 9.8000 9.2000 ;
	    RECT 8.6000 8.8000 9.8000 9.1000 ;
	    RECT 5.4000 8.2000 5.7000 8.8000 ;
	    RECT 5.4000 7.8000 5.8000 8.2000 ;
	    RECT 5.4000 6.2000 5.7000 7.8000 ;
	    RECT 2.2000 5.8000 2.6000 6.2000 ;
	    RECT 3.8000 5.8000 4.2000 6.2000 ;
	    RECT 5.4000 5.8000 5.8000 6.2000 ;
	    RECT 8.6000 6.1000 9.0000 6.2000 ;
	    RECT 9.4000 6.1000 9.8000 6.2000 ;
	    RECT 8.6000 5.8000 9.8000 6.1000 ;
	    RECT 8.6000 4.8000 9.0000 5.2000 ;
	    RECT 8.6000 4.2000 8.9000 4.8000 ;
	    RECT 8.6000 3.8000 9.0000 4.2000 ;
	    RECT 11.8000 3.1000 12.2000 8.9000 ;
	    RECT 12.6000 8.8000 13.0000 9.2000 ;
	    RECT 14.2000 6.2000 14.5000 14.8000 ;
	    RECT 15.8000 14.2000 16.1000 14.8000 ;
	    RECT 15.8000 13.8000 16.2000 14.2000 ;
	    RECT 19.8000 12.8000 20.2000 13.2000 ;
	    RECT 15.8000 8.8000 16.2000 9.2000 ;
	    RECT 15.8000 8.2000 16.1000 8.8000 ;
	    RECT 15.8000 7.8000 16.2000 8.2000 ;
	    RECT 14.2000 5.8000 14.6000 6.2000 ;
	    RECT 15.0000 5.8000 15.4000 6.2000 ;
	    RECT 15.0000 5.2000 15.3000 5.8000 ;
	    RECT 15.0000 4.8000 15.4000 5.2000 ;
	    RECT 16.6000 3.1000 17.0000 8.9000 ;
	    RECT 18.2000 5.1000 18.6000 7.9000 ;
	    RECT 19.8000 6.1000 20.1000 12.8000 ;
	    RECT 20.6000 12.1000 21.0000 17.9000 ;
	    RECT 23.0000 15.1000 23.4000 15.2000 ;
	    RECT 23.8000 15.1000 24.2000 15.2000 ;
	    RECT 23.0000 14.8000 24.2000 15.1000 ;
	    RECT 25.4000 12.1000 25.8000 17.9000 ;
	    RECT 26.2000 14.8000 26.6000 15.2000 ;
	    RECT 26.2000 14.2000 26.5000 14.8000 ;
	    RECT 26.2000 13.8000 26.6000 14.2000 ;
	    RECT 26.2000 9.2000 26.5000 13.8000 ;
	    RECT 27.0000 13.1000 27.4000 15.9000 ;
	    RECT 30.2000 13.1000 30.6000 15.9000 ;
	    RECT 31.0000 14.8000 31.4000 15.2000 ;
	    RECT 31.0000 14.2000 31.3000 14.8000 ;
	    RECT 31.0000 13.8000 31.4000 14.2000 ;
	    RECT 31.8000 12.1000 32.2000 17.9000 ;
	    RECT 35.8000 15.2000 36.1000 22.8000 ;
	    RECT 43.8000 19.2000 44.1000 25.8000 ;
	    RECT 44.6000 23.1000 45.0000 28.9000 ;
	    RECT 45.4000 25.9000 45.8000 26.3000 ;
	    RECT 47.0000 26.2000 47.3000 33.8000 ;
	    RECT 45.4000 25.2000 45.7000 25.9000 ;
	    RECT 47.0000 25.8000 47.4000 26.2000 ;
	    RECT 48.6000 25.8000 49.0000 26.2000 ;
	    RECT 45.4000 24.8000 45.8000 25.2000 ;
	    RECT 46.2000 21.8000 46.6000 22.2000 ;
	    RECT 43.8000 18.8000 44.2000 19.2000 ;
	    RECT 33.4000 15.1000 33.8000 15.2000 ;
	    RECT 34.2000 15.1000 34.6000 15.2000 ;
	    RECT 33.4000 14.8000 34.6000 15.1000 ;
	    RECT 35.8000 14.8000 36.2000 15.2000 ;
	    RECT 36.6000 12.1000 37.0000 17.9000 ;
	    RECT 39.8000 15.8000 40.2000 16.2000 ;
	    RECT 39.8000 15.2000 40.1000 15.8000 ;
	    RECT 39.8000 14.8000 40.2000 15.2000 ;
	    RECT 43.0000 15.1000 43.4000 15.2000 ;
	    RECT 43.8000 15.1000 44.2000 15.2000 ;
	    RECT 43.0000 14.8000 44.2000 15.1000 ;
	    RECT 41.4000 13.8000 41.8000 14.2000 ;
	    RECT 41.4000 12.2000 41.7000 13.8000 ;
	    RECT 43.0000 13.2000 43.3000 14.8000 ;
	    RECT 46.2000 13.2000 46.5000 21.8000 ;
	    RECT 47.0000 15.2000 47.3000 25.8000 ;
	    RECT 48.6000 23.2000 48.9000 25.8000 ;
	    RECT 48.6000 22.8000 49.0000 23.2000 ;
	    RECT 49.4000 23.1000 49.8000 28.9000 ;
	    RECT 47.0000 14.8000 47.4000 15.2000 ;
	    RECT 50.2000 14.2000 50.5000 34.8000 ;
	    RECT 52.6000 32.1000 53.0000 37.9000 ;
	    RECT 53.4000 35.2000 53.7000 53.8000 ;
	    RECT 55.0000 52.8000 55.4000 53.2000 ;
	    RECT 54.2000 48.8000 54.6000 49.2000 ;
	    RECT 54.2000 47.2000 54.5000 48.8000 ;
	    RECT 55.0000 48.2000 55.3000 52.8000 ;
	    RECT 57.4000 51.8000 57.8000 52.2000 ;
	    RECT 59.8000 52.1000 60.2000 57.9000 ;
	    RECT 57.4000 51.2000 57.7000 51.8000 ;
	    RECT 57.4000 50.8000 57.8000 51.2000 ;
	    RECT 57.4000 48.8000 57.8000 49.2000 ;
	    RECT 57.4000 48.2000 57.7000 48.8000 ;
	    RECT 60.6000 48.2000 60.9000 65.8000 ;
	    RECT 61.4000 52.2000 61.7000 66.8000 ;
	    RECT 62.2000 54.2000 62.5000 70.8000 ;
	    RECT 63.0000 65.8000 63.4000 66.2000 ;
	    RECT 64.6000 65.8000 65.0000 66.2000 ;
	    RECT 63.0000 61.2000 63.3000 65.8000 ;
	    RECT 64.6000 65.2000 64.9000 65.8000 ;
	    RECT 63.8000 64.8000 64.2000 65.2000 ;
	    RECT 64.6000 64.8000 65.0000 65.2000 ;
	    RECT 63.8000 64.2000 64.1000 64.8000 ;
	    RECT 65.4000 64.2000 65.7000 73.8000 ;
	    RECT 67.0000 72.1000 67.4000 77.9000 ;
	    RECT 72.6000 76.8000 73.0000 77.2000 ;
	    RECT 72.6000 76.2000 72.9000 76.8000 ;
	    RECT 67.8000 73.8000 68.2000 74.2000 ;
	    RECT 67.8000 71.2000 68.1000 73.8000 ;
	    RECT 68.6000 73.1000 69.0000 75.9000 ;
	    RECT 71.8000 75.8000 72.2000 76.2000 ;
	    RECT 72.6000 75.8000 73.0000 76.2000 ;
	    RECT 71.8000 75.2000 72.1000 75.8000 ;
	    RECT 72.6000 75.2000 72.9000 75.8000 ;
	    RECT 74.2000 75.2000 74.5000 81.8000 ;
	    RECT 69.4000 74.8000 69.8000 75.2000 ;
	    RECT 71.8000 74.8000 72.2000 75.2000 ;
	    RECT 72.6000 74.8000 73.0000 75.2000 ;
	    RECT 74.2000 74.8000 74.6000 75.2000 ;
	    RECT 69.4000 74.2000 69.7000 74.8000 ;
	    RECT 69.4000 73.8000 69.8000 74.2000 ;
	    RECT 71.8000 73.8000 72.2000 74.2000 ;
	    RECT 69.4000 72.8000 69.8000 73.2000 ;
	    RECT 67.8000 70.8000 68.2000 71.2000 ;
	    RECT 69.4000 67.2000 69.7000 72.8000 ;
	    RECT 70.2000 71.8000 70.6000 72.2000 ;
	    RECT 66.2000 67.1000 66.6000 67.2000 ;
	    RECT 67.0000 67.1000 67.4000 67.2000 ;
	    RECT 66.2000 66.8000 67.4000 67.1000 ;
	    RECT 69.4000 66.8000 69.8000 67.2000 ;
	    RECT 67.8000 66.1000 68.2000 66.2000 ;
	    RECT 68.6000 66.1000 69.0000 66.2000 ;
	    RECT 67.8000 65.8000 69.0000 66.1000 ;
	    RECT 69.4000 65.1000 69.8000 65.2000 ;
	    RECT 70.2000 65.1000 70.5000 71.8000 ;
	    RECT 69.4000 64.8000 70.5000 65.1000 ;
	    RECT 63.8000 63.8000 64.2000 64.2000 ;
	    RECT 65.4000 63.8000 65.8000 64.2000 ;
	    RECT 63.0000 60.8000 63.4000 61.2000 ;
	    RECT 65.4000 59.2000 65.7000 63.8000 ;
	    RECT 66.2000 61.8000 66.6000 62.2000 ;
	    RECT 65.4000 58.8000 65.8000 59.2000 ;
	    RECT 63.0000 55.0000 63.4000 55.1000 ;
	    RECT 63.8000 55.0000 64.2000 55.1000 ;
	    RECT 63.0000 54.7000 64.2000 55.0000 ;
	    RECT 62.2000 53.8000 62.6000 54.2000 ;
	    RECT 61.4000 51.8000 61.8000 52.2000 ;
	    RECT 64.6000 52.1000 65.0000 57.9000 ;
	    RECT 66.2000 57.2000 66.5000 61.8000 ;
	    RECT 66.2000 56.8000 66.6000 57.2000 ;
	    RECT 69.4000 56.8000 69.8000 57.2000 ;
	    RECT 66.2000 53.1000 66.6000 55.9000 ;
	    RECT 69.4000 55.2000 69.7000 56.8000 ;
	    RECT 70.2000 56.2000 70.5000 64.8000 ;
	    RECT 71.8000 70.2000 72.1000 73.8000 ;
	    RECT 74.2000 73.2000 74.5000 74.8000 ;
	    RECT 75.0000 74.2000 75.3000 84.8000 ;
	    RECT 77.4000 79.2000 77.7000 85.8000 ;
	    RECT 79.0000 85.1000 79.4000 87.9000 ;
	    RECT 77.4000 78.8000 77.8000 79.2000 ;
	    RECT 79.8000 77.2000 80.1000 91.8000 ;
	    RECT 82.2000 89.2000 82.5000 94.8000 ;
	    RECT 84.6000 93.2000 84.9000 94.8000 ;
	    RECT 84.6000 92.8000 85.0000 93.2000 ;
	    RECT 86.2000 90.2000 86.5000 94.8000 ;
	    RECT 88.6000 94.2000 88.9000 94.8000 ;
	    RECT 89.4000 94.2000 89.7000 104.8000 ;
	    RECT 95.0000 104.2000 95.3000 107.8000 ;
	    RECT 95.8000 107.2000 96.1000 107.8000 ;
	    RECT 99.0000 107.2000 99.3000 107.8000 ;
	    RECT 95.8000 106.8000 96.2000 107.2000 ;
	    RECT 97.4000 106.8000 97.8000 107.2000 ;
	    RECT 99.0000 106.8000 99.4000 107.2000 ;
	    RECT 100.6000 107.1000 101.0000 107.2000 ;
	    RECT 101.4000 107.1000 101.7000 109.8000 ;
	    RECT 103.0000 108.2000 103.3000 111.8000 ;
	    RECT 107.0000 110.2000 107.3000 111.8000 ;
	    RECT 107.0000 109.8000 107.4000 110.2000 ;
	    RECT 111.0000 108.8000 111.4000 109.2000 ;
	    RECT 103.0000 107.8000 103.4000 108.2000 ;
	    RECT 105.4000 107.8000 105.8000 108.2000 ;
	    RECT 100.6000 106.8000 101.7000 107.1000 ;
	    RECT 103.0000 107.1000 103.4000 107.2000 ;
	    RECT 103.8000 107.1000 104.2000 107.2000 ;
	    RECT 103.0000 106.8000 104.2000 107.1000 ;
	    RECT 97.4000 106.2000 97.7000 106.8000 ;
	    RECT 95.8000 105.8000 96.2000 106.2000 ;
	    RECT 97.4000 105.8000 97.8000 106.2000 ;
	    RECT 95.8000 105.2000 96.1000 105.8000 ;
	    RECT 105.4000 105.2000 105.7000 107.8000 ;
	    RECT 111.0000 107.2000 111.3000 108.8000 ;
	    RECT 106.2000 107.1000 106.6000 107.2000 ;
	    RECT 107.0000 107.1000 107.4000 107.2000 ;
	    RECT 106.2000 106.8000 107.4000 107.1000 ;
	    RECT 107.8000 106.8000 108.2000 107.2000 ;
	    RECT 111.0000 106.8000 111.4000 107.2000 ;
	    RECT 107.8000 106.2000 108.1000 106.8000 ;
	    RECT 107.8000 105.8000 108.2000 106.2000 ;
	    RECT 111.0000 106.1000 111.4000 106.2000 ;
	    RECT 111.8000 106.1000 112.1000 111.8000 ;
	    RECT 111.0000 105.8000 112.1000 106.1000 ;
	    RECT 113.4000 106.2000 113.7000 112.8000 ;
	    RECT 114.2000 112.1000 114.6000 112.2000 ;
	    RECT 115.0000 112.1000 115.4000 112.2000 ;
	    RECT 114.2000 111.8000 115.4000 112.1000 ;
	    RECT 115.8000 106.8000 116.2000 107.2000 ;
	    RECT 115.8000 106.2000 116.1000 106.8000 ;
	    RECT 113.4000 105.8000 113.8000 106.2000 ;
	    RECT 115.0000 105.8000 115.4000 106.2000 ;
	    RECT 115.8000 105.8000 116.2000 106.2000 ;
	    RECT 95.8000 104.8000 96.2000 105.2000 ;
	    RECT 96.6000 105.1000 97.0000 105.2000 ;
	    RECT 97.4000 105.1000 97.8000 105.2000 ;
	    RECT 96.6000 104.8000 97.8000 105.1000 ;
	    RECT 105.4000 104.8000 105.8000 105.2000 ;
	    RECT 108.6000 104.8000 109.0000 105.2000 ;
	    RECT 111.8000 104.8000 112.2000 105.2000 ;
	    RECT 95.0000 103.8000 95.4000 104.2000 ;
	    RECT 107.0000 104.1000 107.4000 104.2000 ;
	    RECT 107.8000 104.1000 108.2000 104.2000 ;
	    RECT 107.0000 103.8000 108.2000 104.1000 ;
	    RECT 108.6000 102.2000 108.9000 104.8000 ;
	    RECT 111.8000 104.2000 112.1000 104.8000 ;
	    RECT 111.8000 103.8000 112.2000 104.2000 ;
	    RECT 115.0000 103.2000 115.3000 105.8000 ;
	    RECT 116.6000 104.2000 116.9000 112.8000 ;
	    RECT 118.2000 111.8000 118.6000 112.2000 ;
	    RECT 118.2000 108.2000 118.5000 111.8000 ;
	    RECT 120.6000 109.2000 120.9000 112.8000 ;
	    RECT 123.8000 109.2000 124.1000 112.8000 ;
	    RECT 125.4000 109.2000 125.7000 114.8000 ;
	    RECT 126.2000 113.8000 126.6000 114.2000 ;
	    RECT 126.2000 113.2000 126.5000 113.8000 ;
	    RECT 126.2000 112.8000 126.6000 113.2000 ;
	    RECT 120.6000 108.8000 121.0000 109.2000 ;
	    RECT 123.8000 108.8000 124.2000 109.2000 ;
	    RECT 125.4000 108.8000 125.8000 109.2000 ;
	    RECT 118.2000 107.8000 118.6000 108.2000 ;
	    RECT 119.0000 107.8000 119.4000 108.2000 ;
	    RECT 118.2000 107.2000 118.5000 107.8000 ;
	    RECT 119.0000 107.2000 119.3000 107.8000 ;
	    RECT 118.2000 106.8000 118.6000 107.2000 ;
	    RECT 119.0000 106.8000 119.4000 107.2000 ;
	    RECT 123.0000 107.1000 123.4000 107.2000 ;
	    RECT 123.8000 107.1000 124.2000 107.2000 ;
	    RECT 123.0000 106.8000 124.2000 107.1000 ;
	    RECT 124.6000 106.8000 125.0000 107.2000 ;
	    RECT 122.2000 105.8000 122.6000 106.2000 ;
	    RECT 119.8000 105.1000 120.2000 105.2000 ;
	    RECT 120.6000 105.1000 121.0000 105.2000 ;
	    RECT 119.8000 104.8000 121.0000 105.1000 ;
	    RECT 116.6000 103.8000 117.0000 104.2000 ;
	    RECT 115.0000 102.8000 115.4000 103.2000 ;
	    RECT 94.2000 101.8000 94.6000 102.2000 ;
	    RECT 98.2000 101.8000 98.6000 102.2000 ;
	    RECT 103.8000 101.8000 104.2000 102.2000 ;
	    RECT 108.6000 101.8000 109.0000 102.2000 ;
	    RECT 118.2000 101.8000 118.6000 102.2000 ;
	    RECT 91.8000 94.8000 92.2000 95.2000 ;
	    RECT 88.6000 93.8000 89.0000 94.2000 ;
	    RECT 89.4000 93.8000 89.8000 94.2000 ;
	    RECT 91.8000 91.2000 92.1000 94.8000 ;
	    RECT 93.4000 93.8000 93.8000 94.2000 ;
	    RECT 93.4000 93.2000 93.7000 93.8000 ;
	    RECT 93.4000 92.8000 93.8000 93.2000 ;
	    RECT 91.8000 90.8000 92.2000 91.2000 ;
	    RECT 86.2000 89.8000 86.6000 90.2000 ;
	    RECT 87.8000 89.8000 88.2000 90.2000 ;
	    RECT 88.6000 89.8000 89.0000 90.2000 ;
	    RECT 87.8000 89.2000 88.1000 89.8000 ;
	    RECT 88.6000 89.2000 88.9000 89.8000 ;
	    RECT 93.4000 89.2000 93.7000 92.8000 ;
	    RECT 80.6000 83.1000 81.0000 88.9000 ;
	    RECT 81.4000 88.8000 81.8000 89.2000 ;
	    RECT 82.2000 88.8000 82.6000 89.2000 ;
	    RECT 81.4000 86.3000 81.7000 88.8000 ;
	    RECT 84.6000 87.8000 85.0000 88.2000 ;
	    RECT 81.4000 85.9000 81.8000 86.3000 ;
	    RECT 84.6000 86.2000 84.9000 87.8000 ;
	    RECT 84.6000 85.8000 85.0000 86.2000 ;
	    RECT 75.8000 76.8000 76.2000 77.2000 ;
	    RECT 79.8000 76.8000 80.2000 77.2000 ;
	    RECT 75.8000 76.2000 76.1000 76.8000 ;
	    RECT 75.8000 75.8000 76.2000 76.2000 ;
	    RECT 75.0000 73.8000 75.4000 74.2000 ;
	    RECT 74.2000 72.8000 74.6000 73.2000 ;
	    RECT 73.4000 70.8000 73.8000 71.2000 ;
	    RECT 71.8000 69.8000 72.2000 70.2000 ;
	    RECT 71.8000 68.2000 72.1000 69.8000 ;
	    RECT 71.8000 67.8000 72.2000 68.2000 ;
	    RECT 71.8000 64.2000 72.1000 67.8000 ;
	    RECT 72.6000 65.1000 73.0000 67.9000 ;
	    RECT 73.4000 67.2000 73.7000 70.8000 ;
	    RECT 75.0000 69.2000 75.3000 73.8000 ;
	    RECT 75.8000 72.2000 76.1000 75.8000 ;
	    RECT 76.6000 75.1000 77.0000 75.2000 ;
	    RECT 77.4000 75.1000 77.8000 75.2000 ;
	    RECT 76.6000 74.8000 77.8000 75.1000 ;
	    RECT 78.2000 74.8000 78.6000 75.2000 ;
	    RECT 78.2000 74.2000 78.5000 74.8000 ;
	    RECT 78.2000 73.8000 78.6000 74.2000 ;
	    RECT 75.8000 71.8000 76.2000 72.2000 ;
	    RECT 79.0000 71.8000 79.4000 72.2000 ;
	    RECT 81.4000 72.1000 81.8000 77.9000 ;
	    RECT 84.6000 74.2000 84.9000 85.8000 ;
	    RECT 85.4000 83.1000 85.8000 88.9000 ;
	    RECT 87.8000 88.8000 88.2000 89.2000 ;
	    RECT 88.6000 88.8000 89.0000 89.2000 ;
	    RECT 91.0000 83.1000 91.4000 88.9000 ;
	    RECT 93.4000 88.8000 93.8000 89.2000 ;
	    RECT 94.2000 86.2000 94.5000 101.8000 ;
	    RECT 98.2000 100.2000 98.5000 101.8000 ;
	    RECT 102.2000 100.8000 102.6000 101.2000 ;
	    RECT 98.2000 99.8000 98.6000 100.2000 ;
	    RECT 98.2000 97.8000 98.6000 98.2000 ;
	    RECT 100.6000 97.8000 101.0000 98.2000 ;
	    RECT 95.0000 95.8000 95.4000 96.2000 ;
	    RECT 95.8000 95.8000 96.2000 96.2000 ;
	    RECT 97.4000 95.8000 97.8000 96.2000 ;
	    RECT 95.0000 95.2000 95.3000 95.8000 ;
	    RECT 95.0000 94.8000 95.4000 95.2000 ;
	    RECT 95.8000 94.1000 96.1000 95.8000 ;
	    RECT 97.4000 95.2000 97.7000 95.8000 ;
	    RECT 97.4000 94.8000 97.8000 95.2000 ;
	    RECT 98.2000 94.2000 98.5000 97.8000 ;
	    RECT 100.6000 94.2000 100.9000 97.8000 ;
	    RECT 101.4000 94.8000 101.8000 95.2000 ;
	    RECT 101.4000 94.2000 101.7000 94.8000 ;
	    RECT 95.0000 93.8000 96.1000 94.1000 ;
	    RECT 96.6000 93.8000 97.0000 94.2000 ;
	    RECT 98.2000 93.8000 98.6000 94.2000 ;
	    RECT 99.0000 94.1000 99.4000 94.2000 ;
	    RECT 99.8000 94.1000 100.2000 94.2000 ;
	    RECT 99.0000 93.8000 100.2000 94.1000 ;
	    RECT 100.6000 93.8000 101.0000 94.2000 ;
	    RECT 101.4000 93.8000 101.8000 94.2000 ;
	    RECT 94.2000 85.8000 94.6000 86.2000 ;
	    RECT 85.4000 74.7000 85.8000 75.1000 ;
	    RECT 84.6000 73.8000 85.0000 74.2000 ;
	    RECT 83.8000 72.8000 84.2000 73.2000 ;
	    RECT 79.0000 71.2000 79.3000 71.8000 ;
	    RECT 83.8000 71.2000 84.1000 72.8000 ;
	    RECT 79.0000 70.8000 79.4000 71.2000 ;
	    RECT 83.8000 70.8000 84.2000 71.2000 ;
	    RECT 85.4000 71.1000 85.7000 74.7000 ;
	    RECT 86.2000 72.1000 86.6000 77.9000 ;
	    RECT 95.0000 77.2000 95.3000 93.8000 ;
	    RECT 96.6000 93.2000 96.9000 93.8000 ;
	    RECT 96.6000 92.8000 97.0000 93.2000 ;
	    RECT 98.2000 93.1000 98.6000 93.2000 ;
	    RECT 99.0000 93.1000 99.4000 93.2000 ;
	    RECT 98.2000 92.8000 99.4000 93.1000 ;
	    RECT 100.6000 89.8000 101.0000 90.2000 ;
	    RECT 95.8000 83.1000 96.2000 88.9000 ;
	    RECT 96.6000 87.8000 97.0000 88.2000 ;
	    RECT 96.6000 87.2000 96.9000 87.8000 ;
	    RECT 96.6000 86.8000 97.0000 87.2000 ;
	    RECT 97.4000 85.1000 97.8000 87.9000 ;
	    RECT 98.2000 87.1000 98.6000 87.2000 ;
	    RECT 99.0000 87.1000 99.4000 87.2000 ;
	    RECT 98.2000 86.8000 99.4000 87.1000 ;
	    RECT 98.2000 85.8000 98.6000 86.2000 ;
	    RECT 95.0000 76.8000 95.4000 77.2000 ;
	    RECT 95.0000 76.2000 95.3000 76.8000 ;
	    RECT 87.8000 73.1000 88.2000 75.9000 ;
	    RECT 89.4000 75.8000 89.8000 76.2000 ;
	    RECT 90.2000 75.8000 90.6000 76.2000 ;
	    RECT 95.0000 75.8000 95.4000 76.2000 ;
	    RECT 89.4000 75.2000 89.7000 75.8000 ;
	    RECT 89.4000 74.8000 89.8000 75.2000 ;
	    RECT 90.2000 74.2000 90.5000 75.8000 ;
	    RECT 93.4000 74.8000 93.8000 75.2000 ;
	    RECT 95.0000 75.1000 95.4000 75.2000 ;
	    RECT 95.8000 75.1000 96.2000 75.2000 ;
	    RECT 95.0000 74.8000 96.2000 75.1000 ;
	    RECT 97.4000 74.8000 97.8000 75.2000 ;
	    RECT 90.2000 73.8000 90.6000 74.2000 ;
	    RECT 91.8000 74.1000 92.2000 74.2000 ;
	    RECT 92.6000 74.1000 93.0000 74.2000 ;
	    RECT 91.8000 73.8000 93.0000 74.1000 ;
	    RECT 85.4000 70.8000 86.5000 71.1000 ;
	    RECT 73.4000 66.8000 73.8000 67.2000 ;
	    RECT 71.8000 63.8000 72.2000 64.2000 ;
	    RECT 71.0000 63.1000 71.4000 63.2000 ;
	    RECT 71.8000 63.1000 72.2000 63.2000 ;
	    RECT 74.2000 63.1000 74.6000 68.9000 ;
	    RECT 75.0000 68.8000 75.4000 69.2000 ;
	    RECT 75.8000 68.8000 76.2000 69.2000 ;
	    RECT 75.0000 65.9000 75.4000 66.3000 ;
	    RECT 75.0000 63.2000 75.3000 65.9000 ;
	    RECT 71.0000 62.8000 72.2000 63.1000 ;
	    RECT 75.0000 62.8000 75.4000 63.2000 ;
	    RECT 71.8000 60.8000 72.2000 61.2000 ;
	    RECT 71.8000 59.2000 72.1000 60.8000 ;
	    RECT 71.8000 58.8000 72.2000 59.2000 ;
	    RECT 70.2000 56.1000 70.6000 56.2000 ;
	    RECT 70.2000 55.8000 71.3000 56.1000 ;
	    RECT 67.0000 55.1000 67.4000 55.2000 ;
	    RECT 67.8000 55.1000 68.2000 55.2000 ;
	    RECT 67.0000 54.8000 68.2000 55.1000 ;
	    RECT 68.6000 54.8000 69.0000 55.2000 ;
	    RECT 69.4000 54.8000 69.8000 55.2000 ;
	    RECT 68.6000 54.2000 68.9000 54.8000 ;
	    RECT 67.0000 53.8000 67.4000 54.2000 ;
	    RECT 68.6000 53.8000 69.0000 54.2000 ;
	    RECT 67.0000 53.2000 67.3000 53.8000 ;
	    RECT 67.0000 52.8000 67.4000 53.2000 ;
	    RECT 69.4000 51.8000 69.8000 52.2000 ;
	    RECT 66.2000 49.8000 66.6000 50.2000 ;
	    RECT 66.2000 49.2000 66.5000 49.8000 ;
	    RECT 69.4000 49.2000 69.7000 51.8000 ;
	    RECT 66.2000 48.8000 66.6000 49.2000 ;
	    RECT 69.4000 48.8000 69.8000 49.2000 ;
	    RECT 55.0000 48.1000 55.4000 48.2000 ;
	    RECT 55.8000 48.1000 56.2000 48.2000 ;
	    RECT 55.0000 47.8000 56.2000 48.1000 ;
	    RECT 57.4000 47.8000 57.8000 48.2000 ;
	    RECT 60.6000 47.8000 61.0000 48.2000 ;
	    RECT 68.6000 48.1000 69.0000 48.2000 ;
	    RECT 69.4000 48.1000 69.8000 48.2000 ;
	    RECT 68.6000 47.8000 69.8000 48.1000 ;
	    RECT 70.2000 47.8000 70.6000 48.2000 ;
	    RECT 70.2000 47.2000 70.5000 47.8000 ;
	    RECT 54.2000 46.8000 54.6000 47.2000 ;
	    RECT 62.2000 47.1000 62.6000 47.2000 ;
	    RECT 63.0000 47.1000 63.4000 47.2000 ;
	    RECT 62.2000 46.8000 63.4000 47.1000 ;
	    RECT 65.4000 47.1000 65.8000 47.2000 ;
	    RECT 66.2000 47.1000 66.6000 47.2000 ;
	    RECT 65.4000 46.8000 66.6000 47.1000 ;
	    RECT 70.2000 46.8000 70.6000 47.2000 ;
	    RECT 55.8000 45.8000 56.2000 46.2000 ;
	    RECT 63.0000 45.8000 63.4000 46.2000 ;
	    RECT 64.6000 46.1000 65.0000 46.2000 ;
	    RECT 65.4000 46.1000 65.8000 46.2000 ;
	    RECT 64.6000 45.8000 65.8000 46.1000 ;
	    RECT 69.4000 46.1000 69.8000 46.2000 ;
	    RECT 70.2000 46.1000 70.6000 46.2000 ;
	    RECT 69.4000 45.8000 70.6000 46.1000 ;
	    RECT 55.8000 42.2000 56.1000 45.8000 ;
	    RECT 55.8000 41.8000 56.2000 42.2000 ;
	    RECT 55.8000 36.2000 56.1000 41.8000 ;
	    RECT 63.0000 39.2000 63.3000 45.8000 ;
	    RECT 69.4000 44.8000 69.8000 45.2000 ;
	    RECT 63.8000 42.8000 64.2000 43.2000 ;
	    RECT 67.0000 42.8000 67.4000 43.2000 ;
	    RECT 56.6000 38.8000 57.0000 39.2000 ;
	    RECT 63.0000 38.8000 63.4000 39.2000 ;
	    RECT 55.8000 35.8000 56.2000 36.2000 ;
	    RECT 53.4000 34.8000 53.8000 35.2000 ;
	    RECT 56.6000 35.1000 56.9000 38.8000 ;
	    RECT 56.6000 34.7000 57.0000 35.1000 ;
	    RECT 57.4000 32.1000 57.8000 37.9000 ;
	    RECT 62.2000 36.8000 62.6000 37.2000 ;
	    RECT 62.2000 36.2000 62.5000 36.8000 ;
	    RECT 63.8000 36.2000 64.1000 42.8000 ;
	    RECT 59.0000 33.1000 59.4000 35.9000 ;
	    RECT 62.2000 35.8000 62.6000 36.2000 ;
	    RECT 63.8000 35.8000 64.2000 36.2000 ;
	    RECT 66.2000 35.8000 66.6000 36.2000 ;
	    RECT 63.0000 35.1000 63.4000 35.2000 ;
	    RECT 63.8000 35.1000 64.2000 35.2000 ;
	    RECT 63.0000 34.8000 64.2000 35.1000 ;
	    RECT 55.8000 27.8000 56.2000 28.2000 ;
	    RECT 54.2000 26.8000 54.6000 27.2000 ;
	    RECT 54.2000 26.2000 54.5000 26.8000 ;
	    RECT 51.8000 26.1000 52.2000 26.2000 ;
	    RECT 52.6000 26.1000 53.0000 26.2000 ;
	    RECT 51.8000 25.8000 53.0000 26.1000 ;
	    RECT 54.2000 25.8000 54.6000 26.2000 ;
	    RECT 55.8000 24.2000 56.1000 27.8000 ;
	    RECT 58.2000 25.1000 58.6000 27.9000 ;
	    RECT 55.8000 23.8000 56.2000 24.2000 ;
	    RECT 51.0000 22.1000 51.4000 22.2000 ;
	    RECT 51.8000 22.1000 52.2000 22.2000 ;
	    RECT 51.0000 21.8000 52.2000 22.1000 ;
	    RECT 53.4000 17.1000 53.8000 17.2000 ;
	    RECT 54.2000 17.1000 54.6000 17.2000 ;
	    RECT 53.4000 16.8000 54.6000 17.1000 ;
	    RECT 51.8000 15.9000 52.2000 16.3000 ;
	    RECT 55.1000 15.9000 55.5000 16.3000 ;
	    RECT 51.8000 14.2000 52.1000 15.9000 ;
	    RECT 53.8000 14.2000 54.2000 14.3000 ;
	    RECT 50.2000 13.8000 50.6000 14.2000 ;
	    RECT 51.8000 13.9000 54.2000 14.2000 ;
	    RECT 51.8000 13.5000 52.1000 13.9000 ;
	    RECT 52.5000 13.5000 52.9000 13.6000 ;
	    RECT 54.2000 13.5000 54.6000 13.6000 ;
	    RECT 55.2000 13.5000 55.5000 15.9000 ;
	    RECT 43.0000 12.8000 43.4000 13.2000 ;
	    RECT 46.2000 12.8000 46.6000 13.2000 ;
	    RECT 47.0000 12.8000 47.4000 13.2000 ;
	    RECT 48.6000 13.1000 49.0000 13.2000 ;
	    RECT 49.4000 13.1000 49.8000 13.2000 ;
	    RECT 48.6000 12.8000 49.8000 13.1000 ;
	    RECT 50.2000 12.8000 50.6000 13.2000 ;
	    RECT 51.8000 13.1000 52.2000 13.5000 ;
	    RECT 52.5000 13.2000 54.6000 13.5000 ;
	    RECT 55.1000 13.1000 55.5000 13.5000 ;
	    RECT 55.8000 14.2000 56.1000 23.8000 ;
	    RECT 59.8000 23.1000 60.2000 28.9000 ;
	    RECT 60.6000 26.8000 61.0000 27.2000 ;
	    RECT 60.6000 26.3000 60.9000 26.8000 ;
	    RECT 60.6000 25.9000 61.0000 26.3000 ;
	    RECT 63.8000 25.8000 64.2000 26.2000 ;
	    RECT 63.8000 23.2000 64.1000 25.8000 ;
	    RECT 63.8000 22.8000 64.2000 23.2000 ;
	    RECT 64.6000 23.1000 65.0000 28.9000 ;
	    RECT 66.2000 28.2000 66.5000 35.8000 ;
	    RECT 66.2000 27.8000 66.6000 28.2000 ;
	    RECT 67.0000 28.1000 67.3000 42.8000 ;
	    RECT 69.4000 39.2000 69.7000 44.8000 ;
	    RECT 69.4000 38.8000 69.8000 39.2000 ;
	    RECT 71.0000 36.2000 71.3000 55.8000 ;
	    RECT 71.8000 54.8000 72.2000 55.2000 ;
	    RECT 73.4000 55.1000 73.8000 55.2000 ;
	    RECT 74.2000 55.1000 74.6000 55.2000 ;
	    RECT 73.4000 54.8000 74.6000 55.1000 ;
	    RECT 75.0000 54.8000 75.4000 55.2000 ;
	    RECT 71.8000 51.2000 72.1000 54.8000 ;
	    RECT 72.6000 54.1000 73.0000 54.2000 ;
	    RECT 72.6000 53.8000 73.7000 54.1000 ;
	    RECT 71.8000 50.8000 72.2000 51.2000 ;
	    RECT 71.8000 48.2000 72.1000 50.8000 ;
	    RECT 73.4000 49.2000 73.7000 53.8000 ;
	    RECT 73.4000 48.8000 73.8000 49.2000 ;
	    RECT 71.8000 47.8000 72.2000 48.2000 ;
	    RECT 72.6000 47.8000 73.0000 48.2000 ;
	    RECT 72.6000 46.2000 72.9000 47.8000 ;
	    RECT 75.0000 47.2000 75.3000 54.8000 ;
	    RECT 75.8000 54.2000 76.1000 68.8000 ;
	    RECT 78.2000 65.8000 78.6000 66.2000 ;
	    RECT 78.2000 63.2000 78.5000 65.8000 ;
	    RECT 78.2000 62.8000 78.6000 63.2000 ;
	    RECT 79.0000 63.1000 79.4000 68.9000 ;
	    RECT 79.8000 66.8000 80.2000 67.2000 ;
	    RECT 79.8000 57.1000 80.1000 66.8000 ;
	    RECT 83.8000 66.2000 84.1000 70.8000 ;
	    RECT 86.2000 69.2000 86.5000 70.8000 ;
	    RECT 89.4000 69.8000 89.8000 70.2000 ;
	    RECT 84.6000 68.8000 85.0000 69.2000 ;
	    RECT 86.2000 68.8000 86.6000 69.2000 ;
	    RECT 84.6000 67.2000 84.9000 68.8000 ;
	    RECT 85.4000 67.8000 85.8000 68.2000 ;
	    RECT 85.4000 67.2000 85.7000 67.8000 ;
	    RECT 84.6000 66.8000 85.0000 67.2000 ;
	    RECT 85.4000 66.8000 85.8000 67.2000 ;
	    RECT 87.0000 66.8000 87.4000 67.2000 ;
	    RECT 82.2000 65.8000 82.6000 66.2000 ;
	    RECT 83.8000 65.8000 84.2000 66.2000 ;
	    RECT 82.2000 65.2000 82.5000 65.8000 ;
	    RECT 82.2000 64.8000 82.6000 65.2000 ;
	    RECT 83.8000 65.1000 84.2000 65.2000 ;
	    RECT 87.0000 65.1000 87.3000 66.8000 ;
	    RECT 89.4000 66.2000 89.7000 69.8000 ;
	    RECT 93.4000 68.2000 93.7000 74.8000 ;
	    RECT 97.4000 74.2000 97.7000 74.8000 ;
	    RECT 95.0000 73.8000 95.4000 74.2000 ;
	    RECT 95.8000 73.8000 96.2000 74.2000 ;
	    RECT 97.4000 73.8000 97.8000 74.2000 ;
	    RECT 94.2000 71.8000 94.6000 72.2000 ;
	    RECT 93.4000 67.8000 93.8000 68.2000 ;
	    RECT 90.2000 66.8000 90.6000 67.2000 ;
	    RECT 90.2000 66.2000 90.5000 66.8000 ;
	    RECT 94.2000 66.2000 94.5000 71.8000 ;
	    RECT 87.8000 66.1000 88.2000 66.2000 ;
	    RECT 88.6000 66.1000 89.0000 66.2000 ;
	    RECT 87.8000 65.8000 89.0000 66.1000 ;
	    RECT 89.4000 65.8000 89.8000 66.2000 ;
	    RECT 90.2000 65.8000 90.6000 66.2000 ;
	    RECT 94.2000 65.8000 94.6000 66.2000 ;
	    RECT 89.4000 65.2000 89.7000 65.8000 ;
	    RECT 83.8000 64.8000 87.3000 65.1000 ;
	    RECT 88.6000 64.8000 89.0000 65.2000 ;
	    RECT 89.4000 64.8000 89.8000 65.2000 ;
	    RECT 92.6000 64.8000 93.0000 65.2000 ;
	    RECT 88.6000 64.2000 88.9000 64.8000 ;
	    RECT 92.6000 64.2000 92.9000 64.8000 ;
	    RECT 81.4000 64.1000 81.8000 64.2000 ;
	    RECT 82.2000 64.1000 82.6000 64.2000 ;
	    RECT 81.4000 63.8000 82.6000 64.1000 ;
	    RECT 88.6000 63.8000 89.0000 64.2000 ;
	    RECT 90.2000 64.1000 90.6000 64.2000 ;
	    RECT 91.0000 64.1000 91.4000 64.2000 ;
	    RECT 90.2000 63.8000 91.4000 64.1000 ;
	    RECT 92.6000 63.8000 93.0000 64.2000 ;
	    RECT 84.6000 62.8000 85.0000 63.2000 ;
	    RECT 79.0000 56.8000 80.1000 57.1000 ;
	    RECT 80.6000 58.8000 81.0000 59.2000 ;
	    RECT 80.6000 57.2000 80.9000 58.8000 ;
	    RECT 84.6000 57.2000 84.9000 62.8000 ;
	    RECT 90.2000 59.2000 90.5000 63.8000 ;
	    RECT 95.0000 61.2000 95.3000 73.8000 ;
	    RECT 95.8000 73.2000 96.1000 73.8000 ;
	    RECT 95.8000 72.8000 96.2000 73.2000 ;
	    RECT 96.6000 73.1000 97.0000 73.2000 ;
	    RECT 97.4000 73.1000 97.8000 73.2000 ;
	    RECT 96.6000 72.8000 97.8000 73.1000 ;
	    RECT 98.2000 71.2000 98.5000 85.8000 ;
	    RECT 100.6000 85.2000 100.9000 89.8000 ;
	    RECT 102.2000 87.2000 102.5000 100.8000 ;
	    RECT 103.8000 98.2000 104.1000 101.8000 ;
	    RECT 103.8000 97.8000 104.2000 98.2000 ;
	    RECT 103.0000 92.8000 103.4000 93.2000 ;
	    RECT 103.8000 93.1000 104.2000 95.9000 ;
	    RECT 104.6000 93.8000 105.0000 94.2000 ;
	    RECT 103.0000 90.2000 103.3000 92.8000 ;
	    RECT 103.0000 89.8000 103.4000 90.2000 ;
	    RECT 104.6000 88.2000 104.9000 93.8000 ;
	    RECT 105.4000 92.1000 105.8000 97.9000 ;
	    RECT 106.2000 94.7000 106.6000 95.1000 ;
	    RECT 109.4000 94.8000 109.8000 95.2000 ;
	    RECT 106.2000 94.2000 106.5000 94.7000 ;
	    RECT 109.4000 94.2000 109.7000 94.8000 ;
	    RECT 106.2000 93.8000 106.6000 94.2000 ;
	    RECT 109.4000 93.8000 109.8000 94.2000 ;
	    RECT 110.2000 92.1000 110.6000 97.9000 ;
	    RECT 111.0000 94.8000 111.4000 95.2000 ;
	    RECT 105.4000 90.8000 105.8000 91.2000 ;
	    RECT 105.4000 89.2000 105.7000 90.8000 ;
	    RECT 111.0000 89.2000 111.3000 94.8000 ;
	    RECT 113.4000 94.1000 113.8000 94.2000 ;
	    RECT 114.2000 94.1000 114.6000 94.2000 ;
	    RECT 113.4000 93.8000 114.6000 94.1000 ;
	    RECT 115.0000 93.1000 115.4000 95.9000 ;
	    RECT 113.4000 91.8000 113.8000 92.2000 ;
	    RECT 116.6000 92.1000 117.0000 97.9000 ;
	    RECT 117.4000 94.7000 117.8000 95.1000 ;
	    RECT 117.4000 94.2000 117.7000 94.7000 ;
	    RECT 117.4000 93.8000 117.8000 94.2000 ;
	    RECT 105.4000 88.8000 105.8000 89.2000 ;
	    RECT 107.8000 88.8000 108.2000 89.2000 ;
	    RECT 111.0000 88.8000 111.4000 89.2000 ;
	    RECT 104.6000 87.8000 105.0000 88.2000 ;
	    RECT 107.8000 87.2000 108.1000 88.8000 ;
	    RECT 108.6000 87.8000 109.0000 88.2000 ;
	    RECT 108.6000 87.2000 108.9000 87.8000 ;
	    RECT 101.4000 87.1000 101.8000 87.2000 ;
	    RECT 102.2000 87.1000 102.6000 87.2000 ;
	    RECT 101.4000 86.8000 102.6000 87.1000 ;
	    RECT 107.8000 86.8000 108.2000 87.2000 ;
	    RECT 108.6000 86.8000 109.0000 87.2000 ;
	    RECT 111.8000 86.8000 112.2000 87.2000 ;
	    RECT 112.6000 86.8000 113.0000 87.2000 ;
	    RECT 111.8000 86.2000 112.1000 86.8000 ;
	    RECT 112.6000 86.2000 112.9000 86.8000 ;
	    RECT 113.4000 86.2000 113.7000 91.8000 ;
	    RECT 118.2000 89.2000 118.5000 101.8000 ;
	    RECT 120.6000 94.8000 121.0000 95.2000 ;
	    RECT 120.6000 94.2000 120.9000 94.8000 ;
	    RECT 120.6000 93.8000 121.0000 94.2000 ;
	    RECT 121.4000 92.1000 121.8000 97.9000 ;
	    RECT 122.2000 96.2000 122.5000 105.8000 ;
	    RECT 124.6000 103.2000 124.9000 106.8000 ;
	    RECT 124.6000 102.8000 125.0000 103.2000 ;
	    RECT 126.2000 103.1000 126.6000 108.9000 ;
	    RECT 127.0000 107.2000 127.3000 126.8000 ;
	    RECT 128.6000 125.8000 129.0000 126.2000 ;
	    RECT 128.6000 125.2000 128.9000 125.8000 ;
	    RECT 128.6000 124.8000 129.0000 125.2000 ;
	    RECT 129.4000 125.1000 129.8000 127.9000 ;
	    RECT 130.2000 127.8000 130.6000 128.2000 ;
	    RECT 130.2000 127.2000 130.5000 127.8000 ;
	    RECT 130.2000 126.8000 130.6000 127.2000 ;
	    RECT 128.6000 122.8000 129.0000 123.2000 ;
	    RECT 131.0000 123.1000 131.4000 128.9000 ;
	    RECT 128.6000 117.2000 128.9000 122.8000 ;
	    RECT 132.6000 120.2000 132.9000 141.8000 ;
	    RECT 135.8000 140.2000 136.1000 141.8000 ;
	    RECT 135.8000 139.8000 136.2000 140.2000 ;
	    RECT 143.8000 139.8000 144.2000 140.2000 ;
	    RECT 137.4000 139.1000 137.8000 139.2000 ;
	    RECT 138.2000 139.1000 138.6000 139.2000 ;
	    RECT 137.4000 138.8000 138.6000 139.1000 ;
	    RECT 134.2000 134.8000 134.6000 135.2000 ;
	    RECT 135.0000 134.8000 135.4000 135.2000 ;
	    RECT 134.2000 132.2000 134.5000 134.8000 ;
	    RECT 135.0000 133.2000 135.3000 134.8000 ;
	    RECT 135.0000 132.8000 135.4000 133.2000 ;
	    RECT 134.2000 131.8000 134.6000 132.2000 ;
	    RECT 135.0000 127.2000 135.3000 132.8000 ;
	    RECT 135.8000 132.1000 136.2000 137.9000 ;
	    RECT 137.4000 133.1000 137.8000 135.9000 ;
	    RECT 140.6000 132.1000 141.0000 137.9000 ;
	    RECT 143.8000 135.2000 144.1000 139.8000 ;
	    RECT 141.4000 135.1000 141.8000 135.2000 ;
	    RECT 142.2000 135.1000 142.6000 135.2000 ;
	    RECT 141.4000 134.8000 142.6000 135.1000 ;
	    RECT 143.8000 134.8000 144.2000 135.2000 ;
	    RECT 145.4000 132.1000 145.8000 137.9000 ;
	    RECT 151.8000 137.2000 152.1000 145.8000 ;
	    RECT 155.0000 143.1000 155.4000 148.9000 ;
	    RECT 158.2000 148.8000 158.6000 149.2000 ;
	    RECT 156.6000 145.1000 157.0000 147.9000 ;
	    RECT 159.8000 145.8000 160.2000 146.2000 ;
	    RECT 159.8000 145.2000 160.1000 145.8000 ;
	    RECT 159.8000 144.8000 160.2000 145.2000 ;
	    RECT 162.2000 145.1000 162.6000 147.9000 ;
	    RECT 159.8000 142.2000 160.1000 144.8000 ;
	    RECT 163.8000 143.1000 164.2000 148.9000 ;
	    RECT 167.0000 146.2000 167.3000 153.8000 ;
	    RECT 167.8000 153.1000 168.2000 155.9000 ;
	    RECT 171.8000 155.8000 173.0000 156.1000 ;
	    RECT 179.8000 155.8000 180.2000 156.2000 ;
	    RECT 181.4000 156.1000 181.8000 156.2000 ;
	    RECT 182.2000 156.1000 182.6000 156.2000 ;
	    RECT 181.4000 155.8000 182.6000 156.1000 ;
	    RECT 168.6000 154.8000 169.0000 155.2000 ;
	    RECT 173.4000 154.8000 173.8000 155.2000 ;
	    RECT 175.0000 154.8000 175.4000 155.2000 ;
	    RECT 168.6000 154.2000 168.9000 154.8000 ;
	    RECT 168.6000 153.8000 169.0000 154.2000 ;
	    RECT 170.2000 154.1000 170.6000 154.2000 ;
	    RECT 171.0000 154.1000 171.4000 154.2000 ;
	    RECT 170.2000 153.8000 171.4000 154.1000 ;
	    RECT 168.6000 153.1000 169.0000 153.2000 ;
	    RECT 169.4000 153.1000 169.8000 153.2000 ;
	    RECT 168.6000 152.8000 169.8000 153.1000 ;
	    RECT 173.4000 152.2000 173.7000 154.8000 ;
	    RECT 175.0000 154.2000 175.3000 154.8000 ;
	    RECT 179.8000 154.2000 180.1000 155.8000 ;
	    RECT 175.0000 153.8000 175.4000 154.2000 ;
	    RECT 176.6000 154.1000 177.0000 154.2000 ;
	    RECT 177.4000 154.1000 177.8000 154.2000 ;
	    RECT 176.6000 153.8000 177.8000 154.1000 ;
	    RECT 178.2000 154.1000 178.6000 154.2000 ;
	    RECT 179.0000 154.1000 179.4000 154.2000 ;
	    RECT 178.2000 153.8000 179.4000 154.1000 ;
	    RECT 179.8000 153.8000 180.2000 154.2000 ;
	    RECT 173.4000 151.8000 173.8000 152.2000 ;
	    RECT 175.0000 151.2000 175.3000 153.8000 ;
	    RECT 176.6000 152.8000 177.0000 153.2000 ;
	    RECT 176.6000 152.2000 176.9000 152.8000 ;
	    RECT 179.8000 152.2000 180.1000 153.8000 ;
	    RECT 176.6000 151.8000 177.0000 152.2000 ;
	    RECT 179.8000 151.8000 180.2000 152.2000 ;
	    RECT 180.6000 151.8000 181.0000 152.2000 ;
	    RECT 175.0000 150.8000 175.4000 151.2000 ;
	    RECT 165.4000 146.1000 165.8000 146.2000 ;
	    RECT 166.2000 146.1000 166.6000 146.2000 ;
	    RECT 165.4000 145.8000 166.6000 146.1000 ;
	    RECT 167.0000 145.8000 167.4000 146.2000 ;
	    RECT 159.8000 141.8000 160.2000 142.2000 ;
	    RECT 163.8000 141.8000 164.2000 142.2000 ;
	    RECT 151.8000 136.8000 152.2000 137.2000 ;
	    RECT 147.0000 133.1000 147.4000 135.9000 ;
	    RECT 150.2000 131.8000 150.6000 132.2000 ;
	    RECT 152.6000 132.1000 153.0000 137.9000 ;
	    RECT 156.6000 134.7000 157.0000 135.1000 ;
	    RECT 156.6000 132.2000 156.9000 134.7000 ;
	    RECT 156.6000 131.8000 157.0000 132.2000 ;
	    RECT 157.4000 132.1000 157.8000 137.9000 ;
	    RECT 158.2000 134.8000 158.6000 135.2000 ;
	    RECT 158.2000 134.2000 158.5000 134.8000 ;
	    RECT 158.2000 133.8000 158.6000 134.2000 ;
	    RECT 159.0000 133.1000 159.4000 135.9000 ;
	    RECT 159.0000 131.8000 159.4000 132.2000 ;
	    RECT 133.4000 126.8000 133.8000 127.2000 ;
	    RECT 135.0000 126.8000 135.4000 127.2000 ;
	    RECT 133.4000 126.2000 133.7000 126.8000 ;
	    RECT 133.4000 125.8000 133.8000 126.2000 ;
	    RECT 135.8000 123.1000 136.2000 128.9000 ;
	    RECT 150.2000 128.2000 150.5000 131.8000 ;
	    RECT 159.0000 129.2000 159.3000 131.8000 ;
	    RECT 163.8000 129.2000 164.1000 141.8000 ;
	    RECT 167.0000 139.2000 167.3000 145.8000 ;
	    RECT 168.6000 143.1000 169.0000 148.9000 ;
	    RECT 171.0000 148.8000 171.4000 149.2000 ;
	    RECT 171.0000 148.2000 171.3000 148.8000 ;
	    RECT 171.0000 147.8000 171.4000 148.2000 ;
	    RECT 171.8000 148.1000 172.2000 148.2000 ;
	    RECT 172.6000 148.1000 173.0000 148.2000 ;
	    RECT 171.8000 147.8000 173.0000 148.1000 ;
	    RECT 173.4000 146.8000 173.8000 147.2000 ;
	    RECT 173.4000 146.2000 173.7000 146.8000 ;
	    RECT 173.4000 145.8000 173.8000 146.2000 ;
	    RECT 175.8000 144.8000 176.2000 145.2000 ;
	    RECT 175.8000 142.2000 176.1000 144.8000 ;
	    RECT 175.8000 141.8000 176.2000 142.2000 ;
	    RECT 175.8000 139.2000 176.1000 141.8000 ;
	    RECT 176.6000 140.2000 176.9000 151.8000 ;
	    RECT 178.2000 150.8000 178.6000 151.2000 ;
	    RECT 178.2000 147.2000 178.5000 150.8000 ;
	    RECT 180.6000 149.2000 180.9000 151.8000 ;
	    RECT 181.4000 150.2000 181.7000 155.8000 ;
	    RECT 182.2000 152.8000 182.6000 153.2000 ;
	    RECT 182.2000 152.2000 182.5000 152.8000 ;
	    RECT 182.2000 151.8000 182.6000 152.2000 ;
	    RECT 181.4000 149.8000 181.8000 150.2000 ;
	    RECT 180.6000 148.8000 181.0000 149.2000 ;
	    RECT 180.6000 147.8000 181.0000 148.2000 ;
	    RECT 178.2000 146.8000 178.6000 147.2000 ;
	    RECT 179.0000 146.8000 179.4000 147.2000 ;
	    RECT 180.6000 147.0000 180.9000 147.8000 ;
	    RECT 181.4000 147.2000 181.7000 149.8000 ;
	    RECT 182.2000 148.8000 182.6000 149.2000 ;
	    RECT 182.2000 148.2000 182.5000 148.8000 ;
	    RECT 182.2000 147.8000 182.6000 148.2000 ;
	    RECT 177.4000 145.8000 177.8000 146.2000 ;
	    RECT 177.4000 144.2000 177.7000 145.8000 ;
	    RECT 177.4000 143.8000 177.8000 144.2000 ;
	    RECT 176.6000 139.8000 177.0000 140.2000 ;
	    RECT 178.2000 139.2000 178.5000 146.8000 ;
	    RECT 179.0000 146.2000 179.3000 146.8000 ;
	    RECT 180.6000 146.6000 181.0000 147.0000 ;
	    RECT 181.4000 146.8000 181.8000 147.2000 ;
	    RECT 183.0000 146.2000 183.3000 174.8000 ;
	    RECT 183.8000 173.8000 184.2000 174.2000 ;
	    RECT 185.4000 173.8000 185.8000 174.2000 ;
	    RECT 183.8000 173.2000 184.1000 173.8000 ;
	    RECT 183.8000 172.8000 184.2000 173.2000 ;
	    RECT 185.4000 168.2000 185.7000 173.8000 ;
	    RECT 187.0000 173.2000 187.3000 174.8000 ;
	    RECT 187.0000 172.8000 187.4000 173.2000 ;
	    RECT 190.2000 173.1000 190.6000 175.9000 ;
	    RECT 191.0000 173.8000 191.4000 174.2000 ;
	    RECT 191.0000 172.2000 191.3000 173.8000 ;
	    RECT 191.0000 171.8000 191.4000 172.2000 ;
	    RECT 191.8000 172.1000 192.2000 177.9000 ;
	    RECT 193.4000 174.8000 193.8000 175.2000 ;
	    RECT 185.4000 167.8000 185.8000 168.2000 ;
	    RECT 183.8000 166.8000 184.2000 167.2000 ;
	    RECT 183.8000 166.2000 184.1000 166.8000 ;
	    RECT 183.8000 165.8000 184.2000 166.2000 ;
	    RECT 184.6000 164.8000 185.0000 165.2000 ;
	    RECT 184.6000 159.2000 184.9000 164.8000 ;
	    RECT 187.8000 163.8000 188.2000 164.2000 ;
	    RECT 184.6000 158.8000 185.0000 159.2000 ;
	    RECT 187.8000 156.2000 188.1000 163.8000 ;
	    RECT 188.6000 163.1000 189.0000 168.9000 ;
	    RECT 191.0000 167.2000 191.3000 171.8000 ;
	    RECT 193.4000 170.2000 193.7000 174.8000 ;
	    RECT 196.6000 172.1000 197.0000 177.9000 ;
	    RECT 202.2000 177.8000 202.6000 178.2000 ;
	    RECT 215.0000 178.1000 215.4000 178.2000 ;
	    RECT 215.8000 178.1000 216.2000 178.2000 ;
	    RECT 202.2000 176.2000 202.5000 177.8000 ;
	    RECT 205.4000 176.8000 205.8000 177.2000 ;
	    RECT 205.4000 176.2000 205.7000 176.8000 ;
	    RECT 202.2000 175.8000 202.6000 176.2000 ;
	    RECT 205.4000 175.8000 205.8000 176.2000 ;
	    RECT 200.6000 174.8000 201.0000 175.2000 ;
	    RECT 200.6000 174.2000 200.9000 174.8000 ;
	    RECT 199.0000 174.1000 199.4000 174.2000 ;
	    RECT 199.8000 174.1000 200.2000 174.2000 ;
	    RECT 199.0000 173.8000 200.2000 174.1000 ;
	    RECT 200.6000 173.8000 201.0000 174.2000 ;
	    RECT 203.8000 173.8000 204.2000 174.2000 ;
	    RECT 203.8000 172.2000 204.1000 173.8000 ;
	    RECT 205.4000 172.8000 205.8000 173.2000 ;
	    RECT 206.2000 173.1000 206.6000 175.9000 ;
	    RECT 207.0000 173.8000 207.4000 174.2000 ;
	    RECT 199.0000 171.8000 199.4000 172.2000 ;
	    RECT 203.8000 171.8000 204.2000 172.2000 ;
	    RECT 193.4000 169.8000 193.8000 170.2000 ;
	    RECT 191.0000 166.8000 191.4000 167.2000 ;
	    RECT 191.0000 166.1000 191.4000 166.2000 ;
	    RECT 191.8000 166.1000 192.2000 166.2000 ;
	    RECT 191.0000 165.8000 192.2000 166.1000 ;
	    RECT 193.4000 163.1000 193.8000 168.9000 ;
	    RECT 195.0000 165.1000 195.4000 167.9000 ;
	    RECT 195.8000 165.1000 196.2000 167.9000 ;
	    RECT 197.4000 163.1000 197.8000 168.9000 ;
	    RECT 198.2000 165.9000 198.6000 166.3000 ;
	    RECT 198.2000 165.2000 198.5000 165.9000 ;
	    RECT 199.0000 165.2000 199.3000 171.8000 ;
	    RECT 203.0000 170.8000 203.4000 171.2000 ;
	    RECT 198.2000 164.8000 198.6000 165.2000 ;
	    RECT 199.0000 164.8000 199.4000 165.2000 ;
	    RECT 202.2000 163.1000 202.6000 168.9000 ;
	    RECT 203.0000 164.2000 203.3000 170.8000 ;
	    RECT 205.4000 168.2000 205.7000 172.8000 ;
	    RECT 207.0000 171.2000 207.3000 173.8000 ;
	    RECT 207.8000 172.1000 208.2000 177.9000 ;
	    RECT 208.6000 175.8000 209.0000 176.2000 ;
	    RECT 208.6000 175.1000 208.9000 175.8000 ;
	    RECT 208.6000 174.7000 209.0000 175.1000 ;
	    RECT 212.6000 172.1000 213.0000 177.9000 ;
	    RECT 215.0000 177.8000 216.2000 178.1000 ;
	    RECT 222.2000 176.8000 222.6000 177.2000 ;
	    RECT 222.2000 176.2000 222.5000 176.8000 ;
	    RECT 222.2000 175.8000 222.6000 176.2000 ;
	    RECT 223.0000 175.8000 223.4000 176.2000 ;
	    RECT 223.0000 175.2000 223.3000 175.8000 ;
	    RECT 217.4000 174.8000 217.8000 175.2000 ;
	    RECT 219.0000 175.1000 219.4000 175.2000 ;
	    RECT 219.8000 175.1000 220.2000 175.2000 ;
	    RECT 219.0000 174.8000 220.2000 175.1000 ;
	    RECT 220.6000 174.8000 221.0000 175.2000 ;
	    RECT 222.2000 174.8000 222.6000 175.2000 ;
	    RECT 223.0000 174.8000 223.4000 175.2000 ;
	    RECT 224.6000 175.1000 225.0000 175.2000 ;
	    RECT 225.4000 175.1000 225.8000 175.2000 ;
	    RECT 224.6000 174.8000 225.8000 175.1000 ;
	    RECT 227.8000 174.8000 228.2000 175.2000 ;
	    RECT 217.4000 174.2000 217.7000 174.8000 ;
	    RECT 217.4000 173.8000 217.8000 174.2000 ;
	    RECT 219.0000 174.1000 219.4000 174.2000 ;
	    RECT 219.8000 174.1000 220.2000 174.2000 ;
	    RECT 219.0000 173.8000 220.2000 174.1000 ;
	    RECT 207.0000 170.8000 207.4000 171.2000 ;
	    RECT 206.2000 169.8000 206.6000 170.2000 ;
	    RECT 206.2000 169.2000 206.5000 169.8000 ;
	    RECT 206.2000 168.8000 206.6000 169.2000 ;
	    RECT 207.0000 168.2000 207.3000 170.8000 ;
	    RECT 214.2000 169.8000 214.6000 170.2000 ;
	    RECT 208.6000 168.8000 209.0000 169.2000 ;
	    RECT 208.6000 168.2000 208.9000 168.8000 ;
	    RECT 205.4000 167.8000 205.8000 168.2000 ;
	    RECT 207.0000 167.8000 207.4000 168.2000 ;
	    RECT 208.6000 167.8000 209.0000 168.2000 ;
	    RECT 210.2000 168.1000 210.6000 168.2000 ;
	    RECT 209.4000 167.8000 210.6000 168.1000 ;
	    RECT 203.0000 163.8000 203.4000 164.2000 ;
	    RECT 203.8000 164.1000 204.2000 164.2000 ;
	    RECT 204.6000 164.1000 205.0000 164.2000 ;
	    RECT 203.8000 163.8000 205.0000 164.1000 ;
	    RECT 193.4000 160.8000 193.8000 161.2000 ;
	    RECT 191.0000 157.1000 191.4000 157.2000 ;
	    RECT 191.8000 157.1000 192.2000 157.2000 ;
	    RECT 191.0000 156.8000 192.2000 157.1000 ;
	    RECT 183.8000 155.8000 184.2000 156.2000 ;
	    RECT 187.8000 155.8000 188.2000 156.2000 ;
	    RECT 183.8000 155.2000 184.1000 155.8000 ;
	    RECT 193.4000 155.2000 193.7000 160.8000 ;
	    RECT 195.8000 157.8000 196.2000 158.2000 ;
	    RECT 195.8000 156.2000 196.1000 157.8000 ;
	    RECT 199.8000 156.8000 200.2000 157.2000 ;
	    RECT 199.8000 156.2000 200.1000 156.8000 ;
	    RECT 195.8000 155.8000 196.2000 156.2000 ;
	    RECT 199.8000 155.8000 200.2000 156.2000 ;
	    RECT 183.8000 154.8000 184.2000 155.2000 ;
	    RECT 189.4000 154.8000 189.8000 155.2000 ;
	    RECT 191.8000 155.1000 192.2000 155.2000 ;
	    RECT 192.6000 155.1000 193.0000 155.2000 ;
	    RECT 191.8000 154.8000 193.0000 155.1000 ;
	    RECT 193.4000 154.8000 193.8000 155.2000 ;
	    RECT 199.0000 155.1000 199.4000 155.2000 ;
	    RECT 199.8000 155.1000 200.2000 155.2000 ;
	    RECT 199.0000 154.8000 200.2000 155.1000 ;
	    RECT 187.0000 153.8000 187.4000 154.2000 ;
	    RECT 183.8000 152.8000 184.2000 153.2000 ;
	    RECT 184.6000 152.8000 185.0000 153.2000 ;
	    RECT 183.8000 149.2000 184.1000 152.8000 ;
	    RECT 183.8000 148.8000 184.2000 149.2000 ;
	    RECT 179.0000 145.8000 179.4000 146.2000 ;
	    RECT 181.4000 145.8000 181.8000 146.2000 ;
	    RECT 183.0000 145.8000 183.4000 146.2000 ;
	    RECT 179.0000 144.8000 179.4000 145.2000 ;
	    RECT 167.0000 138.8000 167.4000 139.2000 ;
	    RECT 175.8000 138.8000 176.2000 139.2000 ;
	    RECT 178.2000 138.8000 178.6000 139.2000 ;
	    RECT 177.4000 137.1000 177.8000 137.2000 ;
	    RECT 178.2000 137.1000 178.6000 137.2000 ;
	    RECT 177.4000 136.8000 178.6000 137.1000 ;
	    RECT 169.4000 135.8000 169.8000 136.2000 ;
	    RECT 175.8000 136.1000 176.2000 136.2000 ;
	    RECT 176.6000 136.1000 177.0000 136.2000 ;
	    RECT 175.8000 135.8000 177.0000 136.1000 ;
	    RECT 166.2000 132.8000 166.6000 133.2000 ;
	    RECT 159.0000 128.8000 159.4000 129.2000 ;
	    RECT 163.8000 128.8000 164.2000 129.2000 ;
	    RECT 147.0000 128.1000 147.4000 128.2000 ;
	    RECT 147.8000 128.1000 148.2000 128.2000 ;
	    RECT 147.0000 127.8000 148.2000 128.1000 ;
	    RECT 150.2000 127.8000 150.6000 128.2000 ;
	    RECT 152.6000 127.8000 153.0000 128.2000 ;
	    RECT 153.4000 128.1000 153.8000 128.2000 ;
	    RECT 154.2000 128.1000 154.6000 128.2000 ;
	    RECT 153.4000 127.8000 154.6000 128.1000 ;
	    RECT 158.2000 127.8000 158.6000 128.2000 ;
	    RECT 159.0000 128.1000 159.4000 128.2000 ;
	    RECT 159.8000 128.1000 160.2000 128.2000 ;
	    RECT 159.0000 127.8000 160.2000 128.1000 ;
	    RECT 152.6000 127.2000 152.9000 127.8000 ;
	    RECT 139.8000 126.8000 140.2000 127.2000 ;
	    RECT 140.6000 127.1000 141.0000 127.2000 ;
	    RECT 141.4000 127.1000 141.8000 127.2000 ;
	    RECT 140.6000 126.8000 141.8000 127.1000 ;
	    RECT 144.6000 126.8000 145.0000 127.2000 ;
	    RECT 145.4000 126.8000 145.8000 127.2000 ;
	    RECT 146.2000 127.1000 146.6000 127.2000 ;
	    RECT 147.0000 127.1000 147.4000 127.2000 ;
	    RECT 146.2000 126.8000 147.4000 127.1000 ;
	    RECT 148.6000 126.8000 149.0000 127.2000 ;
	    RECT 152.6000 126.8000 153.0000 127.2000 ;
	    RECT 138.2000 126.1000 138.6000 126.2000 ;
	    RECT 139.0000 126.1000 139.4000 126.2000 ;
	    RECT 138.2000 125.8000 139.4000 126.1000 ;
	    RECT 138.2000 124.2000 138.5000 125.8000 ;
	    RECT 139.0000 124.8000 139.4000 125.2000 ;
	    RECT 138.2000 123.8000 138.6000 124.2000 ;
	    RECT 132.6000 119.8000 133.0000 120.2000 ;
	    RECT 128.6000 116.8000 129.0000 117.2000 ;
	    RECT 129.4000 117.1000 129.8000 117.2000 ;
	    RECT 130.2000 117.1000 130.6000 117.2000 ;
	    RECT 129.4000 116.8000 130.6000 117.1000 ;
	    RECT 131.0000 117.1000 131.4000 117.2000 ;
	    RECT 131.8000 117.1000 132.2000 117.2000 ;
	    RECT 131.0000 116.8000 132.2000 117.1000 ;
	    RECT 134.2000 116.8000 134.6000 117.2000 ;
	    RECT 128.6000 115.2000 128.9000 116.8000 ;
	    RECT 134.2000 116.2000 134.5000 116.8000 ;
	    RECT 139.0000 116.2000 139.3000 124.8000 ;
	    RECT 139.8000 123.2000 140.1000 126.8000 ;
	    RECT 142.2000 124.8000 142.6000 125.2000 ;
	    RECT 142.2000 124.2000 142.5000 124.8000 ;
	    RECT 142.2000 123.8000 142.6000 124.2000 ;
	    RECT 144.6000 123.2000 144.9000 126.8000 ;
	    RECT 145.4000 126.2000 145.7000 126.8000 ;
	    RECT 145.4000 125.8000 145.8000 126.2000 ;
	    RECT 147.0000 126.1000 147.4000 126.2000 ;
	    RECT 147.8000 126.1000 148.2000 126.2000 ;
	    RECT 147.0000 125.8000 148.2000 126.1000 ;
	    RECT 148.6000 123.2000 148.9000 126.8000 ;
	    RECT 154.2000 126.2000 154.5000 127.8000 ;
	    RECT 158.2000 127.2000 158.5000 127.8000 ;
	    RECT 155.0000 126.8000 155.4000 127.2000 ;
	    RECT 158.2000 126.8000 158.6000 127.2000 ;
	    RECT 151.0000 125.8000 151.4000 126.2000 ;
	    RECT 152.6000 125.8000 153.0000 126.2000 ;
	    RECT 154.2000 125.8000 154.6000 126.2000 ;
	    RECT 151.0000 125.2000 151.3000 125.8000 ;
	    RECT 152.6000 125.2000 152.9000 125.8000 ;
	    RECT 151.0000 124.8000 151.4000 125.2000 ;
	    RECT 152.6000 124.8000 153.0000 125.2000 ;
	    RECT 139.8000 122.8000 140.2000 123.2000 ;
	    RECT 144.6000 122.8000 145.0000 123.2000 ;
	    RECT 148.6000 122.8000 149.0000 123.2000 ;
	    RECT 141.4000 119.8000 141.8000 120.2000 ;
	    RECT 144.6000 119.8000 145.0000 120.2000 ;
	    RECT 132.6000 115.8000 133.0000 116.2000 ;
	    RECT 134.2000 115.8000 134.6000 116.2000 ;
	    RECT 135.8000 115.8000 136.2000 116.2000 ;
	    RECT 139.0000 115.8000 139.4000 116.2000 ;
	    RECT 128.6000 114.8000 129.0000 115.2000 ;
	    RECT 130.2000 114.8000 130.6000 115.2000 ;
	    RECT 130.2000 114.2000 130.5000 114.8000 ;
	    RECT 130.2000 113.8000 130.6000 114.2000 ;
	    RECT 131.8000 113.8000 132.2000 114.2000 ;
	    RECT 131.8000 113.2000 132.1000 113.8000 ;
	    RECT 132.6000 113.2000 132.9000 115.8000 ;
	    RECT 135.8000 115.2000 136.1000 115.8000 ;
	    RECT 134.2000 115.1000 134.6000 115.2000 ;
	    RECT 135.0000 115.1000 135.4000 115.2000 ;
	    RECT 134.2000 114.8000 135.4000 115.1000 ;
	    RECT 135.8000 114.8000 136.2000 115.2000 ;
	    RECT 140.6000 114.8000 141.0000 115.2000 ;
	    RECT 134.2000 114.2000 134.5000 114.8000 ;
	    RECT 140.6000 114.2000 140.9000 114.8000 ;
	    RECT 141.4000 114.2000 141.7000 119.8000 ;
	    RECT 144.6000 115.2000 144.9000 119.8000 ;
	    RECT 144.6000 114.8000 145.0000 115.2000 ;
	    RECT 148.6000 114.2000 148.9000 122.8000 ;
	    RECT 153.4000 121.8000 153.8000 122.2000 ;
	    RECT 152.6000 117.8000 153.0000 118.2000 ;
	    RECT 151.8000 116.8000 152.2000 117.2000 ;
	    RECT 151.8000 116.2000 152.1000 116.8000 ;
	    RECT 149.4000 115.8000 149.8000 116.2000 ;
	    RECT 150.2000 115.8000 150.6000 116.2000 ;
	    RECT 151.8000 115.8000 152.2000 116.2000 ;
	    RECT 149.4000 115.2000 149.7000 115.8000 ;
	    RECT 150.2000 115.2000 150.5000 115.8000 ;
	    RECT 149.4000 114.8000 149.8000 115.2000 ;
	    RECT 150.2000 114.8000 150.6000 115.2000 ;
	    RECT 152.6000 114.2000 152.9000 117.8000 ;
	    RECT 153.4000 116.2000 153.7000 121.8000 ;
	    RECT 155.0000 118.2000 155.3000 126.8000 ;
	    RECT 158.2000 125.8000 158.6000 126.2000 ;
	    RECT 158.2000 125.2000 158.5000 125.8000 ;
	    RECT 157.4000 125.1000 157.8000 125.2000 ;
	    RECT 156.6000 124.8000 157.8000 125.1000 ;
	    RECT 158.2000 124.8000 158.6000 125.2000 ;
	    RECT 165.4000 125.1000 165.8000 127.9000 ;
	    RECT 156.6000 124.2000 156.9000 124.8000 ;
	    RECT 156.6000 123.8000 157.0000 124.2000 ;
	    RECT 156.6000 119.2000 156.9000 123.8000 ;
	    RECT 156.6000 118.8000 157.0000 119.2000 ;
	    RECT 159.8000 118.8000 160.2000 119.2000 ;
	    RECT 155.0000 117.8000 155.4000 118.2000 ;
	    RECT 153.4000 115.8000 153.8000 116.2000 ;
	    RECT 134.2000 113.8000 134.6000 114.2000 ;
	    RECT 135.0000 114.1000 135.4000 114.2000 ;
	    RECT 135.8000 114.1000 136.2000 114.2000 ;
	    RECT 135.0000 113.8000 136.2000 114.1000 ;
	    RECT 136.6000 113.8000 137.0000 114.2000 ;
	    RECT 139.8000 113.8000 140.2000 114.2000 ;
	    RECT 140.6000 113.8000 141.0000 114.2000 ;
	    RECT 141.4000 113.8000 141.8000 114.2000 ;
	    RECT 143.8000 114.1000 144.2000 114.2000 ;
	    RECT 144.6000 114.1000 145.0000 114.2000 ;
	    RECT 143.8000 113.8000 145.0000 114.1000 ;
	    RECT 147.0000 113.8000 147.4000 114.2000 ;
	    RECT 148.6000 113.8000 149.0000 114.2000 ;
	    RECT 149.4000 113.8000 149.8000 114.2000 ;
	    RECT 150.2000 113.8000 150.6000 114.2000 ;
	    RECT 152.6000 113.8000 153.0000 114.2000 ;
	    RECT 136.6000 113.2000 136.9000 113.8000 ;
	    RECT 139.8000 113.2000 140.1000 113.8000 ;
	    RECT 147.0000 113.2000 147.3000 113.8000 ;
	    RECT 131.8000 112.8000 132.2000 113.2000 ;
	    RECT 132.6000 112.8000 133.0000 113.2000 ;
	    RECT 136.6000 112.8000 137.0000 113.2000 ;
	    RECT 138.2000 112.8000 138.6000 113.2000 ;
	    RECT 139.8000 112.8000 140.2000 113.2000 ;
	    RECT 141.4000 113.1000 141.8000 113.2000 ;
	    RECT 142.2000 113.1000 142.6000 113.2000 ;
	    RECT 141.4000 112.8000 142.6000 113.1000 ;
	    RECT 146.2000 112.8000 146.6000 113.2000 ;
	    RECT 147.0000 112.8000 147.4000 113.2000 ;
	    RECT 137.4000 111.8000 137.8000 112.2000 ;
	    RECT 133.4000 109.1000 133.8000 109.2000 ;
	    RECT 134.2000 109.1000 134.6000 109.2000 ;
	    RECT 130.2000 107.8000 130.6000 108.2000 ;
	    RECT 127.0000 106.8000 127.4000 107.2000 ;
	    RECT 129.4000 106.8000 129.8000 107.2000 ;
	    RECT 129.4000 106.2000 129.7000 106.8000 ;
	    RECT 130.2000 106.3000 130.5000 107.8000 ;
	    RECT 129.4000 105.8000 129.8000 106.2000 ;
	    RECT 130.2000 105.9000 130.6000 106.3000 ;
	    RECT 127.8000 103.8000 128.2000 104.2000 ;
	    RECT 124.6000 99.2000 124.9000 102.8000 ;
	    RECT 127.8000 99.2000 128.1000 103.8000 ;
	    RECT 124.6000 98.8000 125.0000 99.2000 ;
	    RECT 127.8000 98.8000 128.2000 99.2000 ;
	    RECT 129.4000 97.2000 129.7000 105.8000 ;
	    RECT 131.0000 103.1000 131.4000 108.9000 ;
	    RECT 133.4000 108.8000 134.6000 109.1000 ;
	    RECT 132.6000 105.1000 133.0000 107.9000 ;
	    RECT 135.8000 103.1000 136.2000 108.9000 ;
	    RECT 137.4000 108.2000 137.7000 111.8000 ;
	    RECT 137.4000 107.8000 137.8000 108.2000 ;
	    RECT 136.6000 106.8000 137.0000 107.2000 ;
	    RECT 136.6000 106.2000 136.9000 106.8000 ;
	    RECT 136.6000 105.8000 137.0000 106.2000 ;
	    RECT 138.2000 105.1000 138.5000 112.8000 ;
	    RECT 143.0000 111.8000 143.4000 112.2000 ;
	    RECT 144.6000 111.8000 145.0000 112.2000 ;
	    RECT 143.0000 110.2000 143.3000 111.8000 ;
	    RECT 143.0000 109.8000 143.4000 110.2000 ;
	    RECT 139.0000 106.2000 139.4000 106.3000 ;
	    RECT 139.8000 106.2000 140.2000 106.3000 ;
	    RECT 139.0000 105.9000 140.2000 106.2000 ;
	    RECT 138.2000 104.8000 139.3000 105.1000 ;
	    RECT 129.4000 96.8000 129.8000 97.2000 ;
	    RECT 122.2000 95.8000 122.6000 96.2000 ;
	    RECT 124.6000 94.8000 125.0000 95.2000 ;
	    RECT 123.8000 91.8000 124.2000 92.2000 ;
	    RECT 120.6000 89.8000 121.0000 90.2000 ;
	    RECT 120.6000 89.2000 120.9000 89.8000 ;
	    RECT 114.2000 88.8000 114.6000 89.2000 ;
	    RECT 118.2000 88.8000 118.6000 89.2000 ;
	    RECT 120.6000 88.8000 121.0000 89.2000 ;
	    RECT 114.2000 86.2000 114.5000 88.8000 ;
	    RECT 116.6000 87.8000 117.0000 88.2000 ;
	    RECT 115.0000 86.8000 115.4000 87.2000 ;
	    RECT 115.0000 86.2000 115.3000 86.8000 ;
	    RECT 101.4000 86.1000 101.8000 86.2000 ;
	    RECT 102.2000 86.1000 102.6000 86.2000 ;
	    RECT 101.4000 85.8000 102.6000 86.1000 ;
	    RECT 104.6000 85.8000 105.0000 86.2000 ;
	    RECT 111.8000 85.8000 112.2000 86.2000 ;
	    RECT 112.6000 85.8000 113.0000 86.2000 ;
	    RECT 113.4000 85.8000 113.8000 86.2000 ;
	    RECT 114.2000 85.8000 114.6000 86.2000 ;
	    RECT 115.0000 85.8000 115.4000 86.2000 ;
	    RECT 100.6000 84.8000 101.0000 85.2000 ;
	    RECT 101.4000 79.8000 101.8000 80.2000 ;
	    RECT 101.4000 75.2000 101.7000 79.8000 ;
	    RECT 100.6000 74.8000 101.0000 75.2000 ;
	    RECT 101.4000 74.8000 101.8000 75.2000 ;
	    RECT 100.6000 74.2000 100.9000 74.8000 ;
	    RECT 100.6000 73.8000 101.0000 74.2000 ;
	    RECT 99.0000 71.8000 99.4000 72.2000 ;
	    RECT 98.2000 70.8000 98.6000 71.2000 ;
	    RECT 95.8000 69.1000 96.2000 69.2000 ;
	    RECT 96.6000 69.1000 97.0000 69.2000 ;
	    RECT 95.8000 68.8000 97.0000 69.1000 ;
	    RECT 98.2000 67.2000 98.5000 70.8000 ;
	    RECT 99.0000 70.2000 99.3000 71.8000 ;
	    RECT 99.0000 69.8000 99.4000 70.2000 ;
	    RECT 101.4000 68.1000 101.7000 74.8000 ;
	    RECT 102.2000 73.8000 102.6000 74.2000 ;
	    RECT 103.8000 73.8000 104.2000 74.2000 ;
	    RECT 102.2000 73.2000 102.5000 73.8000 ;
	    RECT 103.8000 73.2000 104.1000 73.8000 ;
	    RECT 102.2000 72.8000 102.6000 73.2000 ;
	    RECT 103.8000 72.8000 104.2000 73.2000 ;
	    RECT 103.0000 71.8000 103.4000 72.2000 ;
	    RECT 101.4000 67.8000 102.5000 68.1000 ;
	    RECT 98.2000 66.8000 98.6000 67.2000 ;
	    RECT 101.4000 66.8000 101.8000 67.2000 ;
	    RECT 101.4000 66.2000 101.7000 66.8000 ;
	    RECT 97.4000 66.1000 97.8000 66.2000 ;
	    RECT 98.2000 66.1000 98.6000 66.2000 ;
	    RECT 97.4000 65.8000 98.6000 66.1000 ;
	    RECT 99.8000 66.1000 100.2000 66.2000 ;
	    RECT 100.6000 66.1000 101.0000 66.2000 ;
	    RECT 99.8000 65.8000 101.0000 66.1000 ;
	    RECT 101.4000 65.8000 101.8000 66.2000 ;
	    RECT 95.0000 60.8000 95.4000 61.2000 ;
	    RECT 90.2000 58.8000 90.6000 59.2000 ;
	    RECT 80.6000 56.8000 81.0000 57.2000 ;
	    RECT 84.6000 56.8000 85.0000 57.2000 ;
	    RECT 76.6000 55.1000 77.0000 55.2000 ;
	    RECT 77.4000 55.1000 77.8000 55.2000 ;
	    RECT 76.6000 54.8000 77.8000 55.1000 ;
	    RECT 79.0000 54.2000 79.3000 56.8000 ;
	    RECT 79.8000 55.8000 80.2000 56.2000 ;
	    RECT 79.8000 55.2000 80.1000 55.8000 ;
	    RECT 79.8000 54.8000 80.2000 55.2000 ;
	    RECT 81.4000 54.8000 81.8000 55.2000 ;
	    RECT 82.2000 54.8000 82.6000 55.2000 ;
	    RECT 75.8000 53.8000 76.2000 54.2000 ;
	    RECT 76.6000 53.8000 77.0000 54.2000 ;
	    RECT 79.0000 53.8000 79.4000 54.2000 ;
	    RECT 76.6000 49.2000 76.9000 53.8000 ;
	    RECT 79.0000 53.2000 79.3000 53.8000 ;
	    RECT 81.4000 53.2000 81.7000 54.8000 ;
	    RECT 79.0000 52.8000 79.4000 53.2000 ;
	    RECT 81.4000 52.8000 81.8000 53.2000 ;
	    RECT 78.2000 51.8000 78.6000 52.2000 ;
	    RECT 76.6000 48.8000 77.0000 49.2000 ;
	    RECT 78.2000 48.1000 78.5000 51.8000 ;
	    RECT 77.4000 47.8000 78.5000 48.1000 ;
	    RECT 79.0000 49.8000 79.4000 50.2000 ;
	    RECT 75.0000 46.8000 75.4000 47.2000 ;
	    RECT 72.6000 45.8000 73.0000 46.2000 ;
	    RECT 74.2000 46.1000 74.6000 46.2000 ;
	    RECT 75.0000 46.1000 75.4000 46.2000 ;
	    RECT 74.2000 45.8000 75.4000 46.1000 ;
	    RECT 75.8000 45.8000 76.2000 46.2000 ;
	    RECT 75.8000 45.2000 76.1000 45.8000 ;
	    RECT 75.8000 44.8000 76.2000 45.2000 ;
	    RECT 76.6000 43.8000 77.0000 44.2000 ;
	    RECT 71.0000 35.8000 71.4000 36.2000 ;
	    RECT 69.4000 35.1000 69.8000 35.2000 ;
	    RECT 70.2000 35.1000 70.6000 35.2000 ;
	    RECT 69.4000 34.8000 70.6000 35.1000 ;
	    RECT 67.8000 31.8000 68.2000 32.2000 ;
	    RECT 67.8000 29.2000 68.1000 31.8000 ;
	    RECT 67.8000 28.8000 68.2000 29.2000 ;
	    RECT 67.0000 27.8000 68.1000 28.1000 ;
	    RECT 67.8000 27.2000 68.1000 27.8000 ;
	    RECT 68.6000 27.8000 69.0000 28.2000 ;
	    RECT 65.4000 26.8000 65.8000 27.2000 ;
	    RECT 67.8000 26.8000 68.2000 27.2000 ;
	    RECT 65.4000 19.2000 65.7000 26.8000 ;
	    RECT 66.2000 24.1000 66.6000 24.2000 ;
	    RECT 67.0000 24.1000 67.4000 24.2000 ;
	    RECT 66.2000 23.8000 67.4000 24.1000 ;
	    RECT 65.4000 18.8000 65.8000 19.2000 ;
	    RECT 67.8000 18.2000 68.1000 26.8000 ;
	    RECT 68.6000 26.2000 68.9000 27.8000 ;
	    RECT 71.0000 26.2000 71.3000 35.8000 ;
	    RECT 71.8000 32.1000 72.2000 32.2000 ;
	    RECT 72.6000 32.1000 73.0000 32.2000 ;
	    RECT 74.2000 32.1000 74.6000 37.9000 ;
	    RECT 76.6000 35.2000 76.9000 43.8000 ;
	    RECT 77.4000 39.2000 77.7000 47.8000 ;
	    RECT 79.0000 47.2000 79.3000 49.8000 ;
	    RECT 82.2000 49.2000 82.5000 54.8000 ;
	    RECT 83.0000 51.8000 83.4000 52.2000 ;
	    RECT 78.2000 46.8000 78.6000 47.2000 ;
	    RECT 79.0000 46.8000 79.4000 47.2000 ;
	    RECT 78.2000 46.2000 78.5000 46.8000 ;
	    RECT 78.2000 45.8000 78.6000 46.2000 ;
	    RECT 79.8000 45.1000 80.2000 47.9000 ;
	    RECT 81.4000 43.1000 81.8000 48.9000 ;
	    RECT 82.2000 48.8000 82.6000 49.2000 ;
	    RECT 83.0000 48.2000 83.3000 51.8000 ;
	    RECT 83.0000 47.8000 83.4000 48.2000 ;
	    RECT 82.2000 45.9000 82.6000 46.3000 ;
	    RECT 82.2000 45.2000 82.5000 45.9000 ;
	    RECT 82.2000 44.8000 82.6000 45.2000 ;
	    RECT 83.0000 43.2000 83.3000 47.8000 ;
	    RECT 84.6000 46.2000 84.9000 56.8000 ;
	    RECT 85.4000 52.1000 85.8000 57.9000 ;
	    RECT 89.4000 54.7000 89.8000 55.1000 ;
	    RECT 89.4000 51.2000 89.7000 54.7000 ;
	    RECT 90.2000 52.1000 90.6000 57.9000 ;
	    RECT 91.0000 54.8000 91.4000 55.2000 ;
	    RECT 91.0000 54.2000 91.3000 54.8000 ;
	    RECT 91.0000 53.8000 91.4000 54.2000 ;
	    RECT 91.8000 53.1000 92.2000 55.9000 ;
	    RECT 95.0000 55.2000 95.3000 60.8000 ;
	    RECT 98.2000 60.2000 98.5000 65.8000 ;
	    RECT 99.0000 61.8000 99.4000 62.2000 ;
	    RECT 98.2000 59.8000 98.6000 60.2000 ;
	    RECT 98.2000 55.2000 98.5000 59.8000 ;
	    RECT 99.0000 56.2000 99.3000 61.8000 ;
	    RECT 99.0000 55.8000 99.4000 56.2000 ;
	    RECT 95.0000 54.8000 95.4000 55.2000 ;
	    RECT 98.2000 54.8000 98.6000 55.2000 ;
	    RECT 99.0000 54.2000 99.3000 55.8000 ;
	    RECT 102.2000 55.2000 102.5000 67.8000 ;
	    RECT 103.0000 57.2000 103.3000 71.8000 ;
	    RECT 104.6000 66.2000 104.9000 85.8000 ;
	    RECT 116.6000 85.2000 116.9000 87.8000 ;
	    RECT 116.6000 84.8000 117.0000 85.2000 ;
	    RECT 115.0000 83.8000 115.4000 84.2000 ;
	    RECT 115.0000 83.2000 115.3000 83.8000 ;
	    RECT 115.0000 82.8000 115.4000 83.2000 ;
	    RECT 117.4000 82.8000 117.8000 83.2000 ;
	    RECT 123.0000 83.1000 123.4000 88.9000 ;
	    RECT 123.8000 85.2000 124.1000 91.8000 ;
	    RECT 124.6000 86.2000 124.9000 94.8000 ;
	    RECT 126.2000 92.8000 126.6000 93.2000 ;
	    RECT 126.2000 90.2000 126.5000 92.8000 ;
	    RECT 127.0000 91.8000 127.4000 92.2000 ;
	    RECT 127.8000 92.1000 128.2000 92.2000 ;
	    RECT 128.6000 92.1000 129.0000 92.2000 ;
	    RECT 130.2000 92.1000 130.6000 97.9000 ;
	    RECT 134.2000 94.7000 134.6000 95.1000 ;
	    RECT 127.8000 91.8000 129.0000 92.1000 ;
	    RECT 131.8000 91.8000 132.2000 92.2000 ;
	    RECT 126.2000 89.8000 126.6000 90.2000 ;
	    RECT 127.0000 88.2000 127.3000 91.8000 ;
	    RECT 127.0000 87.8000 127.4000 88.2000 ;
	    RECT 127.0000 86.8000 127.4000 87.2000 ;
	    RECT 127.0000 86.3000 127.3000 86.8000 ;
	    RECT 124.6000 85.8000 125.0000 86.2000 ;
	    RECT 127.0000 85.9000 127.4000 86.3000 ;
	    RECT 123.8000 84.8000 124.2000 85.2000 ;
	    RECT 105.4000 81.8000 105.8000 82.2000 ;
	    RECT 105.4000 66.2000 105.7000 81.8000 ;
	    RECT 117.4000 79.2000 117.7000 82.8000 ;
	    RECT 117.4000 78.8000 117.8000 79.2000 ;
	    RECT 106.2000 73.1000 106.6000 75.9000 ;
	    RECT 107.0000 71.8000 107.4000 72.2000 ;
	    RECT 107.8000 72.1000 108.2000 77.9000 ;
	    RECT 108.6000 75.8000 109.0000 76.2000 ;
	    RECT 108.6000 75.1000 108.9000 75.8000 ;
	    RECT 111.0000 75.1000 111.4000 75.2000 ;
	    RECT 111.8000 75.1000 112.2000 75.2000 ;
	    RECT 108.6000 74.7000 109.0000 75.1000 ;
	    RECT 111.0000 74.8000 112.2000 75.1000 ;
	    RECT 112.6000 72.1000 113.0000 77.9000 ;
	    RECT 115.8000 74.8000 116.2000 75.2000 ;
	    RECT 118.2000 74.8000 118.6000 75.2000 ;
	    RECT 115.8000 72.2000 116.1000 74.8000 ;
	    RECT 118.2000 74.2000 118.5000 74.8000 ;
	    RECT 118.2000 73.8000 118.6000 74.2000 ;
	    RECT 119.0000 73.1000 119.4000 75.9000 ;
	    RECT 119.8000 74.8000 120.2000 75.2000 ;
	    RECT 115.0000 71.8000 115.4000 72.2000 ;
	    RECT 115.8000 71.8000 116.2000 72.2000 ;
	    RECT 117.4000 71.8000 117.8000 72.2000 ;
	    RECT 107.0000 66.2000 107.3000 71.8000 ;
	    RECT 107.8000 68.8000 108.2000 69.2000 ;
	    RECT 107.8000 66.2000 108.1000 68.8000 ;
	    RECT 111.8000 66.8000 112.2000 67.2000 ;
	    RECT 111.8000 66.2000 112.1000 66.8000 ;
	    RECT 115.0000 66.2000 115.3000 71.8000 ;
	    RECT 117.4000 70.2000 117.7000 71.8000 ;
	    RECT 117.4000 69.8000 117.8000 70.2000 ;
	    RECT 119.8000 69.2000 120.1000 74.8000 ;
	    RECT 120.6000 72.1000 121.0000 77.9000 ;
	    RECT 124.6000 75.2000 124.9000 85.8000 ;
	    RECT 127.8000 83.1000 128.2000 88.9000 ;
	    RECT 130.2000 88.8000 130.6000 89.2000 ;
	    RECT 130.2000 88.2000 130.5000 88.8000 ;
	    RECT 131.8000 88.2000 132.1000 91.8000 ;
	    RECT 129.4000 85.1000 129.8000 87.9000 ;
	    RECT 130.2000 87.8000 130.6000 88.2000 ;
	    RECT 131.8000 87.8000 132.2000 88.2000 ;
	    RECT 134.2000 87.2000 134.5000 94.7000 ;
	    RECT 135.0000 92.1000 135.4000 97.9000 ;
	    RECT 135.8000 93.8000 136.2000 94.2000 ;
	    RECT 135.8000 87.2000 136.1000 93.8000 ;
	    RECT 136.6000 93.1000 137.0000 95.9000 ;
	    RECT 137.4000 94.8000 137.8000 95.2000 ;
	    RECT 130.2000 86.8000 130.6000 87.2000 ;
	    RECT 134.2000 86.8000 134.6000 87.2000 ;
	    RECT 135.8000 86.8000 136.2000 87.2000 ;
	    RECT 130.2000 86.2000 130.5000 86.8000 ;
	    RECT 130.2000 85.8000 130.6000 86.2000 ;
	    RECT 131.8000 85.8000 132.2000 86.2000 ;
	    RECT 135.8000 85.8000 136.2000 86.2000 ;
	    RECT 131.8000 82.2000 132.1000 85.8000 ;
	    RECT 135.8000 82.2000 136.1000 85.8000 ;
	    RECT 136.6000 85.1000 137.0000 87.9000 ;
	    RECT 137.4000 83.2000 137.7000 94.8000 ;
	    RECT 138.2000 93.8000 138.6000 94.2000 ;
	    RECT 139.0000 94.1000 139.3000 104.8000 ;
	    RECT 140.6000 103.1000 141.0000 108.9000 ;
	    RECT 144.6000 108.2000 144.9000 111.8000 ;
	    RECT 142.2000 105.1000 142.6000 107.9000 ;
	    RECT 143.0000 107.8000 143.4000 108.2000 ;
	    RECT 144.6000 107.8000 145.0000 108.2000 ;
	    RECT 143.0000 106.2000 143.3000 107.8000 ;
	    RECT 143.0000 105.8000 143.4000 106.2000 ;
	    RECT 143.8000 106.1000 144.2000 106.2000 ;
	    RECT 144.6000 106.1000 145.0000 106.2000 ;
	    RECT 143.8000 105.8000 145.0000 106.1000 ;
	    RECT 144.6000 104.8000 145.0000 105.2000 ;
	    RECT 144.6000 99.2000 144.9000 104.8000 ;
	    RECT 144.6000 98.8000 145.0000 99.2000 ;
	    RECT 146.2000 97.2000 146.5000 112.8000 ;
	    RECT 147.0000 109.2000 147.3000 112.8000 ;
	    RECT 147.8000 111.8000 148.2000 112.2000 ;
	    RECT 147.0000 108.8000 147.4000 109.2000 ;
	    RECT 147.8000 108.2000 148.1000 111.8000 ;
	    RECT 148.6000 110.8000 149.0000 111.2000 ;
	    RECT 147.8000 107.8000 148.2000 108.2000 ;
	    RECT 148.6000 106.2000 148.9000 110.8000 ;
	    RECT 149.4000 109.2000 149.7000 113.8000 ;
	    RECT 150.2000 113.2000 150.5000 113.8000 ;
	    RECT 150.2000 112.8000 150.6000 113.2000 ;
	    RECT 155.0000 112.8000 155.4000 113.2000 ;
	    RECT 155.0000 112.2000 155.3000 112.8000 ;
	    RECT 155.0000 111.8000 155.4000 112.2000 ;
	    RECT 153.4000 109.8000 153.8000 110.2000 ;
	    RECT 155.8000 109.8000 156.2000 110.2000 ;
	    RECT 149.4000 108.8000 149.8000 109.2000 ;
	    RECT 150.2000 106.8000 150.6000 107.2000 ;
	    RECT 153.4000 107.0000 153.7000 109.8000 ;
	    RECT 155.0000 107.8000 155.4000 108.2000 ;
	    RECT 155.0000 107.2000 155.3000 107.8000 ;
	    RECT 155.8000 107.2000 156.1000 109.8000 ;
	    RECT 159.8000 109.2000 160.1000 118.8000 ;
	    RECT 160.6000 113.1000 161.0000 115.9000 ;
	    RECT 162.2000 112.1000 162.6000 117.9000 ;
	    RECT 163.0000 114.7000 163.4000 115.1000 ;
	    RECT 163.0000 114.2000 163.3000 114.7000 ;
	    RECT 163.0000 113.8000 163.4000 114.2000 ;
	    RECT 164.6000 113.8000 165.0000 114.2000 ;
	    RECT 163.8000 112.8000 164.2000 113.2000 ;
	    RECT 159.8000 108.8000 160.2000 109.2000 ;
	    RECT 163.0000 108.8000 163.4000 109.2000 ;
	    RECT 163.0000 108.2000 163.3000 108.8000 ;
	    RECT 163.8000 108.2000 164.1000 112.8000 ;
	    RECT 158.2000 107.8000 158.6000 108.2000 ;
	    RECT 162.2000 107.8000 162.6000 108.2000 ;
	    RECT 163.0000 107.8000 163.4000 108.2000 ;
	    RECT 163.8000 107.8000 164.2000 108.2000 ;
	    RECT 150.2000 106.2000 150.5000 106.8000 ;
	    RECT 153.4000 106.6000 153.8000 107.0000 ;
	    RECT 155.0000 106.8000 155.4000 107.2000 ;
	    RECT 155.8000 106.8000 156.2000 107.2000 ;
	    RECT 148.6000 105.8000 149.0000 106.2000 ;
	    RECT 150.2000 105.8000 150.6000 106.2000 ;
	    RECT 155.0000 105.2000 155.3000 106.8000 ;
	    RECT 158.2000 106.2000 158.5000 107.8000 ;
	    RECT 162.2000 106.2000 162.5000 107.8000 ;
	    RECT 163.0000 106.8000 163.4000 107.2000 ;
	    RECT 158.2000 105.8000 158.6000 106.2000 ;
	    RECT 162.2000 105.8000 162.6000 106.2000 ;
	    RECT 155.0000 104.8000 155.4000 105.2000 ;
	    RECT 142.2000 96.8000 142.6000 97.2000 ;
	    RECT 145.4000 96.8000 145.8000 97.2000 ;
	    RECT 146.2000 96.8000 146.6000 97.2000 ;
	    RECT 139.8000 96.1000 140.2000 96.2000 ;
	    RECT 140.6000 96.1000 141.0000 96.2000 ;
	    RECT 139.8000 95.8000 141.0000 96.1000 ;
	    RECT 142.2000 95.2000 142.5000 96.8000 ;
	    RECT 142.2000 94.8000 142.6000 95.2000 ;
	    RECT 139.8000 94.1000 140.2000 94.2000 ;
	    RECT 139.0000 93.8000 140.2000 94.1000 ;
	    RECT 143.8000 93.8000 144.2000 94.2000 ;
	    RECT 138.2000 93.2000 138.5000 93.8000 ;
	    RECT 138.2000 92.8000 138.6000 93.2000 ;
	    RECT 139.0000 91.8000 139.4000 92.2000 ;
	    RECT 137.4000 82.8000 137.8000 83.2000 ;
	    RECT 138.2000 83.1000 138.6000 88.9000 ;
	    RECT 139.0000 86.3000 139.3000 91.8000 ;
	    RECT 139.0000 85.9000 139.4000 86.3000 ;
	    RECT 131.8000 81.8000 132.2000 82.2000 ;
	    RECT 135.8000 81.8000 136.2000 82.2000 ;
	    RECT 139.8000 79.2000 140.1000 93.8000 ;
	    RECT 143.8000 93.2000 144.1000 93.8000 ;
	    RECT 142.2000 92.8000 142.6000 93.2000 ;
	    RECT 143.8000 92.8000 144.2000 93.2000 ;
	    RECT 141.4000 85.8000 141.8000 86.2000 ;
	    RECT 141.4000 84.2000 141.7000 85.8000 ;
	    RECT 141.4000 83.8000 141.8000 84.2000 ;
	    RECT 142.2000 79.2000 142.5000 92.8000 ;
	    RECT 145.4000 89.2000 145.7000 96.8000 ;
	    RECT 146.2000 95.8000 146.6000 96.2000 ;
	    RECT 146.2000 89.2000 146.5000 95.8000 ;
	    RECT 152.6000 93.8000 153.0000 94.2000 ;
	    RECT 152.6000 92.2000 152.9000 93.8000 ;
	    RECT 154.2000 93.1000 154.6000 95.9000 ;
	    RECT 155.0000 93.8000 155.4000 94.2000 ;
	    RECT 155.0000 93.2000 155.3000 93.8000 ;
	    RECT 155.0000 92.8000 155.4000 93.2000 ;
	    RECT 152.6000 91.8000 153.0000 92.2000 ;
	    RECT 155.8000 92.1000 156.2000 97.9000 ;
	    RECT 157.4000 95.1000 157.8000 95.2000 ;
	    RECT 158.2000 95.1000 158.6000 95.2000 ;
	    RECT 157.4000 94.8000 158.6000 95.1000 ;
	    RECT 157.4000 92.8000 157.8000 93.2000 ;
	    RECT 143.0000 83.1000 143.4000 88.9000 ;
	    RECT 145.4000 88.8000 145.8000 89.2000 ;
	    RECT 146.2000 88.8000 146.6000 89.2000 ;
	    RECT 145.4000 88.2000 145.7000 88.8000 ;
	    RECT 145.4000 87.8000 145.8000 88.2000 ;
	    RECT 148.6000 83.1000 149.0000 88.9000 ;
	    RECT 152.6000 88.2000 152.9000 91.8000 ;
	    RECT 157.4000 89.2000 157.7000 92.8000 ;
	    RECT 160.6000 92.1000 161.0000 97.9000 ;
	    RECT 161.4000 97.8000 161.8000 98.2000 ;
	    RECT 161.4000 97.2000 161.7000 97.8000 ;
	    RECT 161.4000 96.8000 161.8000 97.2000 ;
	    RECT 162.2000 93.2000 162.5000 105.8000 ;
	    RECT 163.0000 99.2000 163.3000 106.8000 ;
	    RECT 163.8000 105.8000 164.2000 106.2000 ;
	    RECT 163.8000 105.2000 164.1000 105.8000 ;
	    RECT 163.8000 104.8000 164.2000 105.2000 ;
	    RECT 163.0000 98.8000 163.4000 99.2000 ;
	    RECT 164.6000 97.2000 164.9000 113.8000 ;
	    RECT 165.4000 111.8000 165.8000 112.2000 ;
	    RECT 165.4000 109.2000 165.7000 111.8000 ;
	    RECT 165.4000 108.8000 165.8000 109.2000 ;
	    RECT 166.2000 107.2000 166.5000 132.8000 ;
	    RECT 167.0000 123.1000 167.4000 128.9000 ;
	    RECT 167.8000 126.8000 168.2000 127.2000 ;
	    RECT 167.0000 112.1000 167.4000 117.9000 ;
	    RECT 167.8000 117.2000 168.1000 126.8000 ;
	    RECT 168.6000 125.8000 169.0000 126.2000 ;
	    RECT 168.6000 119.2000 168.9000 125.8000 ;
	    RECT 169.4000 119.2000 169.7000 135.8000 ;
	    RECT 179.0000 135.2000 179.3000 144.8000 ;
	    RECT 180.6000 143.8000 181.0000 144.2000 ;
	    RECT 174.2000 135.1000 174.6000 135.2000 ;
	    RECT 175.0000 135.1000 175.4000 135.2000 ;
	    RECT 174.2000 134.8000 175.4000 135.1000 ;
	    RECT 176.6000 134.8000 177.0000 135.2000 ;
	    RECT 179.0000 134.8000 179.4000 135.2000 ;
	    RECT 175.8000 133.8000 176.2000 134.2000 ;
	    RECT 175.8000 129.2000 176.1000 133.8000 ;
	    RECT 176.6000 133.2000 176.9000 134.8000 ;
	    RECT 176.6000 132.8000 177.0000 133.2000 ;
	    RECT 180.6000 129.2000 180.9000 143.8000 ;
	    RECT 181.4000 134.2000 181.7000 145.8000 ;
	    RECT 182.2000 135.1000 182.6000 135.2000 ;
	    RECT 183.0000 135.1000 183.4000 135.2000 ;
	    RECT 182.2000 134.8000 183.4000 135.1000 ;
	    RECT 181.4000 133.8000 181.8000 134.2000 ;
	    RECT 183.0000 134.1000 183.4000 134.2000 ;
	    RECT 183.8000 134.1000 184.2000 134.2000 ;
	    RECT 183.0000 133.8000 184.2000 134.1000 ;
	    RECT 171.8000 123.1000 172.2000 128.9000 ;
	    RECT 174.2000 128.8000 174.6000 129.2000 ;
	    RECT 175.8000 128.8000 176.2000 129.2000 ;
	    RECT 180.6000 128.8000 181.0000 129.2000 ;
	    RECT 174.2000 126.2000 174.5000 128.8000 ;
	    RECT 180.6000 127.8000 181.0000 128.2000 ;
	    RECT 176.6000 127.1000 177.0000 127.2000 ;
	    RECT 177.4000 127.1000 177.8000 127.2000 ;
	    RECT 176.6000 126.8000 177.8000 127.1000 ;
	    RECT 174.2000 125.8000 174.6000 126.2000 ;
	    RECT 175.0000 124.8000 175.4000 125.2000 ;
	    RECT 168.6000 118.8000 169.0000 119.2000 ;
	    RECT 169.4000 118.8000 169.8000 119.2000 ;
	    RECT 167.8000 116.8000 168.2000 117.2000 ;
	    RECT 167.8000 116.2000 168.1000 116.8000 ;
	    RECT 167.8000 115.8000 168.2000 116.2000 ;
	    RECT 169.4000 115.2000 169.7000 118.8000 ;
	    RECT 173.4000 117.8000 173.8000 118.2000 ;
	    RECT 169.4000 114.8000 169.8000 115.2000 ;
	    RECT 173.4000 113.2000 173.7000 117.8000 ;
	    RECT 174.2000 114.8000 174.6000 115.2000 ;
	    RECT 173.4000 112.8000 173.8000 113.2000 ;
	    RECT 174.2000 112.2000 174.5000 114.8000 ;
	    RECT 171.0000 111.8000 171.4000 112.2000 ;
	    RECT 173.4000 111.8000 173.8000 112.2000 ;
	    RECT 174.2000 111.8000 174.6000 112.2000 ;
	    RECT 171.0000 110.2000 171.3000 111.8000 ;
	    RECT 173.4000 111.2000 173.7000 111.8000 ;
	    RECT 173.4000 110.8000 173.8000 111.2000 ;
	    RECT 171.0000 109.8000 171.4000 110.2000 ;
	    RECT 172.6000 108.8000 173.0000 109.2000 ;
	    RECT 171.0000 107.8000 171.4000 108.2000 ;
	    RECT 166.2000 106.8000 166.6000 107.2000 ;
	    RECT 167.0000 107.1000 167.4000 107.2000 ;
	    RECT 167.8000 107.1000 168.2000 107.2000 ;
	    RECT 167.0000 106.8000 168.2000 107.1000 ;
	    RECT 170.2000 106.8000 170.6000 107.2000 ;
	    RECT 166.2000 106.2000 166.5000 106.8000 ;
	    RECT 170.2000 106.2000 170.5000 106.8000 ;
	    RECT 165.4000 105.8000 165.8000 106.2000 ;
	    RECT 166.2000 105.8000 166.6000 106.2000 ;
	    RECT 168.6000 106.1000 169.0000 106.2000 ;
	    RECT 169.4000 106.1000 169.8000 106.2000 ;
	    RECT 168.6000 105.8000 169.8000 106.1000 ;
	    RECT 170.2000 105.8000 170.6000 106.2000 ;
	    RECT 165.4000 104.2000 165.7000 105.8000 ;
	    RECT 171.0000 105.2000 171.3000 107.8000 ;
	    RECT 171.8000 106.8000 172.2000 107.2000 ;
	    RECT 171.8000 106.2000 172.1000 106.8000 ;
	    RECT 171.8000 105.8000 172.2000 106.2000 ;
	    RECT 167.0000 105.1000 167.4000 105.2000 ;
	    RECT 167.8000 105.1000 168.2000 105.2000 ;
	    RECT 167.0000 104.8000 168.2000 105.1000 ;
	    RECT 171.0000 104.8000 171.4000 105.2000 ;
	    RECT 165.4000 103.8000 165.8000 104.2000 ;
	    RECT 166.2000 101.8000 166.6000 102.2000 ;
	    RECT 164.6000 96.8000 165.0000 97.2000 ;
	    RECT 163.8000 95.1000 164.2000 95.2000 ;
	    RECT 164.6000 95.1000 165.0000 95.2000 ;
	    RECT 163.8000 94.8000 165.0000 95.1000 ;
	    RECT 166.2000 94.2000 166.5000 101.8000 ;
	    RECT 168.6000 96.1000 169.0000 96.2000 ;
	    RECT 169.4000 96.1000 169.8000 96.2000 ;
	    RECT 168.6000 95.8000 169.8000 96.1000 ;
	    RECT 171.0000 95.2000 171.3000 104.8000 ;
	    RECT 172.6000 104.2000 172.9000 108.8000 ;
	    RECT 174.2000 107.8000 174.6000 108.2000 ;
	    RECT 174.2000 107.2000 174.5000 107.8000 ;
	    RECT 174.2000 106.8000 174.6000 107.2000 ;
	    RECT 175.0000 105.2000 175.3000 124.8000 ;
	    RECT 176.6000 110.2000 176.9000 126.8000 ;
	    RECT 179.0000 126.1000 179.4000 126.2000 ;
	    RECT 179.8000 126.1000 180.2000 126.2000 ;
	    RECT 179.0000 125.8000 180.2000 126.1000 ;
	    RECT 180.6000 125.2000 180.9000 127.8000 ;
	    RECT 180.6000 124.8000 181.0000 125.2000 ;
	    RECT 178.2000 122.8000 178.6000 123.2000 ;
	    RECT 178.2000 122.2000 178.5000 122.8000 ;
	    RECT 178.2000 121.8000 178.6000 122.2000 ;
	    RECT 178.2000 113.2000 178.5000 121.8000 ;
	    RECT 181.4000 117.2000 181.7000 133.8000 ;
	    RECT 182.2000 127.1000 182.6000 127.2000 ;
	    RECT 183.0000 127.1000 183.4000 127.2000 ;
	    RECT 182.2000 126.8000 183.4000 127.1000 ;
	    RECT 183.8000 121.8000 184.2000 122.2000 ;
	    RECT 183.8000 118.2000 184.1000 121.8000 ;
	    RECT 181.4000 116.8000 181.8000 117.2000 ;
	    RECT 179.0000 115.1000 179.4000 115.2000 ;
	    RECT 179.8000 115.1000 180.2000 115.2000 ;
	    RECT 179.0000 114.8000 180.2000 115.1000 ;
	    RECT 180.6000 114.8000 181.0000 115.2000 ;
	    RECT 180.6000 114.2000 180.9000 114.8000 ;
	    RECT 179.8000 113.8000 180.2000 114.2000 ;
	    RECT 180.6000 113.8000 181.0000 114.2000 ;
	    RECT 178.2000 112.8000 178.6000 113.2000 ;
	    RECT 177.4000 111.8000 177.8000 112.2000 ;
	    RECT 176.6000 109.8000 177.0000 110.2000 ;
	    RECT 177.4000 109.2000 177.7000 111.8000 ;
	    RECT 178.2000 109.8000 178.6000 110.2000 ;
	    RECT 177.4000 108.8000 177.8000 109.2000 ;
	    RECT 177.4000 106.8000 177.8000 107.2000 ;
	    RECT 177.4000 106.2000 177.7000 106.8000 ;
	    RECT 178.2000 106.2000 178.5000 109.8000 ;
	    RECT 179.8000 109.2000 180.1000 113.8000 ;
	    RECT 181.4000 113.1000 181.8000 115.9000 ;
	    RECT 182.2000 115.8000 182.6000 116.2000 ;
	    RECT 182.2000 114.2000 182.5000 115.8000 ;
	    RECT 182.2000 113.8000 182.6000 114.2000 ;
	    RECT 183.0000 112.1000 183.4000 117.9000 ;
	    RECT 183.8000 117.8000 184.2000 118.2000 ;
	    RECT 183.8000 114.7000 184.2000 115.1000 ;
	    RECT 183.8000 114.2000 184.1000 114.7000 ;
	    RECT 183.8000 113.8000 184.2000 114.2000 ;
	    RECT 183.8000 109.8000 184.2000 110.2000 ;
	    RECT 179.0000 108.8000 179.4000 109.2000 ;
	    RECT 179.8000 108.8000 180.2000 109.2000 ;
	    RECT 179.0000 108.2000 179.3000 108.8000 ;
	    RECT 179.0000 107.8000 179.4000 108.2000 ;
	    RECT 180.6000 106.8000 181.0000 107.2000 ;
	    RECT 182.2000 107.1000 182.6000 107.2000 ;
	    RECT 183.0000 107.1000 183.4000 107.2000 ;
	    RECT 182.2000 106.8000 183.4000 107.1000 ;
	    RECT 177.4000 105.8000 177.8000 106.2000 ;
	    RECT 178.2000 105.8000 178.6000 106.2000 ;
	    RECT 178.2000 105.2000 178.5000 105.8000 ;
	    RECT 175.0000 104.8000 175.4000 105.2000 ;
	    RECT 178.2000 104.8000 178.6000 105.2000 ;
	    RECT 175.0000 104.2000 175.3000 104.8000 ;
	    RECT 172.6000 103.8000 173.0000 104.2000 ;
	    RECT 175.0000 103.8000 175.4000 104.2000 ;
	    RECT 175.8000 104.1000 176.2000 104.2000 ;
	    RECT 176.6000 104.1000 177.0000 104.2000 ;
	    RECT 175.8000 103.8000 177.0000 104.1000 ;
	    RECT 180.6000 104.1000 180.9000 106.8000 ;
	    RECT 181.4000 105.8000 181.8000 106.2000 ;
	    RECT 182.2000 106.1000 182.6000 106.2000 ;
	    RECT 183.0000 106.1000 183.4000 106.2000 ;
	    RECT 182.2000 105.8000 183.4000 106.1000 ;
	    RECT 181.4000 105.2000 181.7000 105.8000 ;
	    RECT 181.4000 104.8000 181.8000 105.2000 ;
	    RECT 182.2000 105.1000 182.6000 105.2000 ;
	    RECT 183.0000 105.1000 183.4000 105.2000 ;
	    RECT 182.2000 104.8000 183.4000 105.1000 ;
	    RECT 180.6000 103.8000 181.7000 104.1000 ;
	    RECT 171.8000 101.8000 172.2000 102.2000 ;
	    RECT 177.4000 101.8000 177.8000 102.2000 ;
	    RECT 171.8000 95.2000 172.1000 101.8000 ;
	    RECT 177.4000 98.2000 177.7000 101.8000 ;
	    RECT 175.0000 96.8000 175.4000 97.2000 ;
	    RECT 167.8000 95.1000 168.2000 95.2000 ;
	    RECT 168.6000 95.1000 169.0000 95.2000 ;
	    RECT 167.8000 94.8000 169.0000 95.1000 ;
	    RECT 171.0000 94.8000 171.4000 95.2000 ;
	    RECT 171.8000 94.8000 172.2000 95.2000 ;
	    RECT 166.2000 93.8000 166.6000 94.2000 ;
	    RECT 162.2000 92.8000 162.6000 93.2000 ;
	    RECT 164.6000 93.1000 165.0000 93.2000 ;
	    RECT 165.4000 93.1000 165.8000 93.2000 ;
	    RECT 164.6000 92.8000 165.8000 93.1000 ;
	    RECT 164.6000 91.8000 165.0000 92.2000 ;
	    RECT 152.6000 87.8000 153.0000 88.2000 ;
	    RECT 152.6000 86.8000 153.0000 87.2000 ;
	    RECT 152.6000 86.3000 152.9000 86.8000 ;
	    RECT 152.6000 85.9000 153.0000 86.3000 ;
	    RECT 152.6000 83.8000 153.0000 84.2000 ;
	    RECT 152.6000 79.2000 152.9000 83.8000 ;
	    RECT 153.4000 83.1000 153.8000 88.9000 ;
	    RECT 157.4000 88.8000 157.8000 89.2000 ;
	    RECT 159.8000 88.8000 160.2000 89.2000 ;
	    RECT 155.0000 85.1000 155.4000 87.9000 ;
	    RECT 155.8000 87.8000 156.2000 88.2000 ;
	    RECT 159.0000 87.8000 159.4000 88.2000 ;
	    RECT 155.8000 87.2000 156.1000 87.8000 ;
	    RECT 159.0000 87.2000 159.3000 87.8000 ;
	    RECT 155.8000 86.8000 156.2000 87.2000 ;
	    RECT 159.0000 86.8000 159.4000 87.2000 ;
	    RECT 139.8000 78.8000 140.2000 79.2000 ;
	    RECT 142.2000 78.8000 142.6000 79.2000 ;
	    RECT 152.6000 78.8000 153.0000 79.2000 ;
	    RECT 121.4000 74.7000 121.8000 75.1000 ;
	    RECT 124.6000 74.8000 125.0000 75.2000 ;
	    RECT 121.4000 74.2000 121.7000 74.7000 ;
	    RECT 124.6000 74.2000 124.9000 74.8000 ;
	    RECT 121.4000 73.8000 121.8000 74.2000 ;
	    RECT 124.6000 73.8000 125.0000 74.2000 ;
	    RECT 125.4000 72.1000 125.8000 77.9000 ;
	    RECT 127.8000 71.8000 128.2000 72.2000 ;
	    RECT 128.6000 72.1000 129.0000 72.2000 ;
	    RECT 129.4000 72.1000 129.8000 72.2000 ;
	    RECT 131.0000 72.1000 131.4000 77.9000 ;
	    RECT 135.0000 74.7000 135.4000 75.1000 ;
	    RECT 128.6000 71.8000 129.8000 72.1000 ;
	    RECT 120.6000 70.8000 121.0000 71.2000 ;
	    RECT 125.4000 70.8000 125.8000 71.2000 ;
	    RECT 119.8000 68.8000 120.2000 69.2000 ;
	    RECT 119.0000 67.8000 119.4000 68.2000 ;
	    RECT 119.0000 67.2000 119.3000 67.8000 ;
	    RECT 120.6000 67.2000 120.9000 70.8000 ;
	    RECT 123.0000 69.8000 123.4000 70.2000 ;
	    RECT 119.0000 66.8000 119.4000 67.2000 ;
	    RECT 120.6000 66.8000 121.0000 67.2000 ;
	    RECT 104.6000 65.8000 105.0000 66.2000 ;
	    RECT 105.4000 65.8000 105.8000 66.2000 ;
	    RECT 107.0000 65.8000 107.4000 66.2000 ;
	    RECT 107.8000 65.8000 108.2000 66.2000 ;
	    RECT 111.8000 65.8000 112.2000 66.2000 ;
	    RECT 112.6000 65.8000 113.0000 66.2000 ;
	    RECT 115.0000 65.8000 115.4000 66.2000 ;
	    RECT 116.6000 65.8000 117.0000 66.2000 ;
	    RECT 118.2000 65.8000 118.6000 66.2000 ;
	    RECT 104.6000 65.2000 104.9000 65.8000 ;
	    RECT 107.8000 65.2000 108.1000 65.8000 ;
	    RECT 104.6000 64.8000 105.0000 65.2000 ;
	    RECT 107.8000 64.8000 108.2000 65.2000 ;
	    RECT 105.4000 63.8000 105.8000 64.2000 ;
	    RECT 105.4000 63.2000 105.7000 63.8000 ;
	    RECT 105.4000 62.8000 105.8000 63.2000 ;
	    RECT 109.4000 59.1000 109.8000 59.2000 ;
	    RECT 110.2000 59.1000 110.6000 59.2000 ;
	    RECT 109.4000 58.8000 110.6000 59.1000 ;
	    RECT 112.6000 58.2000 112.9000 65.8000 ;
	    RECT 114.2000 64.8000 114.6000 65.2000 ;
	    RECT 114.2000 64.2000 114.5000 64.8000 ;
	    RECT 114.2000 63.8000 114.6000 64.2000 ;
	    RECT 116.6000 62.2000 116.9000 65.8000 ;
	    RECT 118.2000 65.2000 118.5000 65.8000 ;
	    RECT 118.2000 64.8000 118.6000 65.2000 ;
	    RECT 117.4000 63.8000 117.8000 64.2000 ;
	    RECT 117.4000 63.2000 117.7000 63.8000 ;
	    RECT 117.4000 62.8000 117.8000 63.2000 ;
	    RECT 116.6000 61.8000 117.0000 62.2000 ;
	    RECT 108.6000 57.8000 109.0000 58.2000 ;
	    RECT 103.0000 56.8000 103.4000 57.2000 ;
	    RECT 106.2000 56.8000 106.6000 57.2000 ;
	    RECT 103.0000 56.1000 103.4000 56.2000 ;
	    RECT 103.8000 56.1000 104.2000 56.2000 ;
	    RECT 103.0000 55.8000 104.2000 56.1000 ;
	    RECT 99.8000 55.1000 100.2000 55.2000 ;
	    RECT 100.6000 55.1000 101.0000 55.2000 ;
	    RECT 99.8000 54.8000 101.0000 55.1000 ;
	    RECT 102.2000 54.8000 102.6000 55.2000 ;
	    RECT 102.2000 54.2000 102.5000 54.8000 ;
	    RECT 99.0000 53.8000 99.4000 54.2000 ;
	    RECT 102.2000 53.8000 102.6000 54.2000 ;
	    RECT 93.4000 52.8000 93.8000 53.2000 ;
	    RECT 93.4000 52.2000 93.7000 52.8000 ;
	    RECT 93.4000 51.8000 93.8000 52.2000 ;
	    RECT 96.6000 51.8000 97.0000 52.2000 ;
	    RECT 101.4000 51.8000 101.8000 52.2000 ;
	    RECT 103.8000 51.8000 104.2000 52.2000 ;
	    RECT 105.4000 51.8000 105.8000 52.2000 ;
	    RECT 89.4000 50.8000 89.8000 51.2000 ;
	    RECT 87.8000 49.1000 88.2000 49.2000 ;
	    RECT 88.6000 49.1000 89.0000 49.2000 ;
	    RECT 83.8000 45.8000 84.2000 46.2000 ;
	    RECT 84.6000 45.8000 85.0000 46.2000 ;
	    RECT 83.0000 42.8000 83.4000 43.2000 ;
	    RECT 82.2000 39.8000 82.6000 40.2000 ;
	    RECT 77.4000 38.8000 77.8000 39.2000 ;
	    RECT 78.2000 36.8000 78.6000 37.2000 ;
	    RECT 76.6000 34.8000 77.0000 35.2000 ;
	    RECT 78.2000 35.1000 78.5000 36.8000 ;
	    RECT 78.2000 34.7000 78.6000 35.1000 ;
	    RECT 78.2000 32.8000 78.6000 33.2000 ;
	    RECT 71.8000 31.8000 73.0000 32.1000 ;
	    RECT 76.6000 31.8000 77.0000 32.2000 ;
	    RECT 72.6000 28.8000 73.0000 29.2000 ;
	    RECT 72.6000 28.2000 72.9000 28.8000 ;
	    RECT 72.6000 27.8000 73.0000 28.2000 ;
	    RECT 68.6000 25.8000 69.0000 26.2000 ;
	    RECT 70.2000 25.8000 70.6000 26.2000 ;
	    RECT 71.0000 25.8000 71.4000 26.2000 ;
	    RECT 70.2000 25.2000 70.5000 25.8000 ;
	    RECT 70.2000 24.8000 70.6000 25.2000 ;
	    RECT 71.8000 24.8000 72.2000 25.2000 ;
	    RECT 73.4000 25.1000 73.8000 27.9000 ;
	    RECT 71.8000 24.2000 72.1000 24.8000 ;
	    RECT 71.8000 23.8000 72.2000 24.2000 ;
	    RECT 75.0000 23.1000 75.4000 28.9000 ;
	    RECT 75.8000 25.9000 76.2000 26.3000 ;
	    RECT 75.8000 25.2000 76.1000 25.9000 ;
	    RECT 75.8000 24.8000 76.2000 25.2000 ;
	    RECT 68.6000 21.8000 69.0000 22.2000 ;
	    RECT 67.8000 17.8000 68.2000 18.2000 ;
	    RECT 63.0000 16.8000 63.4000 17.2000 ;
	    RECT 63.0000 16.2000 63.3000 16.8000 ;
	    RECT 59.0000 15.8000 59.4000 16.2000 ;
	    RECT 63.0000 15.8000 63.4000 16.2000 ;
	    RECT 63.8000 15.8000 64.2000 16.2000 ;
	    RECT 65.4000 15.8000 65.8000 16.2000 ;
	    RECT 59.0000 15.2000 59.3000 15.8000 ;
	    RECT 63.8000 15.2000 64.1000 15.8000 ;
	    RECT 65.4000 15.2000 65.7000 15.8000 ;
	    RECT 68.6000 15.2000 68.9000 21.8000 ;
	    RECT 69.4000 16.8000 69.8000 17.2000 ;
	    RECT 69.4000 16.2000 69.7000 16.8000 ;
	    RECT 69.4000 15.8000 69.8000 16.2000 ;
	    RECT 71.0000 16.1000 71.4000 16.2000 ;
	    RECT 71.8000 16.1000 72.2000 16.2000 ;
	    RECT 71.0000 15.8000 72.2000 16.1000 ;
	    RECT 59.0000 14.8000 59.4000 15.2000 ;
	    RECT 61.4000 14.8000 61.8000 15.2000 ;
	    RECT 63.0000 14.8000 63.4000 15.2000 ;
	    RECT 63.8000 14.8000 64.2000 15.2000 ;
	    RECT 65.4000 14.8000 65.8000 15.2000 ;
	    RECT 67.0000 15.1000 67.4000 15.2000 ;
	    RECT 67.8000 15.1000 68.2000 15.2000 ;
	    RECT 67.0000 14.8000 68.2000 15.1000 ;
	    RECT 68.6000 14.8000 69.0000 15.2000 ;
	    RECT 70.2000 15.1000 70.6000 15.2000 ;
	    RECT 71.0000 15.1000 71.4000 15.2000 ;
	    RECT 70.2000 14.8000 71.4000 15.1000 ;
	    RECT 75.0000 14.8000 75.4000 15.2000 ;
	    RECT 55.8000 13.8000 56.2000 14.2000 ;
	    RECT 59.8000 13.8000 60.2000 14.2000 ;
	    RECT 60.6000 13.8000 61.0000 14.2000 ;
	    RECT 47.0000 12.2000 47.3000 12.8000 ;
	    RECT 50.2000 12.2000 50.5000 12.8000 ;
	    RECT 39.0000 12.1000 39.4000 12.2000 ;
	    RECT 39.8000 12.1000 40.2000 12.2000 ;
	    RECT 39.0000 11.8000 40.2000 12.1000 ;
	    RECT 41.4000 11.8000 41.8000 12.2000 ;
	    RECT 47.0000 11.8000 47.4000 12.2000 ;
	    RECT 50.2000 11.8000 50.6000 12.2000 ;
	    RECT 52.6000 11.8000 53.0000 12.2000 ;
	    RECT 47.0000 10.2000 47.3000 11.8000 ;
	    RECT 47.0000 9.8000 47.4000 10.2000 ;
	    RECT 26.2000 8.8000 26.6000 9.2000 ;
	    RECT 24.6000 7.8000 25.0000 8.2000 ;
	    RECT 24.6000 7.2000 24.9000 7.8000 ;
	    RECT 24.6000 6.8000 25.0000 7.2000 ;
	    RECT 20.6000 6.1000 21.0000 6.2000 ;
	    RECT 19.8000 5.8000 21.0000 6.1000 ;
	    RECT 21.4000 6.1000 21.8000 6.2000 ;
	    RECT 22.2000 6.1000 22.6000 6.2000 ;
	    RECT 21.4000 5.8000 22.6000 6.1000 ;
	    RECT 22.2000 4.8000 22.6000 5.2000 ;
	    RECT 25.4000 5.1000 25.8000 7.9000 ;
	    RECT 22.2000 4.2000 22.5000 4.8000 ;
	    RECT 22.2000 3.8000 22.6000 4.2000 ;
	    RECT 27.0000 3.1000 27.4000 8.9000 ;
	    RECT 27.8000 8.8000 28.2000 9.2000 ;
	    RECT 27.8000 8.2000 28.1000 8.8000 ;
	    RECT 27.8000 7.8000 28.2000 8.2000 ;
	    RECT 27.8000 5.9000 28.2000 6.3000 ;
	    RECT 27.8000 5.2000 28.1000 5.9000 ;
	    RECT 27.8000 4.8000 28.2000 5.2000 ;
	    RECT 31.8000 3.1000 32.2000 8.9000 ;
	    RECT 34.2000 8.8000 34.6000 9.2000 ;
	    RECT 34.2000 8.2000 34.5000 8.8000 ;
	    RECT 34.2000 7.8000 34.6000 8.2000 ;
	    RECT 40.6000 7.8000 41.0000 8.2000 ;
	    RECT 40.6000 7.2000 40.9000 7.8000 ;
	    RECT 39.0000 6.8000 39.4000 7.2000 ;
	    RECT 40.6000 6.8000 41.0000 7.2000 ;
	    RECT 39.0000 6.2000 39.3000 6.8000 ;
	    RECT 37.4000 6.1000 37.8000 6.2000 ;
	    RECT 38.2000 6.1000 38.6000 6.2000 ;
	    RECT 37.4000 5.8000 38.6000 6.1000 ;
	    RECT 39.0000 5.8000 39.4000 6.2000 ;
	    RECT 41.4000 5.1000 41.8000 7.9000 ;
	    RECT 43.0000 3.1000 43.4000 8.9000 ;
	    RECT 43.8000 8.8000 44.2000 9.2000 ;
	    RECT 43.8000 8.2000 44.1000 8.8000 ;
	    RECT 43.8000 7.8000 44.2000 8.2000 ;
	    RECT 43.8000 5.9000 44.2000 6.3000 ;
	    RECT 43.8000 5.2000 44.1000 5.9000 ;
	    RECT 43.8000 4.8000 44.2000 5.2000 ;
	    RECT 47.8000 3.1000 48.2000 8.9000 ;
	    RECT 50.2000 8.8000 50.6000 9.2000 ;
	    RECT 50.2000 8.2000 50.5000 8.8000 ;
	    RECT 50.2000 7.8000 50.6000 8.2000 ;
	    RECT 52.6000 7.2000 52.9000 11.8000 ;
	    RECT 55.8000 9.2000 56.1000 13.8000 ;
	    RECT 56.6000 13.1000 57.0000 13.2000 ;
	    RECT 57.4000 13.1000 57.8000 13.2000 ;
	    RECT 56.6000 12.8000 57.8000 13.1000 ;
	    RECT 58.2000 9.8000 58.6000 10.2000 ;
	    RECT 55.8000 8.8000 56.2000 9.2000 ;
	    RECT 54.1000 7.5000 54.5000 7.9000 ;
	    RECT 55.0000 7.5000 57.1000 7.8000 ;
	    RECT 57.4000 7.5000 57.8000 7.9000 ;
	    RECT 52.6000 7.1000 53.0000 7.2000 ;
	    RECT 53.4000 7.1000 53.8000 7.2000 ;
	    RECT 52.6000 6.8000 53.8000 7.1000 ;
	    RECT 54.1000 5.1000 54.4000 7.5000 ;
	    RECT 55.0000 7.4000 55.4000 7.5000 ;
	    RECT 56.7000 7.4000 57.1000 7.5000 ;
	    RECT 57.5000 7.1000 57.8000 7.5000 ;
	    RECT 55.4000 6.8000 57.8000 7.1000 ;
	    RECT 58.2000 7.2000 58.5000 9.8000 ;
	    RECT 58.2000 6.8000 58.6000 7.2000 ;
	    RECT 55.4000 6.7000 55.8000 6.8000 ;
	    RECT 57.5000 5.1000 57.8000 6.8000 ;
	    RECT 59.8000 6.2000 60.1000 13.8000 ;
	    RECT 60.6000 8.2000 60.9000 13.8000 ;
	    RECT 61.4000 9.2000 61.7000 14.8000 ;
	    RECT 63.0000 14.2000 63.3000 14.8000 ;
	    RECT 68.6000 14.2000 68.9000 14.8000 ;
	    RECT 63.0000 13.8000 63.4000 14.2000 ;
	    RECT 65.4000 14.1000 65.8000 14.2000 ;
	    RECT 66.2000 14.1000 66.6000 14.2000 ;
	    RECT 65.4000 13.8000 66.6000 14.1000 ;
	    RECT 68.6000 13.8000 69.0000 14.2000 ;
	    RECT 71.8000 14.1000 72.2000 14.2000 ;
	    RECT 72.6000 14.1000 73.0000 14.2000 ;
	    RECT 71.8000 13.8000 73.0000 14.1000 ;
	    RECT 67.0000 13.1000 67.4000 13.2000 ;
	    RECT 67.8000 13.1000 68.2000 13.2000 ;
	    RECT 67.0000 12.8000 68.2000 13.1000 ;
	    RECT 75.0000 12.2000 75.3000 14.8000 ;
	    RECT 76.6000 13.2000 76.9000 31.8000 ;
	    RECT 78.2000 26.2000 78.5000 32.8000 ;
	    RECT 79.0000 32.1000 79.4000 37.9000 ;
	    RECT 80.6000 33.1000 81.0000 35.9000 ;
	    RECT 82.2000 35.2000 82.5000 39.8000 ;
	    RECT 83.8000 39.2000 84.1000 45.8000 ;
	    RECT 86.2000 43.1000 86.6000 48.9000 ;
	    RECT 87.8000 48.8000 89.0000 49.1000 ;
	    RECT 91.8000 48.8000 92.2000 49.2000 ;
	    RECT 89.4000 47.8000 89.8000 48.2000 ;
	    RECT 90.2000 47.8000 90.6000 48.2000 ;
	    RECT 89.4000 45.2000 89.7000 47.8000 ;
	    RECT 90.2000 47.2000 90.5000 47.8000 ;
	    RECT 91.8000 47.2000 92.1000 48.8000 ;
	    RECT 92.6000 47.8000 93.0000 48.2000 ;
	    RECT 92.6000 47.2000 92.9000 47.8000 ;
	    RECT 90.2000 46.8000 90.6000 47.2000 ;
	    RECT 91.0000 46.8000 91.4000 47.2000 ;
	    RECT 91.8000 46.8000 92.2000 47.2000 ;
	    RECT 92.6000 46.8000 93.0000 47.2000 ;
	    RECT 91.0000 46.2000 91.3000 46.8000 ;
	    RECT 93.4000 46.2000 93.7000 51.8000 ;
	    RECT 94.2000 50.8000 94.6000 51.2000 ;
	    RECT 94.2000 49.2000 94.5000 50.8000 ;
	    RECT 96.6000 49.2000 96.9000 51.8000 ;
	    RECT 101.4000 50.1000 101.7000 51.8000 ;
	    RECT 101.4000 49.8000 102.5000 50.1000 ;
	    RECT 94.2000 48.8000 94.6000 49.2000 ;
	    RECT 96.6000 48.8000 97.0000 49.2000 ;
	    RECT 101.4000 48.8000 101.8000 49.2000 ;
	    RECT 95.0000 48.1000 95.4000 48.2000 ;
	    RECT 95.8000 48.1000 96.2000 48.2000 ;
	    RECT 95.0000 47.8000 96.2000 48.1000 ;
	    RECT 98.2000 48.1000 98.6000 48.2000 ;
	    RECT 99.0000 48.1000 99.4000 48.2000 ;
	    RECT 98.2000 47.8000 99.4000 48.1000 ;
	    RECT 101.4000 47.2000 101.7000 48.8000 ;
	    RECT 96.6000 47.1000 97.0000 47.2000 ;
	    RECT 98.2000 47.1000 98.6000 47.2000 ;
	    RECT 96.6000 46.8000 98.6000 47.1000 ;
	    RECT 101.4000 46.8000 101.8000 47.2000 ;
	    RECT 91.0000 45.8000 91.4000 46.2000 ;
	    RECT 91.8000 46.1000 92.2000 46.2000 ;
	    RECT 92.6000 46.1000 93.0000 46.2000 ;
	    RECT 91.8000 45.8000 93.0000 46.1000 ;
	    RECT 93.4000 45.8000 93.8000 46.2000 ;
	    RECT 95.8000 45.8000 96.2000 46.2000 ;
	    RECT 95.8000 45.2000 96.1000 45.8000 ;
	    RECT 87.0000 44.8000 87.4000 45.2000 ;
	    RECT 89.4000 44.8000 89.8000 45.2000 ;
	    RECT 95.8000 44.8000 96.2000 45.2000 ;
	    RECT 87.0000 39.2000 87.3000 44.8000 ;
	    RECT 99.0000 43.8000 99.4000 44.2000 ;
	    RECT 98.2000 41.8000 98.6000 42.2000 ;
	    RECT 83.8000 38.8000 84.2000 39.2000 ;
	    RECT 87.0000 38.8000 87.4000 39.2000 ;
	    RECT 83.0000 37.8000 83.4000 38.2000 ;
	    RECT 86.2000 37.8000 86.6000 38.2000 ;
	    RECT 83.0000 37.2000 83.3000 37.8000 ;
	    RECT 86.2000 37.2000 86.5000 37.8000 ;
	    RECT 98.2000 37.2000 98.5000 41.8000 ;
	    RECT 83.0000 36.8000 83.4000 37.2000 ;
	    RECT 86.2000 36.8000 86.6000 37.2000 ;
	    RECT 98.2000 36.8000 98.6000 37.2000 ;
	    RECT 85.4000 35.8000 85.8000 36.2000 ;
	    RECT 85.4000 35.2000 85.7000 35.8000 ;
	    RECT 99.0000 35.2000 99.3000 43.8000 ;
	    RECT 101.4000 36.1000 101.8000 36.2000 ;
	    RECT 102.2000 36.1000 102.5000 49.8000 ;
	    RECT 103.0000 46.8000 103.4000 47.2000 ;
	    RECT 103.0000 46.2000 103.3000 46.8000 ;
	    RECT 103.0000 45.8000 103.4000 46.2000 ;
	    RECT 101.4000 35.8000 102.5000 36.1000 ;
	    RECT 81.4000 34.8000 81.8000 35.2000 ;
	    RECT 82.2000 34.8000 82.6000 35.2000 ;
	    RECT 84.6000 34.8000 85.0000 35.2000 ;
	    RECT 85.4000 34.8000 85.8000 35.2000 ;
	    RECT 91.0000 34.8000 91.4000 35.2000 ;
	    RECT 95.0000 34.8000 95.4000 35.2000 ;
	    RECT 97.4000 34.8000 97.8000 35.2000 ;
	    RECT 99.0000 34.8000 99.4000 35.2000 ;
	    RECT 99.8000 34.8000 100.2000 35.2000 ;
	    RECT 101.4000 34.8000 101.8000 35.2000 ;
	    RECT 103.0000 35.1000 103.4000 35.2000 ;
	    RECT 103.8000 35.1000 104.1000 51.8000 ;
	    RECT 105.4000 47.2000 105.7000 51.8000 ;
	    RECT 105.4000 46.8000 105.8000 47.2000 ;
	    RECT 105.4000 45.8000 105.8000 46.2000 ;
	    RECT 105.4000 45.2000 105.7000 45.8000 ;
	    RECT 105.4000 44.8000 105.8000 45.2000 ;
	    RECT 104.6000 43.8000 105.0000 44.2000 ;
	    RECT 104.6000 39.2000 104.9000 43.8000 ;
	    RECT 105.4000 42.8000 105.8000 43.2000 ;
	    RECT 104.6000 38.8000 105.0000 39.2000 ;
	    RECT 103.0000 34.8000 104.1000 35.1000 ;
	    RECT 81.4000 29.1000 81.7000 34.8000 ;
	    RECT 84.6000 29.2000 84.9000 34.8000 ;
	    RECT 91.0000 31.2000 91.3000 34.8000 ;
	    RECT 95.0000 33.2000 95.3000 34.8000 ;
	    RECT 96.6000 33.8000 97.0000 34.2000 ;
	    RECT 92.6000 33.1000 93.0000 33.2000 ;
	    RECT 93.4000 33.1000 93.8000 33.2000 ;
	    RECT 92.6000 32.8000 93.8000 33.1000 ;
	    RECT 95.0000 32.8000 95.4000 33.2000 ;
	    RECT 95.0000 32.2000 95.3000 32.8000 ;
	    RECT 91.8000 31.8000 92.2000 32.2000 ;
	    RECT 95.0000 31.8000 95.4000 32.2000 ;
	    RECT 91.0000 30.8000 91.4000 31.2000 ;
	    RECT 82.2000 29.1000 82.6000 29.2000 ;
	    RECT 78.2000 25.8000 78.6000 26.2000 ;
	    RECT 78.2000 25.2000 78.5000 25.8000 ;
	    RECT 78.2000 24.8000 78.6000 25.2000 ;
	    RECT 78.2000 23.2000 78.5000 24.8000 ;
	    RECT 78.2000 22.8000 78.6000 23.2000 ;
	    RECT 79.8000 23.1000 80.2000 28.9000 ;
	    RECT 81.4000 28.8000 82.6000 29.1000 ;
	    RECT 83.0000 29.1000 83.4000 29.2000 ;
	    RECT 83.8000 29.1000 84.2000 29.2000 ;
	    RECT 83.0000 28.8000 84.2000 29.1000 ;
	    RECT 84.6000 28.8000 85.0000 29.2000 ;
	    RECT 91.8000 29.1000 92.1000 31.8000 ;
	    RECT 85.4000 23.1000 85.8000 28.9000 ;
	    RECT 86.2000 25.8000 86.6000 26.2000 ;
	    RECT 89.4000 25.9000 89.8000 26.3000 ;
	    RECT 86.2000 25.2000 86.5000 25.8000 ;
	    RECT 89.4000 25.2000 89.7000 25.9000 ;
	    RECT 86.2000 24.8000 86.6000 25.2000 ;
	    RECT 89.4000 24.8000 89.8000 25.2000 ;
	    RECT 90.2000 23.1000 90.6000 28.9000 ;
	    RECT 91.8000 28.8000 92.9000 29.1000 ;
	    RECT 92.6000 28.2000 92.9000 28.8000 ;
	    RECT 91.8000 25.1000 92.2000 27.9000 ;
	    RECT 92.6000 27.8000 93.0000 28.2000 ;
	    RECT 96.6000 27.2000 96.9000 33.8000 ;
	    RECT 97.4000 33.2000 97.7000 34.8000 ;
	    RECT 98.2000 33.8000 98.6000 34.2000 ;
	    RECT 99.0000 33.8000 99.4000 34.2000 ;
	    RECT 97.4000 32.8000 97.8000 33.2000 ;
	    RECT 97.4000 28.2000 97.7000 32.8000 ;
	    RECT 98.2000 31.2000 98.5000 33.8000 ;
	    RECT 99.0000 33.2000 99.3000 33.8000 ;
	    RECT 99.0000 32.8000 99.4000 33.2000 ;
	    RECT 99.0000 31.8000 99.4000 32.2000 ;
	    RECT 98.2000 30.8000 98.6000 31.2000 ;
	    RECT 99.0000 29.2000 99.3000 31.8000 ;
	    RECT 99.0000 28.8000 99.4000 29.2000 ;
	    RECT 99.8000 28.2000 100.1000 34.8000 ;
	    RECT 101.4000 34.2000 101.7000 34.8000 ;
	    RECT 101.4000 33.8000 101.8000 34.2000 ;
	    RECT 102.2000 33.8000 102.6000 34.2000 ;
	    RECT 102.2000 32.2000 102.5000 33.8000 ;
	    RECT 103.8000 33.2000 104.1000 34.8000 ;
	    RECT 103.8000 32.8000 104.2000 33.2000 ;
	    RECT 102.2000 31.8000 102.6000 32.2000 ;
	    RECT 103.8000 31.8000 104.2000 32.2000 ;
	    RECT 101.4000 29.1000 101.8000 29.2000 ;
	    RECT 102.2000 29.1000 102.6000 29.2000 ;
	    RECT 101.4000 28.8000 102.6000 29.1000 ;
	    RECT 97.4000 27.8000 97.8000 28.2000 ;
	    RECT 99.8000 27.8000 100.2000 28.2000 ;
	    RECT 99.8000 27.2000 100.1000 27.8000 ;
	    RECT 103.8000 27.2000 104.1000 31.8000 ;
	    RECT 105.4000 31.2000 105.7000 42.8000 ;
	    RECT 106.2000 36.2000 106.5000 56.8000 ;
	    RECT 108.6000 55.2000 108.9000 57.8000 ;
	    RECT 108.6000 54.8000 109.0000 55.2000 ;
	    RECT 110.2000 53.8000 110.6000 54.2000 ;
	    RECT 107.8000 48.1000 108.2000 48.2000 ;
	    RECT 108.6000 48.1000 109.0000 48.2000 ;
	    RECT 107.8000 47.8000 109.0000 48.1000 ;
	    RECT 108.6000 45.1000 109.0000 45.2000 ;
	    RECT 109.4000 45.1000 109.8000 45.2000 ;
	    RECT 108.6000 44.8000 109.8000 45.1000 ;
	    RECT 109.4000 41.8000 109.8000 42.2000 ;
	    RECT 106.2000 35.8000 106.6000 36.2000 ;
	    RECT 107.0000 33.1000 107.4000 35.9000 ;
	    RECT 106.2000 31.8000 106.6000 32.2000 ;
	    RECT 108.6000 32.1000 109.0000 37.9000 ;
	    RECT 109.4000 35.1000 109.7000 41.8000 ;
	    RECT 109.4000 34.7000 109.8000 35.1000 ;
	    RECT 110.2000 32.2000 110.5000 53.8000 ;
	    RECT 111.8000 52.1000 112.2000 57.9000 ;
	    RECT 112.6000 57.8000 113.0000 58.2000 ;
	    RECT 115.0000 55.0000 115.4000 55.1000 ;
	    RECT 115.8000 55.0000 116.2000 55.1000 ;
	    RECT 115.0000 54.7000 116.2000 55.0000 ;
	    RECT 112.6000 53.8000 113.0000 54.2000 ;
	    RECT 111.0000 46.1000 111.4000 46.2000 ;
	    RECT 111.8000 46.1000 112.2000 46.2000 ;
	    RECT 111.0000 45.8000 112.2000 46.1000 ;
	    RECT 111.0000 44.8000 111.4000 45.2000 ;
	    RECT 111.0000 44.2000 111.3000 44.8000 ;
	    RECT 111.0000 43.8000 111.4000 44.2000 ;
	    RECT 112.6000 35.2000 112.9000 53.8000 ;
	    RECT 116.6000 52.1000 117.0000 57.9000 ;
	    RECT 117.4000 53.8000 117.8000 54.2000 ;
	    RECT 115.8000 43.1000 116.2000 48.9000 ;
	    RECT 117.4000 47.2000 117.7000 53.8000 ;
	    RECT 118.2000 53.1000 118.6000 55.9000 ;
	    RECT 119.0000 53.2000 119.3000 66.8000 ;
	    RECT 120.6000 66.1000 121.0000 66.2000 ;
	    RECT 121.4000 66.1000 121.8000 66.2000 ;
	    RECT 120.6000 65.8000 121.8000 66.1000 ;
	    RECT 122.2000 63.8000 122.6000 64.2000 ;
	    RECT 122.2000 59.2000 122.5000 63.8000 ;
	    RECT 122.2000 58.8000 122.6000 59.2000 ;
	    RECT 123.0000 58.2000 123.3000 69.8000 ;
	    RECT 125.4000 69.2000 125.7000 70.8000 ;
	    RECT 125.4000 68.8000 125.8000 69.2000 ;
	    RECT 127.8000 68.2000 128.1000 71.8000 ;
	    RECT 125.4000 67.8000 125.8000 68.2000 ;
	    RECT 127.8000 67.8000 128.2000 68.2000 ;
	    RECT 123.8000 67.1000 124.2000 67.2000 ;
	    RECT 124.6000 67.1000 125.0000 67.2000 ;
	    RECT 123.8000 66.8000 125.0000 67.1000 ;
	    RECT 123.8000 65.8000 124.2000 66.2000 ;
	    RECT 123.8000 64.2000 124.1000 65.8000 ;
	    RECT 125.4000 65.2000 125.7000 67.8000 ;
	    RECT 127.0000 67.1000 127.4000 67.2000 ;
	    RECT 127.8000 67.1000 128.2000 67.2000 ;
	    RECT 127.0000 66.8000 128.2000 67.1000 ;
	    RECT 127.0000 65.8000 127.4000 66.2000 ;
	    RECT 127.8000 65.8000 128.2000 66.2000 ;
	    RECT 125.4000 64.8000 125.8000 65.2000 ;
	    RECT 127.0000 64.2000 127.3000 65.8000 ;
	    RECT 123.8000 63.8000 124.2000 64.2000 ;
	    RECT 127.0000 63.8000 127.4000 64.2000 ;
	    RECT 123.8000 61.8000 124.2000 62.2000 ;
	    RECT 123.0000 57.8000 123.4000 58.2000 ;
	    RECT 123.0000 57.2000 123.3000 57.8000 ;
	    RECT 123.8000 57.2000 124.1000 61.8000 ;
	    RECT 127.8000 61.2000 128.1000 65.8000 ;
	    RECT 127.8000 60.8000 128.2000 61.2000 ;
	    RECT 120.6000 56.8000 121.0000 57.2000 ;
	    RECT 123.0000 56.8000 123.4000 57.2000 ;
	    RECT 123.8000 56.8000 124.2000 57.2000 ;
	    RECT 127.0000 57.1000 127.4000 57.2000 ;
	    RECT 127.8000 57.1000 128.2000 57.2000 ;
	    RECT 127.0000 56.8000 128.2000 57.1000 ;
	    RECT 119.8000 54.8000 120.2000 55.2000 ;
	    RECT 119.8000 54.2000 120.1000 54.8000 ;
	    RECT 120.6000 54.2000 120.9000 56.8000 ;
	    RECT 123.0000 55.8000 123.4000 56.2000 ;
	    RECT 123.0000 55.2000 123.3000 55.8000 ;
	    RECT 128.6000 55.2000 128.9000 71.8000 ;
	    RECT 135.0000 71.2000 135.3000 74.7000 ;
	    RECT 135.8000 72.1000 136.2000 77.9000 ;
	    RECT 136.6000 74.8000 137.0000 75.2000 ;
	    RECT 136.6000 74.2000 136.9000 74.8000 ;
	    RECT 136.6000 73.8000 137.0000 74.2000 ;
	    RECT 137.4000 73.1000 137.8000 75.9000 ;
	    RECT 143.8000 75.8000 144.2000 76.2000 ;
	    RECT 138.2000 74.8000 138.6000 75.2000 ;
	    RECT 135.0000 70.8000 135.4000 71.2000 ;
	    RECT 138.2000 69.2000 138.5000 74.8000 ;
	    RECT 143.8000 73.2000 144.1000 75.8000 ;
	    RECT 155.8000 75.2000 156.1000 86.8000 ;
	    RECT 159.8000 86.2000 160.1000 88.8000 ;
	    RECT 164.6000 88.2000 164.9000 91.8000 ;
	    RECT 165.4000 88.8000 165.8000 89.2000 ;
	    RECT 162.2000 88.1000 162.6000 88.2000 ;
	    RECT 163.0000 88.1000 163.4000 88.2000 ;
	    RECT 162.2000 87.8000 163.4000 88.1000 ;
	    RECT 164.6000 87.8000 165.0000 88.2000 ;
	    RECT 160.6000 87.1000 161.0000 87.2000 ;
	    RECT 161.4000 87.1000 161.8000 87.2000 ;
	    RECT 160.6000 86.8000 161.8000 87.1000 ;
	    RECT 164.6000 86.8000 165.0000 87.2000 ;
	    RECT 159.8000 85.8000 160.2000 86.2000 ;
	    RECT 160.6000 86.1000 161.0000 86.2000 ;
	    RECT 161.4000 86.1000 161.8000 86.2000 ;
	    RECT 160.6000 85.8000 161.8000 86.1000 ;
	    RECT 158.2000 85.1000 158.6000 85.2000 ;
	    RECT 159.0000 85.1000 159.4000 85.2000 ;
	    RECT 158.2000 84.8000 159.4000 85.1000 ;
	    RECT 161.4000 75.8000 161.8000 76.2000 ;
	    RECT 161.4000 75.2000 161.7000 75.8000 ;
	    RECT 144.6000 74.8000 145.0000 75.2000 ;
	    RECT 155.8000 74.8000 156.2000 75.2000 ;
	    RECT 160.6000 74.8000 161.0000 75.2000 ;
	    RECT 161.4000 74.8000 161.8000 75.2000 ;
	    RECT 162.2000 74.8000 162.6000 75.2000 ;
	    RECT 163.8000 74.8000 164.2000 75.2000 ;
	    RECT 144.6000 74.2000 144.9000 74.8000 ;
	    RECT 160.6000 74.2000 160.9000 74.8000 ;
	    RECT 144.6000 73.8000 145.0000 74.2000 ;
	    RECT 160.6000 73.8000 161.0000 74.2000 ;
	    RECT 143.8000 72.8000 144.2000 73.2000 ;
	    RECT 139.0000 71.8000 139.4000 72.2000 ;
	    RECT 139.8000 71.8000 140.2000 72.2000 ;
	    RECT 152.6000 71.8000 153.0000 72.2000 ;
	    RECT 135.0000 69.1000 135.4000 69.2000 ;
	    RECT 135.8000 69.1000 136.2000 69.2000 ;
	    RECT 135.0000 68.8000 136.2000 69.1000 ;
	    RECT 138.2000 68.8000 138.6000 69.2000 ;
	    RECT 133.4000 67.1000 133.8000 67.2000 ;
	    RECT 134.2000 67.1000 134.6000 67.2000 ;
	    RECT 133.4000 66.8000 134.6000 67.1000 ;
	    RECT 135.0000 66.8000 135.4000 67.2000 ;
	    RECT 131.8000 65.8000 132.2000 66.2000 ;
	    RECT 129.4000 63.8000 129.8000 64.2000 ;
	    RECT 121.4000 54.8000 121.8000 55.2000 ;
	    RECT 122.2000 54.8000 122.6000 55.2000 ;
	    RECT 123.0000 54.8000 123.4000 55.2000 ;
	    RECT 123.8000 54.8000 124.2000 55.2000 ;
	    RECT 125.4000 54.8000 125.8000 55.2000 ;
	    RECT 127.0000 54.8000 127.4000 55.2000 ;
	    RECT 128.6000 54.8000 129.0000 55.2000 ;
	    RECT 121.4000 54.2000 121.7000 54.8000 ;
	    RECT 119.8000 53.8000 120.2000 54.2000 ;
	    RECT 120.6000 53.8000 121.0000 54.2000 ;
	    RECT 121.4000 53.8000 121.8000 54.2000 ;
	    RECT 119.0000 52.8000 119.4000 53.2000 ;
	    RECT 119.0000 48.2000 119.3000 52.8000 ;
	    RECT 122.2000 49.2000 122.5000 54.8000 ;
	    RECT 123.8000 54.2000 124.1000 54.8000 ;
	    RECT 125.4000 54.2000 125.7000 54.8000 ;
	    RECT 127.0000 54.2000 127.3000 54.8000 ;
	    RECT 123.8000 53.8000 124.2000 54.2000 ;
	    RECT 125.4000 53.8000 125.8000 54.2000 ;
	    RECT 127.0000 53.8000 127.4000 54.2000 ;
	    RECT 127.8000 54.1000 128.2000 54.2000 ;
	    RECT 128.6000 54.1000 129.0000 54.2000 ;
	    RECT 127.8000 53.8000 129.0000 54.1000 ;
	    RECT 127.0000 53.1000 127.4000 53.2000 ;
	    RECT 127.8000 53.1000 128.2000 53.2000 ;
	    RECT 127.0000 52.8000 128.2000 53.1000 ;
	    RECT 119.0000 47.8000 119.4000 48.2000 ;
	    RECT 117.4000 46.8000 117.8000 47.2000 ;
	    RECT 119.8000 46.8000 120.2000 47.2000 ;
	    RECT 119.8000 46.3000 120.1000 46.8000 ;
	    RECT 119.8000 45.9000 120.2000 46.3000 ;
	    RECT 120.6000 43.1000 121.0000 48.9000 ;
	    RECT 122.2000 48.8000 122.6000 49.2000 ;
	    RECT 121.4000 46.8000 121.8000 47.2000 ;
	    RECT 121.4000 44.2000 121.7000 46.8000 ;
	    RECT 122.2000 45.1000 122.6000 47.9000 ;
	    RECT 123.8000 47.8000 124.2000 48.2000 ;
	    RECT 127.0000 48.1000 127.4000 48.2000 ;
	    RECT 127.8000 48.1000 128.2000 48.2000 ;
	    RECT 127.0000 47.8000 128.2000 48.1000 ;
	    RECT 123.0000 46.8000 123.4000 47.2000 ;
	    RECT 121.4000 43.8000 121.8000 44.2000 ;
	    RECT 123.0000 43.2000 123.3000 46.8000 ;
	    RECT 123.0000 42.8000 123.4000 43.2000 ;
	    RECT 123.8000 39.2000 124.1000 47.8000 ;
	    RECT 127.8000 46.8000 128.2000 47.2000 ;
	    RECT 126.2000 46.1000 126.6000 46.2000 ;
	    RECT 127.0000 46.1000 127.4000 46.2000 ;
	    RECT 126.2000 45.8000 127.4000 46.1000 ;
	    RECT 127.8000 45.2000 128.1000 46.8000 ;
	    RECT 128.6000 46.2000 128.9000 53.8000 ;
	    RECT 129.4000 53.2000 129.7000 63.8000 ;
	    RECT 130.2000 61.8000 130.6000 62.2000 ;
	    RECT 130.2000 56.2000 130.5000 61.8000 ;
	    RECT 131.8000 60.2000 132.1000 65.8000 ;
	    RECT 135.0000 62.2000 135.3000 66.8000 ;
	    RECT 139.0000 65.2000 139.3000 71.8000 ;
	    RECT 139.8000 69.2000 140.1000 71.8000 ;
	    RECT 143.8000 70.8000 144.2000 71.2000 ;
	    RECT 143.8000 69.2000 144.1000 70.8000 ;
	    RECT 139.8000 68.8000 140.2000 69.2000 ;
	    RECT 143.8000 68.8000 144.2000 69.2000 ;
	    RECT 144.6000 68.8000 145.0000 69.2000 ;
	    RECT 151.0000 68.8000 151.4000 69.2000 ;
	    RECT 144.6000 68.2000 144.9000 68.8000 ;
	    RECT 151.0000 68.2000 151.3000 68.8000 ;
	    RECT 139.8000 67.8000 142.5000 68.1000 ;
	    RECT 144.6000 67.8000 145.0000 68.2000 ;
	    RECT 151.0000 67.8000 151.4000 68.2000 ;
	    RECT 139.8000 67.2000 140.1000 67.8000 ;
	    RECT 142.2000 67.2000 142.5000 67.8000 ;
	    RECT 152.6000 67.2000 152.9000 71.8000 ;
	    RECT 139.8000 66.8000 140.2000 67.2000 ;
	    RECT 140.6000 67.1000 141.0000 67.2000 ;
	    RECT 141.4000 67.1000 141.8000 67.2000 ;
	    RECT 140.6000 66.8000 141.8000 67.1000 ;
	    RECT 142.2000 66.8000 142.6000 67.2000 ;
	    RECT 144.6000 67.1000 145.0000 67.2000 ;
	    RECT 145.4000 67.1000 145.8000 67.2000 ;
	    RECT 144.6000 66.8000 145.8000 67.1000 ;
	    RECT 151.0000 66.8000 151.4000 67.2000 ;
	    RECT 152.6000 66.8000 153.0000 67.2000 ;
	    RECT 151.0000 66.2000 151.3000 66.8000 ;
	    RECT 139.8000 66.1000 140.2000 66.2000 ;
	    RECT 140.6000 66.1000 141.0000 66.2000 ;
	    RECT 139.8000 65.8000 141.0000 66.1000 ;
	    RECT 142.2000 65.8000 142.6000 66.2000 ;
	    RECT 145.4000 66.1000 145.8000 66.2000 ;
	    RECT 146.2000 66.1000 146.6000 66.2000 ;
	    RECT 145.4000 65.8000 146.6000 66.1000 ;
	    RECT 148.6000 65.8000 149.0000 66.2000 ;
	    RECT 151.0000 65.8000 151.4000 66.2000 ;
	    RECT 139.0000 64.8000 139.4000 65.2000 ;
	    RECT 135.0000 61.8000 135.4000 62.2000 ;
	    RECT 131.8000 59.8000 132.2000 60.2000 ;
	    RECT 142.2000 59.2000 142.5000 65.8000 ;
	    RECT 147.8000 64.8000 148.2000 65.2000 ;
	    RECT 147.8000 64.2000 148.1000 64.8000 ;
	    RECT 147.8000 63.8000 148.2000 64.2000 ;
	    RECT 148.6000 59.2000 148.9000 65.8000 ;
	    RECT 151.0000 64.1000 151.4000 64.2000 ;
	    RECT 151.8000 64.1000 152.2000 64.2000 ;
	    RECT 151.0000 63.8000 152.2000 64.1000 ;
	    RECT 154.2000 63.1000 154.6000 68.9000 ;
	    RECT 155.0000 66.8000 155.4000 67.2000 ;
	    RECT 155.0000 66.2000 155.3000 66.8000 ;
	    RECT 155.0000 65.8000 155.4000 66.2000 ;
	    RECT 155.8000 65.8000 156.2000 66.2000 ;
	    RECT 155.8000 65.2000 156.1000 65.8000 ;
	    RECT 155.8000 64.8000 156.2000 65.2000 ;
	    RECT 159.0000 63.1000 159.4000 68.9000 ;
	    RECT 160.6000 65.1000 161.0000 67.9000 ;
	    RECT 162.2000 67.2000 162.5000 74.8000 ;
	    RECT 163.8000 74.2000 164.1000 74.8000 ;
	    RECT 164.6000 74.2000 164.9000 86.8000 ;
	    RECT 165.4000 86.2000 165.7000 88.8000 ;
	    RECT 166.2000 88.1000 166.6000 88.2000 ;
	    RECT 167.0000 88.1000 167.4000 88.2000 ;
	    RECT 166.2000 87.8000 167.4000 88.1000 ;
	    RECT 165.4000 85.8000 165.8000 86.2000 ;
	    RECT 167.0000 76.2000 167.3000 87.8000 ;
	    RECT 167.0000 75.8000 167.4000 76.2000 ;
	    RECT 163.8000 73.8000 164.2000 74.2000 ;
	    RECT 164.6000 73.8000 165.0000 74.2000 ;
	    RECT 166.2000 73.1000 166.6000 73.2000 ;
	    RECT 167.0000 73.1000 167.4000 73.2000 ;
	    RECT 167.8000 73.1000 168.2000 75.9000 ;
	    RECT 168.6000 75.2000 168.9000 94.8000 ;
	    RECT 169.4000 94.1000 169.8000 94.2000 ;
	    RECT 170.2000 94.1000 170.6000 94.2000 ;
	    RECT 169.4000 93.8000 170.6000 94.1000 ;
	    RECT 169.4000 91.8000 169.8000 92.2000 ;
	    RECT 169.4000 89.2000 169.7000 91.8000 ;
	    RECT 169.4000 88.8000 169.8000 89.2000 ;
	    RECT 171.0000 87.1000 171.3000 94.8000 ;
	    RECT 171.8000 94.2000 172.1000 94.8000 ;
	    RECT 171.8000 93.8000 172.2000 94.2000 ;
	    RECT 172.6000 93.1000 173.0000 93.2000 ;
	    RECT 173.4000 93.1000 173.8000 93.2000 ;
	    RECT 174.2000 93.1000 174.6000 95.9000 ;
	    RECT 175.0000 94.2000 175.3000 96.8000 ;
	    RECT 175.0000 93.8000 175.4000 94.2000 ;
	    RECT 172.6000 92.8000 173.8000 93.1000 ;
	    RECT 172.6000 91.8000 173.0000 92.2000 ;
	    RECT 172.6000 90.2000 172.9000 91.8000 ;
	    RECT 172.6000 89.8000 173.0000 90.2000 ;
	    RECT 171.8000 87.8000 172.2000 88.2000 ;
	    RECT 171.8000 87.2000 172.1000 87.8000 ;
	    RECT 171.8000 87.1000 172.2000 87.2000 ;
	    RECT 171.0000 86.8000 172.2000 87.1000 ;
	    RECT 170.2000 85.8000 170.6000 86.2000 ;
	    RECT 170.2000 85.2000 170.5000 85.8000 ;
	    RECT 170.2000 84.8000 170.6000 85.2000 ;
	    RECT 172.6000 85.1000 173.0000 87.9000 ;
	    RECT 173.4000 86.8000 173.8000 87.2000 ;
	    RECT 168.6000 74.8000 169.0000 75.2000 ;
	    RECT 166.2000 72.8000 167.4000 73.1000 ;
	    RECT 163.0000 71.8000 163.4000 72.2000 ;
	    RECT 164.6000 71.8000 165.0000 72.2000 ;
	    RECT 161.4000 66.8000 161.8000 67.2000 ;
	    RECT 162.2000 66.8000 162.6000 67.2000 ;
	    RECT 159.0000 61.8000 159.4000 62.2000 ;
	    RECT 161.4000 62.1000 161.7000 66.8000 ;
	    RECT 161.4000 61.8000 162.5000 62.1000 ;
	    RECT 159.0000 59.2000 159.3000 61.8000 ;
	    RECT 142.2000 58.8000 142.6000 59.2000 ;
	    RECT 143.8000 59.1000 144.2000 59.2000 ;
	    RECT 144.6000 59.1000 145.0000 59.2000 ;
	    RECT 143.8000 58.8000 145.0000 59.1000 ;
	    RECT 148.6000 58.8000 149.0000 59.2000 ;
	    RECT 159.0000 58.8000 159.4000 59.2000 ;
	    RECT 130.2000 55.8000 130.6000 56.2000 ;
	    RECT 131.0000 55.8000 131.4000 56.2000 ;
	    RECT 129.4000 52.8000 129.8000 53.2000 ;
	    RECT 129.4000 47.2000 129.7000 52.8000 ;
	    RECT 131.0000 47.2000 131.3000 55.8000 ;
	    RECT 131.8000 55.1000 132.2000 55.2000 ;
	    RECT 132.6000 55.1000 133.0000 55.2000 ;
	    RECT 131.8000 54.8000 133.0000 55.1000 ;
	    RECT 134.2000 54.8000 134.6000 55.2000 ;
	    RECT 134.2000 54.2000 134.5000 54.8000 ;
	    RECT 131.8000 53.8000 132.2000 54.2000 ;
	    RECT 132.6000 54.1000 133.0000 54.2000 ;
	    RECT 133.4000 54.1000 133.8000 54.2000 ;
	    RECT 132.6000 53.8000 133.8000 54.1000 ;
	    RECT 134.2000 53.8000 134.6000 54.2000 ;
	    RECT 131.8000 53.2000 132.1000 53.8000 ;
	    RECT 131.8000 52.8000 132.2000 53.2000 ;
	    RECT 133.4000 53.1000 133.8000 53.2000 ;
	    RECT 134.2000 53.1000 134.6000 53.2000 ;
	    RECT 135.0000 53.1000 135.4000 55.9000 ;
	    RECT 133.4000 52.8000 134.6000 53.1000 ;
	    RECT 136.6000 52.1000 137.0000 57.9000 ;
	    RECT 137.4000 55.0000 137.8000 55.1000 ;
	    RECT 138.2000 55.0000 138.6000 55.1000 ;
	    RECT 137.4000 54.7000 138.6000 55.0000 ;
	    RECT 140.6000 54.8000 141.0000 55.2000 ;
	    RECT 140.6000 54.2000 140.9000 54.8000 ;
	    RECT 140.6000 53.8000 141.0000 54.2000 ;
	    RECT 141.4000 52.1000 141.8000 57.9000 ;
	    RECT 145.4000 57.8000 145.8000 58.2000 ;
	    RECT 145.4000 57.2000 145.7000 57.8000 ;
	    RECT 143.8000 57.1000 144.2000 57.2000 ;
	    RECT 144.6000 57.1000 145.0000 57.2000 ;
	    RECT 143.8000 56.8000 145.0000 57.1000 ;
	    RECT 145.4000 56.8000 145.8000 57.2000 ;
	    RECT 147.8000 56.8000 148.2000 57.2000 ;
	    RECT 147.8000 56.2000 148.1000 56.8000 ;
	    RECT 159.0000 56.2000 159.3000 58.8000 ;
	    RECT 146.2000 55.8000 146.6000 56.2000 ;
	    RECT 147.0000 55.8000 147.4000 56.2000 ;
	    RECT 147.8000 55.8000 148.2000 56.2000 ;
	    RECT 148.6000 55.8000 149.0000 56.2000 ;
	    RECT 154.2000 55.8000 154.6000 56.2000 ;
	    RECT 159.0000 55.8000 159.4000 56.2000 ;
	    RECT 146.2000 55.2000 146.5000 55.8000 ;
	    RECT 143.8000 54.8000 144.2000 55.2000 ;
	    RECT 146.2000 54.8000 146.6000 55.2000 ;
	    RECT 129.4000 46.8000 129.8000 47.2000 ;
	    RECT 130.2000 47.1000 130.6000 47.2000 ;
	    RECT 131.0000 47.1000 131.4000 47.2000 ;
	    RECT 130.2000 46.8000 131.4000 47.1000 ;
	    RECT 128.6000 45.8000 129.0000 46.2000 ;
	    RECT 130.2000 45.8000 130.6000 46.2000 ;
	    RECT 131.0000 46.1000 131.4000 46.2000 ;
	    RECT 131.8000 46.1000 132.2000 46.2000 ;
	    RECT 131.0000 45.8000 132.2000 46.1000 ;
	    RECT 133.4000 45.8000 133.8000 46.2000 ;
	    RECT 130.2000 45.2000 130.5000 45.8000 ;
	    RECT 133.4000 45.2000 133.7000 45.8000 ;
	    RECT 124.6000 45.1000 125.0000 45.2000 ;
	    RECT 125.4000 45.1000 125.8000 45.2000 ;
	    RECT 124.6000 44.8000 125.8000 45.1000 ;
	    RECT 127.8000 44.8000 128.2000 45.2000 ;
	    RECT 130.2000 44.8000 130.6000 45.2000 ;
	    RECT 133.4000 44.8000 133.8000 45.2000 ;
	    RECT 135.0000 44.8000 135.4000 45.2000 ;
	    RECT 141.4000 45.1000 141.8000 47.9000 ;
	    RECT 124.6000 42.8000 125.0000 43.2000 ;
	    RECT 124.6000 39.2000 124.9000 42.8000 ;
	    RECT 115.0000 39.1000 115.4000 39.2000 ;
	    RECT 115.8000 39.1000 116.2000 39.2000 ;
	    RECT 115.0000 38.8000 116.2000 39.1000 ;
	    RECT 123.8000 38.8000 124.2000 39.2000 ;
	    RECT 124.6000 38.8000 125.0000 39.2000 ;
	    RECT 112.6000 34.8000 113.0000 35.2000 ;
	    RECT 110.2000 31.8000 110.6000 32.2000 ;
	    RECT 113.4000 32.1000 113.8000 37.9000 ;
	    RECT 119.0000 37.8000 119.4000 38.2000 ;
	    RECT 119.0000 36.2000 119.3000 37.8000 ;
	    RECT 123.8000 37.2000 124.1000 38.8000 ;
	    RECT 123.8000 36.8000 124.2000 37.2000 ;
	    RECT 119.0000 35.8000 119.4000 36.2000 ;
	    RECT 120.6000 35.8000 121.0000 36.2000 ;
	    RECT 123.8000 36.1000 124.2000 36.2000 ;
	    RECT 124.6000 36.1000 125.0000 36.2000 ;
	    RECT 123.8000 35.8000 125.0000 36.1000 ;
	    RECT 117.4000 34.8000 117.8000 35.2000 ;
	    RECT 119.0000 35.1000 119.4000 35.2000 ;
	    RECT 119.8000 35.1000 120.2000 35.2000 ;
	    RECT 119.0000 34.8000 120.2000 35.1000 ;
	    RECT 116.6000 33.8000 117.0000 34.2000 ;
	    RECT 116.6000 33.2000 116.9000 33.8000 ;
	    RECT 116.6000 32.8000 117.0000 33.2000 ;
	    RECT 105.4000 30.8000 105.8000 31.2000 ;
	    RECT 104.6000 27.8000 105.0000 28.2000 ;
	    RECT 104.6000 27.2000 104.9000 27.8000 ;
	    RECT 105.4000 27.2000 105.7000 30.8000 ;
	    RECT 96.6000 26.8000 97.0000 27.2000 ;
	    RECT 98.2000 26.8000 98.6000 27.2000 ;
	    RECT 99.8000 26.8000 100.2000 27.2000 ;
	    RECT 100.6000 26.8000 101.0000 27.2000 ;
	    RECT 103.8000 26.8000 104.2000 27.2000 ;
	    RECT 104.6000 26.8000 105.0000 27.2000 ;
	    RECT 105.4000 26.8000 105.8000 27.2000 ;
	    RECT 95.0000 25.8000 95.4000 26.2000 ;
	    RECT 97.4000 25.8000 97.8000 26.2000 ;
	    RECT 95.0000 25.2000 95.3000 25.8000 ;
	    RECT 93.4000 24.8000 93.8000 25.2000 ;
	    RECT 94.2000 24.8000 94.6000 25.2000 ;
	    RECT 95.0000 24.8000 95.4000 25.2000 ;
	    RECT 93.4000 24.2000 93.7000 24.8000 ;
	    RECT 93.4000 23.8000 93.8000 24.2000 ;
	    RECT 91.8000 22.8000 92.2000 23.2000 ;
	    RECT 78.2000 19.2000 78.5000 22.8000 ;
	    RECT 85.4000 21.8000 85.8000 22.2000 ;
	    RECT 85.4000 19.2000 85.7000 21.8000 ;
	    RECT 89.4000 20.8000 89.8000 21.2000 ;
	    RECT 89.4000 19.2000 89.7000 20.8000 ;
	    RECT 91.8000 19.2000 92.1000 22.8000 ;
	    RECT 94.2000 19.2000 94.5000 24.8000 ;
	    RECT 97.4000 22.2000 97.7000 25.8000 ;
	    RECT 98.2000 23.2000 98.5000 26.8000 ;
	    RECT 98.2000 22.8000 98.6000 23.2000 ;
	    RECT 100.6000 22.2000 100.9000 26.8000 ;
	    RECT 101.4000 25.1000 101.8000 25.2000 ;
	    RECT 102.2000 25.1000 102.6000 25.2000 ;
	    RECT 101.4000 24.8000 102.6000 25.1000 ;
	    RECT 97.4000 21.8000 97.8000 22.2000 ;
	    RECT 100.6000 21.8000 101.0000 22.2000 ;
	    RECT 78.2000 18.8000 78.6000 19.2000 ;
	    RECT 85.4000 18.8000 85.8000 19.2000 ;
	    RECT 89.4000 18.8000 89.8000 19.2000 ;
	    RECT 91.8000 18.8000 92.2000 19.2000 ;
	    RECT 94.2000 18.8000 94.6000 19.2000 ;
	    RECT 82.2000 15.8000 82.6000 16.2000 ;
	    RECT 87.0000 15.8000 87.4000 16.2000 ;
	    RECT 90.2000 16.1000 90.6000 16.2000 ;
	    RECT 91.0000 16.1000 91.4000 16.2000 ;
	    RECT 90.2000 15.8000 91.4000 16.1000 ;
	    RECT 95.8000 15.8000 96.2000 16.2000 ;
	    RECT 78.2000 13.8000 78.6000 14.2000 ;
	    RECT 76.6000 12.8000 77.0000 13.2000 ;
	    RECT 74.2000 11.8000 74.6000 12.2000 ;
	    RECT 75.0000 11.8000 75.4000 12.2000 ;
	    RECT 64.6000 9.8000 65.0000 10.2000 ;
	    RECT 61.4000 8.8000 61.8000 9.2000 ;
	    RECT 63.8000 8.8000 64.2000 9.2000 ;
	    RECT 63.8000 8.2000 64.1000 8.8000 ;
	    RECT 60.6000 7.8000 61.0000 8.2000 ;
	    RECT 63.8000 7.8000 64.2000 8.2000 ;
	    RECT 63.8000 6.2000 64.1000 7.8000 ;
	    RECT 64.6000 7.2000 64.9000 9.8000 ;
	    RECT 74.2000 9.2000 74.5000 11.8000 ;
	    RECT 67.0000 9.1000 67.4000 9.2000 ;
	    RECT 67.8000 9.1000 68.2000 9.2000 ;
	    RECT 67.0000 8.8000 68.2000 9.1000 ;
	    RECT 74.2000 8.8000 74.6000 9.2000 ;
	    RECT 65.4000 7.5000 65.8000 7.9000 ;
	    RECT 68.5000 7.8000 68.9000 7.9000 ;
	    RECT 66.1000 7.5000 68.9000 7.8000 ;
	    RECT 64.6000 6.8000 65.0000 7.2000 ;
	    RECT 65.4000 7.1000 65.7000 7.5000 ;
	    RECT 66.1000 7.4000 66.5000 7.5000 ;
	    RECT 67.8000 7.4000 68.2000 7.5000 ;
	    RECT 65.4000 6.8000 68.2000 7.1000 ;
	    RECT 59.8000 5.8000 60.2000 6.2000 ;
	    RECT 63.8000 5.8000 64.2000 6.2000 ;
	    RECT 54.1000 4.7000 54.5000 5.1000 ;
	    RECT 57.4000 4.7000 57.8000 5.1000 ;
	    RECT 65.4000 5.1000 65.7000 6.8000 ;
	    RECT 67.9000 6.1000 68.2000 6.8000 ;
	    RECT 67.9000 5.7000 68.3000 6.1000 ;
	    RECT 68.6000 5.1000 68.9000 7.5000 ;
	    RECT 71.1000 7.8000 71.5000 7.9000 ;
	    RECT 71.1000 7.5000 73.9000 7.8000 ;
	    RECT 74.2000 7.5000 74.6000 7.9000 ;
	    RECT 69.4000 6.8000 69.8000 7.2000 ;
	    RECT 70.2000 6.8000 70.6000 7.2000 ;
	    RECT 69.4000 6.2000 69.7000 6.8000 ;
	    RECT 70.2000 6.2000 70.5000 6.8000 ;
	    RECT 69.4000 5.8000 69.8000 6.2000 ;
	    RECT 70.2000 5.8000 70.6000 6.2000 ;
	    RECT 65.4000 4.7000 65.8000 5.1000 ;
	    RECT 68.5000 4.7000 68.9000 5.1000 ;
	    RECT 71.1000 5.1000 71.4000 7.5000 ;
	    RECT 71.8000 7.4000 72.2000 7.5000 ;
	    RECT 73.5000 7.4000 73.9000 7.5000 ;
	    RECT 74.3000 7.1000 74.6000 7.5000 ;
	    RECT 71.8000 6.8000 74.6000 7.1000 ;
	    RECT 75.0000 7.8000 75.4000 8.2000 ;
	    RECT 75.0000 7.2000 75.3000 7.8000 ;
	    RECT 75.0000 6.8000 75.4000 7.2000 ;
	    RECT 71.8000 6.1000 72.1000 6.8000 ;
	    RECT 71.7000 5.7000 72.1000 6.1000 ;
	    RECT 74.3000 5.1000 74.6000 6.8000 ;
	    RECT 76.6000 6.2000 76.9000 12.8000 ;
	    RECT 78.2000 8.2000 78.5000 13.8000 ;
	    RECT 80.6000 12.8000 81.0000 13.2000 ;
	    RECT 77.4000 7.8000 77.8000 8.2000 ;
	    RECT 78.2000 7.8000 78.6000 8.2000 ;
	    RECT 79.8000 7.8000 80.2000 8.2000 ;
	    RECT 77.4000 7.2000 77.7000 7.8000 ;
	    RECT 79.8000 7.2000 80.1000 7.8000 ;
	    RECT 77.4000 6.8000 77.8000 7.2000 ;
	    RECT 78.2000 6.8000 78.6000 7.2000 ;
	    RECT 79.8000 6.8000 80.2000 7.2000 ;
	    RECT 78.2000 6.2000 78.5000 6.8000 ;
	    RECT 80.6000 6.2000 80.9000 12.8000 ;
	    RECT 82.2000 9.2000 82.5000 15.8000 ;
	    RECT 87.0000 15.2000 87.3000 15.8000 ;
	    RECT 84.6000 14.8000 85.0000 15.2000 ;
	    RECT 87.0000 14.8000 87.4000 15.2000 ;
	    RECT 91.8000 15.1000 92.2000 15.2000 ;
	    RECT 92.6000 15.1000 93.0000 15.2000 ;
	    RECT 91.8000 14.8000 93.0000 15.1000 ;
	    RECT 93.4000 15.1000 93.8000 15.2000 ;
	    RECT 94.2000 15.1000 94.6000 15.2000 ;
	    RECT 93.4000 14.8000 94.6000 15.1000 ;
	    RECT 95.0000 14.8000 95.4000 15.2000 ;
	    RECT 84.6000 14.2000 84.9000 14.8000 ;
	    RECT 84.6000 13.8000 85.0000 14.2000 ;
	    RECT 84.6000 12.8000 85.0000 13.2000 ;
	    RECT 86.2000 12.8000 86.6000 13.2000 ;
	    RECT 82.2000 8.8000 82.6000 9.2000 ;
	    RECT 83.8000 7.8000 84.2000 8.2000 ;
	    RECT 82.2000 6.8000 82.6000 7.2000 ;
	    RECT 83.0000 6.8000 83.4000 7.2000 ;
	    RECT 82.2000 6.2000 82.5000 6.8000 ;
	    RECT 76.6000 5.8000 77.0000 6.2000 ;
	    RECT 78.2000 5.8000 78.6000 6.2000 ;
	    RECT 80.6000 5.8000 81.0000 6.2000 ;
	    RECT 81.4000 6.1000 81.8000 6.2000 ;
	    RECT 82.2000 6.1000 82.6000 6.2000 ;
	    RECT 81.4000 5.8000 82.6000 6.1000 ;
	    RECT 71.1000 4.7000 71.5000 5.1000 ;
	    RECT 74.2000 4.7000 74.6000 5.1000 ;
	    RECT 83.0000 5.2000 83.3000 6.8000 ;
	    RECT 83.8000 6.2000 84.1000 7.8000 ;
	    RECT 84.6000 7.2000 84.9000 12.8000 ;
	    RECT 86.2000 10.2000 86.5000 12.8000 ;
	    RECT 87.0000 11.2000 87.3000 14.8000 ;
	    RECT 95.0000 14.2000 95.3000 14.8000 ;
	    RECT 87.8000 14.1000 88.2000 14.2000 ;
	    RECT 88.6000 14.1000 89.0000 14.2000 ;
	    RECT 87.8000 13.8000 89.0000 14.1000 ;
	    RECT 95.0000 13.8000 95.4000 14.2000 ;
	    RECT 89.4000 13.1000 89.8000 13.2000 ;
	    RECT 90.2000 13.1000 90.6000 13.2000 ;
	    RECT 89.4000 12.8000 90.6000 13.1000 ;
	    RECT 92.6000 12.8000 93.0000 13.2000 ;
	    RECT 94.2000 13.1000 94.6000 13.2000 ;
	    RECT 95.0000 13.1000 95.4000 13.2000 ;
	    RECT 94.2000 12.8000 95.4000 13.1000 ;
	    RECT 88.6000 11.8000 89.0000 12.2000 ;
	    RECT 87.0000 10.8000 87.4000 11.2000 ;
	    RECT 86.2000 9.8000 86.6000 10.2000 ;
	    RECT 88.6000 8.2000 88.9000 11.8000 ;
	    RECT 89.4000 9.8000 89.8000 10.2000 ;
	    RECT 89.4000 9.2000 89.7000 9.8000 ;
	    RECT 92.6000 9.2000 92.9000 12.8000 ;
	    RECT 89.4000 8.8000 89.8000 9.2000 ;
	    RECT 91.0000 8.8000 91.4000 9.2000 ;
	    RECT 92.6000 8.8000 93.0000 9.2000 ;
	    RECT 94.2000 8.8000 94.6000 9.2000 ;
	    RECT 88.6000 7.8000 89.0000 8.2000 ;
	    RECT 91.0000 7.2000 91.3000 8.8000 ;
	    RECT 91.8000 7.8000 92.2000 8.2000 ;
	    RECT 91.8000 7.2000 92.1000 7.8000 ;
	    RECT 94.2000 7.2000 94.5000 8.8000 ;
	    RECT 84.6000 6.8000 85.0000 7.2000 ;
	    RECT 85.4000 7.1000 85.8000 7.2000 ;
	    RECT 86.2000 7.1000 86.6000 7.2000 ;
	    RECT 85.4000 6.8000 86.6000 7.1000 ;
	    RECT 91.0000 6.8000 91.4000 7.2000 ;
	    RECT 91.8000 6.8000 92.2000 7.2000 ;
	    RECT 93.4000 6.8000 93.8000 7.2000 ;
	    RECT 94.2000 6.8000 94.6000 7.2000 ;
	    RECT 83.8000 5.8000 84.2000 6.2000 ;
	    RECT 86.2000 5.8000 86.6000 6.2000 ;
	    RECT 87.0000 5.8000 87.4000 6.2000 ;
	    RECT 89.4000 5.8000 89.8000 6.2000 ;
	    RECT 86.2000 5.2000 86.5000 5.8000 ;
	    RECT 87.0000 5.2000 87.3000 5.8000 ;
	    RECT 89.4000 5.2000 89.7000 5.8000 ;
	    RECT 93.4000 5.2000 93.7000 6.8000 ;
	    RECT 94.2000 6.1000 94.6000 6.2000 ;
	    RECT 95.0000 6.1000 95.4000 6.2000 ;
	    RECT 94.2000 5.8000 95.4000 6.1000 ;
	    RECT 95.8000 5.2000 96.1000 15.8000 ;
	    RECT 98.2000 13.8000 98.6000 14.2000 ;
	    RECT 99.8000 13.8000 100.2000 14.2000 ;
	    RECT 102.2000 14.1000 102.6000 14.2000 ;
	    RECT 103.0000 14.1000 103.4000 14.2000 ;
	    RECT 102.2000 13.8000 103.4000 14.1000 ;
	    RECT 98.2000 13.2000 98.5000 13.8000 ;
	    RECT 99.8000 13.2000 100.1000 13.8000 ;
	    RECT 98.2000 12.8000 98.6000 13.2000 ;
	    RECT 99.8000 12.8000 100.2000 13.2000 ;
	    RECT 100.6000 13.1000 101.0000 13.2000 ;
	    RECT 101.4000 13.1000 101.8000 13.2000 ;
	    RECT 100.6000 12.8000 101.8000 13.1000 ;
	    RECT 98.2000 10.8000 98.6000 11.2000 ;
	    RECT 98.2000 9.2000 98.5000 10.8000 ;
	    RECT 98.2000 8.8000 98.6000 9.2000 ;
	    RECT 103.8000 8.2000 104.1000 26.8000 ;
	    RECT 105.4000 26.2000 105.7000 26.8000 ;
	    RECT 105.4000 25.8000 105.8000 26.2000 ;
	    RECT 106.2000 25.2000 106.5000 31.8000 ;
	    RECT 117.4000 29.2000 117.7000 34.8000 ;
	    RECT 120.6000 34.2000 120.9000 35.8000 ;
	    RECT 121.4000 35.1000 121.8000 35.2000 ;
	    RECT 122.2000 35.1000 122.6000 35.2000 ;
	    RECT 121.4000 34.8000 122.6000 35.1000 ;
	    RECT 123.0000 35.1000 123.4000 35.2000 ;
	    RECT 123.0000 34.8000 124.1000 35.1000 ;
	    RECT 119.0000 34.1000 119.4000 34.2000 ;
	    RECT 119.8000 34.1000 120.2000 34.2000 ;
	    RECT 119.0000 33.8000 120.2000 34.1000 ;
	    RECT 120.6000 33.8000 121.0000 34.2000 ;
	    RECT 121.4000 34.1000 121.8000 34.2000 ;
	    RECT 122.2000 34.1000 122.6000 34.2000 ;
	    RECT 121.4000 33.8000 122.6000 34.1000 ;
	    RECT 122.2000 33.2000 122.5000 33.8000 ;
	    RECT 122.2000 32.8000 122.6000 33.2000 ;
	    RECT 123.8000 29.2000 124.1000 34.8000 ;
	    RECT 124.6000 34.8000 125.0000 35.2000 ;
	    RECT 124.6000 34.2000 124.9000 34.8000 ;
	    RECT 124.6000 33.8000 125.0000 34.2000 ;
	    RECT 108.6000 28.8000 109.0000 29.2000 ;
	    RECT 108.6000 28.2000 108.9000 28.8000 ;
	    RECT 107.8000 27.8000 108.2000 28.2000 ;
	    RECT 108.6000 27.8000 109.0000 28.2000 ;
	    RECT 111.0000 28.1000 111.4000 28.2000 ;
	    RECT 111.8000 28.1000 112.2000 28.2000 ;
	    RECT 111.0000 27.8000 112.2000 28.1000 ;
	    RECT 107.8000 26.2000 108.1000 27.8000 ;
	    RECT 110.2000 27.1000 110.6000 27.2000 ;
	    RECT 111.0000 27.1000 111.4000 27.2000 ;
	    RECT 110.2000 26.8000 111.4000 27.1000 ;
	    RECT 107.0000 25.8000 107.4000 26.2000 ;
	    RECT 107.8000 25.8000 108.2000 26.2000 ;
	    RECT 107.0000 25.2000 107.3000 25.8000 ;
	    RECT 106.2000 24.8000 106.6000 25.2000 ;
	    RECT 107.0000 24.8000 107.4000 25.2000 ;
	    RECT 111.8000 24.8000 112.2000 25.2000 ;
	    RECT 112.6000 25.1000 113.0000 27.9000 ;
	    RECT 111.8000 24.2000 112.1000 24.8000 ;
	    RECT 111.8000 23.8000 112.2000 24.2000 ;
	    RECT 114.2000 23.1000 114.6000 28.9000 ;
	    RECT 117.4000 28.8000 117.8000 29.2000 ;
	    RECT 121.4000 29.1000 121.8000 29.2000 ;
	    RECT 122.2000 29.1000 122.6000 29.2000 ;
	    RECT 115.0000 25.9000 115.4000 26.3000 ;
	    RECT 115.0000 25.2000 115.3000 25.9000 ;
	    RECT 118.2000 25.8000 118.6000 26.2000 ;
	    RECT 118.2000 25.2000 118.5000 25.8000 ;
	    RECT 115.0000 24.8000 115.4000 25.2000 ;
	    RECT 118.2000 24.8000 118.6000 25.2000 ;
	    RECT 119.0000 23.1000 119.4000 28.9000 ;
	    RECT 121.4000 28.8000 122.6000 29.1000 ;
	    RECT 123.8000 28.8000 124.2000 29.2000 ;
	    RECT 122.2000 28.1000 122.6000 28.2000 ;
	    RECT 123.0000 28.1000 123.4000 28.2000 ;
	    RECT 122.2000 27.8000 123.4000 28.1000 ;
	    RECT 119.0000 21.8000 119.4000 22.2000 ;
	    RECT 109.4000 16.1000 109.8000 16.2000 ;
	    RECT 110.2000 16.1000 110.6000 16.2000 ;
	    RECT 109.4000 15.8000 110.6000 16.1000 ;
	    RECT 118.2000 15.8000 118.6000 16.2000 ;
	    RECT 118.2000 15.2000 118.5000 15.8000 ;
	    RECT 111.8000 14.8000 112.2000 15.2000 ;
	    RECT 115.8000 15.1000 116.2000 15.2000 ;
	    RECT 116.6000 15.1000 117.0000 15.2000 ;
	    RECT 115.8000 14.8000 117.0000 15.1000 ;
	    RECT 118.2000 14.8000 118.6000 15.2000 ;
	    RECT 111.8000 14.2000 112.1000 14.8000 ;
	    RECT 105.4000 13.8000 105.8000 14.2000 ;
	    RECT 111.0000 13.8000 111.4000 14.2000 ;
	    RECT 111.8000 13.8000 112.2000 14.2000 ;
	    RECT 115.8000 13.8000 116.2000 14.2000 ;
	    RECT 105.4000 13.2000 105.7000 13.8000 ;
	    RECT 104.6000 12.8000 105.0000 13.2000 ;
	    RECT 105.4000 12.8000 105.8000 13.2000 ;
	    RECT 104.6000 11.2000 104.9000 12.8000 ;
	    RECT 111.0000 12.2000 111.3000 13.8000 ;
	    RECT 115.8000 13.2000 116.1000 13.8000 ;
	    RECT 119.0000 13.2000 119.3000 21.8000 ;
	    RECT 122.2000 15.8000 122.6000 16.2000 ;
	    RECT 122.2000 15.2000 122.5000 15.8000 ;
	    RECT 122.2000 14.8000 122.6000 15.2000 ;
	    RECT 122.2000 14.1000 122.6000 14.2000 ;
	    RECT 123.0000 14.1000 123.4000 14.2000 ;
	    RECT 122.2000 13.8000 123.4000 14.1000 ;
	    RECT 124.6000 13.2000 124.9000 33.8000 ;
	    RECT 127.0000 33.1000 127.4000 35.9000 ;
	    RECT 125.4000 30.8000 125.8000 31.2000 ;
	    RECT 125.4000 27.2000 125.7000 30.8000 ;
	    RECT 126.2000 28.8000 126.6000 29.2000 ;
	    RECT 126.2000 28.2000 126.5000 28.8000 ;
	    RECT 127.8000 28.2000 128.1000 44.8000 ;
	    RECT 135.0000 44.2000 135.3000 44.8000 ;
	    RECT 135.0000 43.8000 135.4000 44.2000 ;
	    RECT 143.0000 43.1000 143.4000 48.9000 ;
	    RECT 143.8000 48.2000 144.1000 54.8000 ;
	    RECT 147.0000 48.2000 147.3000 55.8000 ;
	    RECT 148.6000 55.2000 148.9000 55.8000 ;
	    RECT 148.6000 54.8000 149.0000 55.2000 ;
	    RECT 153.4000 54.8000 153.8000 55.2000 ;
	    RECT 143.8000 47.8000 144.2000 48.2000 ;
	    RECT 147.0000 47.8000 147.4000 48.2000 ;
	    RECT 143.8000 45.9000 144.2000 46.3000 ;
	    RECT 143.8000 45.2000 144.1000 45.9000 ;
	    RECT 143.8000 44.8000 144.2000 45.2000 ;
	    RECT 147.8000 43.1000 148.2000 48.9000 ;
	    RECT 151.0000 45.1000 151.4000 47.9000 ;
	    RECT 152.6000 43.1000 153.0000 48.9000 ;
	    RECT 153.4000 44.2000 153.7000 54.8000 ;
	    RECT 154.2000 54.2000 154.5000 55.8000 ;
	    RECT 157.4000 54.8000 157.8000 55.2000 ;
	    RECT 154.2000 53.8000 154.6000 54.2000 ;
	    RECT 155.8000 53.1000 156.2000 53.2000 ;
	    RECT 156.6000 53.1000 157.0000 53.2000 ;
	    RECT 155.8000 52.8000 157.0000 53.1000 ;
	    RECT 155.0000 51.8000 155.4000 52.2000 ;
	    RECT 155.0000 46.2000 155.3000 51.8000 ;
	    RECT 157.4000 50.2000 157.7000 54.8000 ;
	    RECT 158.2000 53.8000 158.6000 54.2000 ;
	    RECT 158.2000 53.2000 158.5000 53.8000 ;
	    RECT 158.2000 52.8000 158.6000 53.2000 ;
	    RECT 161.4000 53.1000 161.8000 55.9000 ;
	    RECT 162.2000 55.2000 162.5000 61.8000 ;
	    RECT 163.0000 60.2000 163.3000 71.8000 ;
	    RECT 163.8000 61.8000 164.2000 62.2000 ;
	    RECT 163.0000 59.8000 163.4000 60.2000 ;
	    RECT 162.2000 54.8000 162.6000 55.2000 ;
	    RECT 162.2000 54.2000 162.5000 54.8000 ;
	    RECT 162.2000 53.8000 162.6000 54.2000 ;
	    RECT 163.0000 52.1000 163.4000 57.9000 ;
	    RECT 163.8000 55.1000 164.1000 61.8000 ;
	    RECT 163.8000 54.7000 164.2000 55.1000 ;
	    RECT 157.4000 49.8000 157.8000 50.2000 ;
	    RECT 159.8000 49.8000 160.2000 50.2000 ;
	    RECT 159.8000 49.2000 160.1000 49.8000 ;
	    RECT 155.0000 45.8000 155.4000 46.2000 ;
	    RECT 155.8000 45.8000 156.2000 46.2000 ;
	    RECT 153.4000 43.8000 153.8000 44.2000 ;
	    RECT 128.6000 32.1000 129.0000 37.9000 ;
	    RECT 129.4000 34.7000 129.8000 35.1000 ;
	    RECT 132.6000 34.8000 133.0000 35.2000 ;
	    RECT 129.4000 34.2000 129.7000 34.7000 ;
	    RECT 129.4000 33.8000 129.8000 34.2000 ;
	    RECT 131.8000 30.8000 132.2000 31.2000 ;
	    RECT 130.2000 29.8000 130.6000 30.2000 ;
	    RECT 128.6000 29.1000 129.0000 29.2000 ;
	    RECT 129.4000 29.1000 129.8000 29.2000 ;
	    RECT 128.6000 28.8000 129.8000 29.1000 ;
	    RECT 126.2000 27.8000 126.6000 28.2000 ;
	    RECT 127.8000 27.8000 128.2000 28.2000 ;
	    RECT 125.4000 26.8000 125.8000 27.2000 ;
	    RECT 125.4000 26.1000 125.8000 26.2000 ;
	    RECT 126.2000 26.1000 126.6000 26.2000 ;
	    RECT 125.4000 25.8000 126.6000 26.1000 ;
	    RECT 127.8000 26.1000 128.2000 26.2000 ;
	    RECT 128.6000 26.1000 129.0000 26.2000 ;
	    RECT 127.8000 25.8000 129.0000 26.1000 ;
	    RECT 130.2000 25.2000 130.5000 29.8000 ;
	    RECT 131.0000 28.8000 131.4000 29.2000 ;
	    RECT 131.0000 28.2000 131.3000 28.8000 ;
	    RECT 131.8000 28.2000 132.1000 30.8000 ;
	    RECT 132.6000 30.2000 132.9000 34.8000 ;
	    RECT 133.4000 32.1000 133.8000 37.9000 ;
	    RECT 139.0000 36.8000 139.4000 37.2000 ;
	    RECT 139.0000 36.2000 139.3000 36.8000 ;
	    RECT 139.0000 35.8000 139.4000 36.2000 ;
	    RECT 139.8000 35.8000 140.2000 36.2000 ;
	    RECT 139.8000 35.2000 140.1000 35.8000 ;
	    RECT 137.4000 35.1000 137.8000 35.2000 ;
	    RECT 138.2000 35.1000 138.6000 35.2000 ;
	    RECT 137.4000 34.8000 138.6000 35.1000 ;
	    RECT 139.8000 34.8000 140.2000 35.2000 ;
	    RECT 134.2000 33.8000 134.6000 34.2000 ;
	    RECT 136.6000 33.8000 137.0000 34.2000 ;
	    RECT 140.6000 34.1000 141.0000 34.2000 ;
	    RECT 141.4000 34.1000 141.8000 34.2000 ;
	    RECT 140.6000 33.8000 141.8000 34.1000 ;
	    RECT 132.6000 29.8000 133.0000 30.2000 ;
	    RECT 132.6000 29.1000 133.0000 29.2000 ;
	    RECT 133.4000 29.1000 133.8000 29.2000 ;
	    RECT 132.6000 28.8000 133.8000 29.1000 ;
	    RECT 131.0000 27.8000 131.4000 28.2000 ;
	    RECT 131.8000 27.8000 132.2000 28.2000 ;
	    RECT 131.0000 27.1000 131.4000 27.2000 ;
	    RECT 131.8000 27.1000 132.2000 27.2000 ;
	    RECT 131.0000 26.8000 132.2000 27.1000 ;
	    RECT 134.2000 26.2000 134.5000 33.8000 ;
	    RECT 136.6000 33.2000 136.9000 33.8000 ;
	    RECT 136.6000 32.8000 137.0000 33.2000 ;
	    RECT 139.0000 32.8000 139.4000 33.2000 ;
	    RECT 141.4000 33.1000 141.8000 33.2000 ;
	    RECT 142.2000 33.1000 142.6000 33.2000 ;
	    RECT 143.0000 33.1000 143.4000 35.9000 ;
	    RECT 141.4000 32.8000 142.6000 33.1000 ;
	    RECT 135.8000 31.8000 136.2000 32.2000 ;
	    RECT 135.8000 31.2000 136.1000 31.8000 ;
	    RECT 135.8000 30.8000 136.2000 31.2000 ;
	    RECT 139.0000 28.2000 139.3000 32.8000 ;
	    RECT 144.6000 32.1000 145.0000 37.9000 ;
	    RECT 145.4000 36.8000 145.8000 37.2000 ;
	    RECT 145.4000 35.1000 145.7000 36.8000 ;
	    RECT 145.4000 34.7000 145.8000 35.1000 ;
	    RECT 145.4000 32.8000 145.8000 33.2000 ;
	    RECT 145.4000 30.2000 145.7000 32.8000 ;
	    RECT 149.4000 32.1000 149.8000 37.9000 ;
	    RECT 154.2000 35.8000 154.6000 36.2000 ;
	    RECT 154.2000 34.2000 154.5000 35.8000 ;
	    RECT 155.8000 35.2000 156.1000 45.8000 ;
	    RECT 157.4000 43.1000 157.8000 48.9000 ;
	    RECT 159.8000 48.8000 160.2000 49.2000 ;
	    RECT 158.2000 44.8000 158.6000 45.2000 ;
	    RECT 156.6000 36.1000 157.0000 36.2000 ;
	    RECT 157.4000 36.1000 157.8000 36.2000 ;
	    RECT 156.6000 35.8000 157.8000 36.1000 ;
	    RECT 155.8000 34.8000 156.2000 35.2000 ;
	    RECT 151.8000 33.8000 152.2000 34.2000 ;
	    RECT 152.6000 33.8000 153.0000 34.2000 ;
	    RECT 154.2000 33.8000 154.6000 34.2000 ;
	    RECT 151.8000 32.2000 152.1000 33.8000 ;
	    RECT 151.8000 31.8000 152.2000 32.2000 ;
	    RECT 152.6000 31.2000 152.9000 33.8000 ;
	    RECT 158.2000 33.2000 158.5000 44.8000 ;
	    RECT 163.0000 42.1000 163.4000 42.2000 ;
	    RECT 163.8000 42.1000 164.2000 42.2000 ;
	    RECT 163.0000 41.8000 164.2000 42.1000 ;
	    RECT 159.0000 34.8000 159.4000 35.2000 ;
	    RECT 158.2000 32.8000 158.6000 33.2000 ;
	    RECT 155.8000 32.1000 156.2000 32.2000 ;
	    RECT 156.6000 32.1000 157.0000 32.2000 ;
	    RECT 155.8000 31.8000 157.0000 32.1000 ;
	    RECT 157.4000 31.8000 157.8000 32.2000 ;
	    RECT 152.6000 30.8000 153.0000 31.2000 ;
	    RECT 145.4000 29.8000 145.8000 30.2000 ;
	    RECT 141.4000 28.8000 141.8000 29.2000 ;
	    RECT 139.0000 27.8000 139.4000 28.2000 ;
	    RECT 140.6000 27.8000 141.0000 28.2000 ;
	    RECT 139.0000 27.2000 139.3000 27.8000 ;
	    RECT 140.6000 27.2000 140.9000 27.8000 ;
	    RECT 135.0000 27.1000 135.4000 27.2000 ;
	    RECT 135.8000 27.1000 136.2000 27.2000 ;
	    RECT 135.0000 26.8000 136.2000 27.1000 ;
	    RECT 139.0000 26.8000 139.4000 27.2000 ;
	    RECT 140.6000 27.1000 141.0000 27.2000 ;
	    RECT 141.4000 27.1000 141.7000 28.8000 ;
	    RECT 140.6000 26.8000 141.7000 27.1000 ;
	    RECT 134.2000 25.8000 134.6000 26.2000 ;
	    RECT 135.8000 26.1000 136.2000 26.2000 ;
	    RECT 136.6000 26.1000 137.0000 26.2000 ;
	    RECT 135.8000 25.8000 137.0000 26.1000 ;
	    RECT 130.2000 24.8000 130.6000 25.2000 ;
	    RECT 135.8000 25.1000 136.2000 25.2000 ;
	    RECT 136.6000 25.1000 137.0000 25.2000 ;
	    RECT 135.8000 24.8000 137.0000 25.1000 ;
	    RECT 138.2000 24.8000 138.6000 25.2000 ;
	    RECT 112.6000 13.1000 113.0000 13.2000 ;
	    RECT 113.4000 13.1000 113.8000 13.2000 ;
	    RECT 112.6000 12.8000 113.8000 13.1000 ;
	    RECT 115.8000 12.8000 116.2000 13.2000 ;
	    RECT 116.6000 12.8000 117.0000 13.2000 ;
	    RECT 119.0000 12.8000 119.4000 13.2000 ;
	    RECT 123.0000 12.8000 123.4000 13.2000 ;
	    RECT 123.8000 13.1000 124.2000 13.2000 ;
	    RECT 124.6000 13.1000 125.0000 13.2000 ;
	    RECT 123.8000 12.8000 125.0000 13.1000 ;
	    RECT 111.0000 11.8000 111.4000 12.2000 ;
	    RECT 104.6000 10.8000 105.0000 11.2000 ;
	    RECT 116.6000 10.2000 116.9000 12.8000 ;
	    RECT 117.4000 11.8000 117.8000 12.2000 ;
	    RECT 120.6000 12.1000 121.0000 12.2000 ;
	    RECT 121.4000 12.1000 121.8000 12.2000 ;
	    RECT 120.6000 11.8000 121.8000 12.1000 ;
	    RECT 110.2000 9.8000 110.6000 10.2000 ;
	    RECT 112.6000 9.8000 113.0000 10.2000 ;
	    RECT 116.6000 9.8000 117.0000 10.2000 ;
	    RECT 105.4000 8.8000 105.8000 9.2000 ;
	    RECT 105.4000 8.2000 105.7000 8.8000 ;
	    RECT 110.2000 8.2000 110.5000 9.8000 ;
	    RECT 111.0000 8.8000 111.4000 9.2000 ;
	    RECT 97.4000 8.1000 97.8000 8.2000 ;
	    RECT 98.2000 8.1000 98.6000 8.2000 ;
	    RECT 97.4000 7.8000 98.6000 8.1000 ;
	    RECT 100.6000 7.8000 101.0000 8.2000 ;
	    RECT 102.2000 8.1000 102.6000 8.2000 ;
	    RECT 103.0000 8.1000 103.4000 8.2000 ;
	    RECT 102.2000 7.8000 103.4000 8.1000 ;
	    RECT 103.8000 7.8000 104.2000 8.2000 ;
	    RECT 105.4000 7.8000 105.8000 8.2000 ;
	    RECT 110.2000 7.8000 110.6000 8.2000 ;
	    RECT 100.6000 7.2000 100.9000 7.8000 ;
	    RECT 96.6000 6.8000 97.0000 7.2000 ;
	    RECT 98.2000 7.1000 98.6000 7.2000 ;
	    RECT 99.0000 7.1000 99.4000 7.2000 ;
	    RECT 98.2000 6.8000 99.4000 7.1000 ;
	    RECT 99.8000 6.8000 100.2000 7.2000 ;
	    RECT 100.6000 6.8000 101.0000 7.2000 ;
	    RECT 102.2000 7.1000 102.6000 7.2000 ;
	    RECT 103.0000 7.1000 103.4000 7.2000 ;
	    RECT 102.2000 6.8000 103.4000 7.1000 ;
	    RECT 103.8000 7.1000 104.1000 7.8000 ;
	    RECT 111.0000 7.2000 111.3000 8.8000 ;
	    RECT 111.8000 7.5000 112.2000 7.9000 ;
	    RECT 112.6000 7.8000 112.9000 9.8000 ;
	    RECT 117.4000 9.2000 117.7000 11.8000 ;
	    RECT 123.0000 9.2000 123.3000 12.8000 ;
	    RECT 124.6000 12.1000 125.0000 12.2000 ;
	    RECT 127.0000 12.1000 127.4000 17.9000 ;
	    RECT 130.2000 14.2000 130.5000 24.8000 ;
	    RECT 138.2000 24.2000 138.5000 24.8000 ;
	    RECT 138.2000 23.8000 138.6000 24.2000 ;
	    RECT 143.8000 23.1000 144.2000 28.9000 ;
	    RECT 145.4000 27.2000 145.7000 29.8000 ;
	    RECT 145.4000 26.8000 145.8000 27.2000 ;
	    RECT 147.0000 25.8000 147.4000 26.2000 ;
	    RECT 147.0000 25.2000 147.3000 25.8000 ;
	    RECT 147.0000 24.8000 147.4000 25.2000 ;
	    RECT 148.6000 23.1000 149.0000 28.9000 ;
	    RECT 153.4000 28.8000 153.8000 29.2000 ;
	    RECT 153.4000 28.2000 153.7000 28.8000 ;
	    RECT 149.4000 27.8000 149.8000 28.2000 ;
	    RECT 149.4000 27.2000 149.7000 27.8000 ;
	    RECT 149.4000 26.8000 149.8000 27.2000 ;
	    RECT 150.2000 25.1000 150.6000 27.9000 ;
	    RECT 151.0000 27.8000 151.4000 28.2000 ;
	    RECT 153.4000 27.8000 153.8000 28.2000 ;
	    RECT 151.0000 26.2000 151.3000 27.8000 ;
	    RECT 151.8000 26.8000 152.2000 27.2000 ;
	    RECT 152.6000 27.1000 153.0000 27.2000 ;
	    RECT 153.4000 27.1000 153.8000 27.2000 ;
	    RECT 152.6000 26.8000 153.8000 27.1000 ;
	    RECT 151.8000 26.2000 152.1000 26.8000 ;
	    RECT 151.0000 25.8000 151.4000 26.2000 ;
	    RECT 151.8000 25.8000 152.2000 26.2000 ;
	    RECT 153.4000 25.8000 153.8000 26.2000 ;
	    RECT 153.4000 25.2000 153.7000 25.8000 ;
	    RECT 153.4000 24.8000 153.8000 25.2000 ;
	    RECT 154.2000 25.1000 154.6000 27.9000 ;
	    RECT 155.8000 23.1000 156.2000 28.9000 ;
	    RECT 157.4000 28.2000 157.7000 31.8000 ;
	    RECT 157.4000 27.8000 157.8000 28.2000 ;
	    RECT 156.6000 25.9000 157.0000 26.3000 ;
	    RECT 159.0000 26.2000 159.3000 34.8000 ;
	    RECT 160.6000 32.1000 161.0000 32.2000 ;
	    RECT 161.4000 32.1000 161.8000 32.2000 ;
	    RECT 163.0000 32.1000 163.4000 37.9000 ;
	    RECT 164.6000 37.2000 164.9000 71.8000 ;
	    RECT 165.4000 68.1000 165.8000 68.2000 ;
	    RECT 166.2000 68.1000 166.6000 68.2000 ;
	    RECT 165.4000 67.8000 166.6000 68.1000 ;
	    RECT 165.4000 58.8000 165.8000 59.2000 ;
	    RECT 165.4000 48.2000 165.7000 58.8000 ;
	    RECT 166.2000 54.2000 166.5000 67.8000 ;
	    RECT 167.0000 55.2000 167.3000 72.8000 ;
	    RECT 169.4000 72.1000 169.8000 77.9000 ;
	    RECT 173.4000 75.2000 173.7000 86.8000 ;
	    RECT 174.2000 83.1000 174.6000 88.9000 ;
	    RECT 175.0000 88.2000 175.3000 93.8000 ;
	    RECT 175.8000 92.1000 176.2000 97.9000 ;
	    RECT 177.4000 97.8000 177.8000 98.2000 ;
	    RECT 177.4000 94.8000 177.8000 95.2000 ;
	    RECT 177.4000 94.2000 177.7000 94.8000 ;
	    RECT 177.4000 93.8000 177.8000 94.2000 ;
	    RECT 180.6000 92.1000 181.0000 97.9000 ;
	    RECT 181.4000 93.2000 181.7000 103.8000 ;
	    RECT 183.0000 96.8000 183.4000 97.2000 ;
	    RECT 183.0000 95.2000 183.3000 96.8000 ;
	    RECT 183.0000 94.8000 183.4000 95.2000 ;
	    RECT 183.8000 94.2000 184.1000 109.8000 ;
	    RECT 184.6000 109.2000 184.9000 152.8000 ;
	    RECT 185.4000 148.8000 185.8000 149.2000 ;
	    RECT 186.2000 148.8000 186.6000 149.2000 ;
	    RECT 185.4000 148.2000 185.7000 148.8000 ;
	    RECT 186.2000 148.2000 186.5000 148.8000 ;
	    RECT 185.4000 147.8000 185.8000 148.2000 ;
	    RECT 186.2000 147.8000 186.6000 148.2000 ;
	    RECT 185.4000 147.1000 185.8000 147.2000 ;
	    RECT 186.2000 147.1000 186.6000 147.2000 ;
	    RECT 185.4000 146.8000 186.6000 147.1000 ;
	    RECT 186.2000 141.8000 186.6000 142.2000 ;
	    RECT 185.4000 134.8000 185.8000 135.2000 ;
	    RECT 185.4000 126.2000 185.7000 134.8000 ;
	    RECT 186.2000 129.2000 186.5000 141.8000 ;
	    RECT 187.0000 140.2000 187.3000 153.8000 ;
	    RECT 189.4000 152.2000 189.7000 154.8000 ;
	    RECT 190.2000 153.8000 190.6000 154.2000 ;
	    RECT 189.4000 151.8000 189.8000 152.2000 ;
	    RECT 187.8000 149.8000 188.2000 150.2000 ;
	    RECT 187.8000 146.2000 188.1000 149.8000 ;
	    RECT 188.6000 146.8000 189.0000 147.2000 ;
	    RECT 188.6000 146.2000 188.9000 146.8000 ;
	    RECT 187.8000 145.8000 188.2000 146.2000 ;
	    RECT 188.6000 145.8000 189.0000 146.2000 ;
	    RECT 189.4000 145.8000 189.8000 146.2000 ;
	    RECT 189.4000 145.2000 189.7000 145.8000 ;
	    RECT 187.8000 144.8000 188.2000 145.2000 ;
	    RECT 189.4000 144.8000 189.8000 145.2000 ;
	    RECT 187.8000 144.2000 188.1000 144.8000 ;
	    RECT 187.8000 143.8000 188.2000 144.2000 ;
	    RECT 187.0000 139.8000 187.4000 140.2000 ;
	    RECT 190.2000 135.2000 190.5000 153.8000 ;
	    RECT 192.6000 153.2000 192.9000 154.8000 ;
	    RECT 193.4000 154.2000 193.7000 154.8000 ;
	    RECT 193.4000 153.8000 193.8000 154.2000 ;
	    RECT 197.4000 154.1000 197.8000 154.2000 ;
	    RECT 198.2000 154.1000 198.6000 154.2000 ;
	    RECT 197.4000 153.8000 198.6000 154.1000 ;
	    RECT 199.0000 154.1000 199.4000 154.2000 ;
	    RECT 199.8000 154.1000 200.2000 154.2000 ;
	    RECT 199.0000 153.8000 200.2000 154.1000 ;
	    RECT 201.4000 153.8000 201.8000 154.2000 ;
	    RECT 192.6000 152.8000 193.0000 153.2000 ;
	    RECT 198.2000 153.1000 198.6000 153.2000 ;
	    RECT 199.0000 153.1000 199.4000 153.2000 ;
	    RECT 198.2000 152.8000 199.4000 153.1000 ;
	    RECT 191.8000 151.8000 192.2000 152.2000 ;
	    RECT 191.8000 148.2000 192.1000 151.8000 ;
	    RECT 193.4000 150.8000 193.8000 151.2000 ;
	    RECT 191.8000 147.8000 192.2000 148.2000 ;
	    RECT 191.0000 146.8000 191.4000 147.2000 ;
	    RECT 191.0000 146.2000 191.3000 146.8000 ;
	    RECT 191.8000 146.2000 192.1000 147.8000 ;
	    RECT 193.4000 147.2000 193.7000 150.8000 ;
	    RECT 197.4000 149.1000 197.8000 149.2000 ;
	    RECT 198.2000 149.1000 198.6000 149.2000 ;
	    RECT 197.4000 148.8000 198.6000 149.1000 ;
	    RECT 193.4000 146.8000 193.8000 147.2000 ;
	    RECT 193.4000 146.2000 193.7000 146.8000 ;
	    RECT 191.0000 145.8000 191.4000 146.2000 ;
	    RECT 191.8000 145.8000 192.2000 146.2000 ;
	    RECT 193.4000 145.8000 193.8000 146.2000 ;
	    RECT 194.2000 145.8000 194.6000 146.2000 ;
	    RECT 195.8000 146.1000 196.2000 146.2000 ;
	    RECT 196.6000 146.1000 197.0000 146.2000 ;
	    RECT 195.8000 145.8000 197.0000 146.1000 ;
	    RECT 191.0000 144.8000 191.4000 145.2000 ;
	    RECT 191.0000 144.2000 191.3000 144.8000 ;
	    RECT 191.0000 143.8000 191.4000 144.2000 ;
	    RECT 187.8000 135.1000 188.2000 135.2000 ;
	    RECT 188.6000 135.1000 189.0000 135.2000 ;
	    RECT 187.8000 134.8000 189.0000 135.1000 ;
	    RECT 190.2000 134.8000 190.6000 135.2000 ;
	    RECT 187.0000 131.8000 187.4000 132.2000 ;
	    RECT 190.2000 131.8000 190.6000 132.2000 ;
	    RECT 186.2000 128.8000 186.6000 129.2000 ;
	    RECT 185.4000 125.8000 185.8000 126.2000 ;
	    RECT 185.4000 125.1000 185.8000 125.2000 ;
	    RECT 186.2000 125.1000 186.6000 125.2000 ;
	    RECT 185.4000 124.8000 186.6000 125.1000 ;
	    RECT 185.4000 111.8000 185.8000 112.2000 ;
	    RECT 184.6000 108.8000 185.0000 109.2000 ;
	    RECT 185.4000 107.2000 185.7000 111.8000 ;
	    RECT 187.0000 111.2000 187.3000 131.8000 ;
	    RECT 188.6000 127.1000 189.0000 127.2000 ;
	    RECT 189.4000 127.1000 189.8000 127.2000 ;
	    RECT 188.6000 126.8000 189.8000 127.1000 ;
	    RECT 190.2000 125.1000 190.5000 131.8000 ;
	    RECT 191.8000 131.2000 192.1000 145.8000 ;
	    RECT 194.2000 145.2000 194.5000 145.8000 ;
	    RECT 194.2000 144.8000 194.6000 145.2000 ;
	    RECT 192.6000 143.1000 193.0000 143.2000 ;
	    RECT 193.4000 143.1000 193.8000 143.2000 ;
	    RECT 199.8000 143.1000 200.2000 148.9000 ;
	    RECT 192.6000 142.8000 193.8000 143.1000 ;
	    RECT 201.4000 141.2000 201.7000 153.8000 ;
	    RECT 202.2000 153.1000 202.6000 155.9000 ;
	    RECT 203.0000 154.2000 203.3000 163.8000 ;
	    RECT 203.0000 153.8000 203.4000 154.2000 ;
	    RECT 203.0000 147.2000 203.3000 153.8000 ;
	    RECT 203.8000 152.1000 204.2000 157.9000 ;
	    RECT 204.6000 154.7000 205.0000 155.1000 ;
	    RECT 204.6000 154.2000 204.9000 154.7000 ;
	    RECT 204.6000 153.8000 205.0000 154.2000 ;
	    RECT 205.4000 153.2000 205.7000 167.8000 ;
	    RECT 208.6000 167.1000 209.0000 167.2000 ;
	    RECT 209.4000 167.1000 209.7000 167.8000 ;
	    RECT 214.2000 167.2000 214.5000 169.8000 ;
	    RECT 217.4000 167.2000 217.7000 173.8000 ;
	    RECT 219.0000 172.8000 219.4000 173.2000 ;
	    RECT 219.0000 172.2000 219.3000 172.8000 ;
	    RECT 220.6000 172.2000 220.9000 174.8000 ;
	    RECT 222.2000 174.2000 222.5000 174.8000 ;
	    RECT 227.8000 174.2000 228.1000 174.8000 ;
	    RECT 222.2000 173.8000 222.6000 174.2000 ;
	    RECT 223.0000 174.1000 223.4000 174.2000 ;
	    RECT 223.8000 174.1000 224.2000 174.2000 ;
	    RECT 223.0000 173.8000 224.2000 174.1000 ;
	    RECT 224.6000 173.8000 225.0000 174.2000 ;
	    RECT 225.4000 174.1000 225.8000 174.2000 ;
	    RECT 226.2000 174.1000 226.6000 174.2000 ;
	    RECT 225.4000 173.8000 226.6000 174.1000 ;
	    RECT 227.8000 173.8000 228.2000 174.2000 ;
	    RECT 224.6000 172.2000 224.9000 173.8000 ;
	    RECT 227.0000 173.1000 227.4000 173.2000 ;
	    RECT 227.8000 173.1000 228.2000 173.2000 ;
	    RECT 228.6000 173.1000 229.0000 175.9000 ;
	    RECT 229.4000 173.8000 229.8000 174.2000 ;
	    RECT 227.0000 172.8000 228.2000 173.1000 ;
	    RECT 219.0000 171.8000 219.4000 172.2000 ;
	    RECT 220.6000 171.8000 221.0000 172.2000 ;
	    RECT 222.2000 171.8000 222.6000 172.2000 ;
	    RECT 224.6000 171.8000 225.0000 172.2000 ;
	    RECT 218.2000 168.8000 218.6000 169.2000 ;
	    RECT 218.2000 168.2000 218.5000 168.8000 ;
	    RECT 218.2000 167.8000 218.6000 168.2000 ;
	    RECT 208.6000 166.8000 209.7000 167.1000 ;
	    RECT 210.2000 166.8000 210.6000 167.2000 ;
	    RECT 214.2000 166.8000 214.6000 167.2000 ;
	    RECT 216.6000 167.1000 217.0000 167.2000 ;
	    RECT 217.4000 167.1000 217.8000 167.2000 ;
	    RECT 216.6000 166.8000 217.8000 167.1000 ;
	    RECT 210.2000 166.2000 210.5000 166.8000 ;
	    RECT 218.2000 166.2000 218.5000 167.8000 ;
	    RECT 207.8000 166.1000 208.2000 166.2000 ;
	    RECT 208.6000 166.1000 209.0000 166.2000 ;
	    RECT 207.8000 165.8000 209.0000 166.1000 ;
	    RECT 210.2000 165.8000 210.6000 166.2000 ;
	    RECT 214.2000 166.1000 214.6000 166.2000 ;
	    RECT 215.0000 166.1000 215.4000 166.2000 ;
	    RECT 214.2000 165.8000 215.4000 166.1000 ;
	    RECT 218.2000 165.8000 218.6000 166.2000 ;
	    RECT 210.2000 161.2000 210.5000 165.8000 ;
	    RECT 215.0000 165.1000 215.4000 165.2000 ;
	    RECT 215.8000 165.1000 216.2000 165.2000 ;
	    RECT 215.0000 164.8000 216.2000 165.1000 ;
	    RECT 219.0000 162.2000 219.3000 171.8000 ;
	    RECT 220.6000 169.8000 221.0000 170.2000 ;
	    RECT 220.6000 169.2000 220.9000 169.8000 ;
	    RECT 220.6000 168.8000 221.0000 169.2000 ;
	    RECT 222.2000 167.2000 222.5000 171.8000 ;
	    RECT 223.0000 168.8000 223.4000 169.2000 ;
	    RECT 227.0000 168.8000 227.4000 169.2000 ;
	    RECT 223.0000 167.2000 223.3000 168.8000 ;
	    RECT 227.0000 168.2000 227.3000 168.8000 ;
	    RECT 229.4000 168.2000 229.7000 173.8000 ;
	    RECT 230.2000 172.1000 230.6000 177.9000 ;
	    RECT 231.0000 175.0000 231.4000 175.1000 ;
	    RECT 231.8000 175.0000 232.2000 175.1000 ;
	    RECT 231.0000 174.7000 232.2000 175.0000 ;
	    RECT 235.0000 172.1000 235.4000 177.9000 ;
	    RECT 250.2000 177.8000 250.6000 178.2000 ;
	    RECT 238.2000 176.8000 238.6000 177.2000 ;
	    RECT 238.2000 176.2000 238.5000 176.8000 ;
	    RECT 238.2000 175.8000 238.6000 176.2000 ;
	    RECT 239.8000 175.8000 240.2000 176.2000 ;
	    RECT 238.2000 174.2000 238.5000 175.8000 ;
	    RECT 239.8000 175.2000 240.1000 175.8000 ;
	    RECT 239.8000 174.8000 240.2000 175.2000 ;
	    RECT 243.0000 174.8000 243.4000 175.2000 ;
	    RECT 247.0000 174.8000 247.4000 175.2000 ;
	    RECT 243.0000 174.2000 243.3000 174.8000 ;
	    RECT 247.0000 174.2000 247.3000 174.8000 ;
	    RECT 250.2000 174.4000 250.5000 177.8000 ;
	    RECT 254.2000 175.8000 254.6000 176.2000 ;
	    RECT 252.6000 174.8000 253.0000 175.2000 ;
	    RECT 238.2000 174.1000 238.6000 174.2000 ;
	    RECT 239.0000 174.1000 239.4000 174.2000 ;
	    RECT 238.2000 173.8000 239.4000 174.1000 ;
	    RECT 240.6000 173.8000 241.0000 174.2000 ;
	    RECT 242.2000 173.8000 242.6000 174.2000 ;
	    RECT 243.0000 173.8000 243.4000 174.2000 ;
	    RECT 247.0000 173.8000 247.4000 174.2000 ;
	    RECT 248.6000 174.1000 249.0000 174.2000 ;
	    RECT 249.4000 174.1000 249.8000 174.2000 ;
	    RECT 248.6000 173.8000 249.8000 174.1000 ;
	    RECT 250.2000 174.0000 250.6000 174.4000 ;
	    RECT 240.6000 173.2000 240.9000 173.8000 ;
	    RECT 242.2000 173.2000 242.5000 173.8000 ;
	    RECT 240.6000 172.8000 241.0000 173.2000 ;
	    RECT 242.2000 172.8000 242.6000 173.2000 ;
	    RECT 243.0000 172.8000 243.4000 173.2000 ;
	    RECT 245.4000 173.1000 245.8000 173.2000 ;
	    RECT 246.2000 173.1000 246.6000 173.2000 ;
	    RECT 245.4000 172.8000 246.6000 173.1000 ;
	    RECT 243.0000 172.2000 243.3000 172.8000 ;
	    RECT 239.0000 172.1000 239.4000 172.2000 ;
	    RECT 239.8000 172.1000 240.2000 172.2000 ;
	    RECT 239.0000 171.8000 240.2000 172.1000 ;
	    RECT 243.0000 171.8000 243.4000 172.2000 ;
	    RECT 245.4000 172.1000 245.8000 172.2000 ;
	    RECT 246.2000 172.1000 246.6000 172.2000 ;
	    RECT 245.4000 171.8000 246.6000 172.1000 ;
	    RECT 247.0000 169.2000 247.3000 173.8000 ;
	    RECT 250.2000 173.2000 250.5000 174.0000 ;
	    RECT 248.6000 173.1000 249.0000 173.2000 ;
	    RECT 249.4000 173.1000 249.8000 173.2000 ;
	    RECT 248.6000 172.8000 249.8000 173.1000 ;
	    RECT 250.2000 172.8000 250.6000 173.2000 ;
	    RECT 247.8000 171.8000 248.2000 172.2000 ;
	    RECT 251.8000 171.8000 252.2000 172.2000 ;
	    RECT 247.8000 169.2000 248.1000 171.8000 ;
	    RECT 235.0000 169.1000 235.4000 169.2000 ;
	    RECT 235.8000 169.1000 236.2000 169.2000 ;
	    RECT 235.0000 168.8000 236.2000 169.1000 ;
	    RECT 239.0000 168.8000 239.4000 169.2000 ;
	    RECT 239.8000 169.1000 240.2000 169.2000 ;
	    RECT 240.6000 169.1000 241.0000 169.2000 ;
	    RECT 239.8000 168.8000 241.0000 169.1000 ;
	    RECT 245.4000 168.8000 245.8000 169.2000 ;
	    RECT 247.0000 168.8000 247.4000 169.2000 ;
	    RECT 247.8000 168.8000 248.2000 169.2000 ;
	    RECT 227.0000 167.8000 227.4000 168.2000 ;
	    RECT 229.4000 167.8000 229.8000 168.2000 ;
	    RECT 239.0000 167.2000 239.3000 168.8000 ;
	    RECT 245.4000 167.2000 245.7000 168.8000 ;
	    RECT 222.2000 166.8000 222.6000 167.2000 ;
	    RECT 223.0000 166.8000 223.4000 167.2000 ;
	    RECT 227.0000 166.8000 227.4000 167.2000 ;
	    RECT 228.6000 167.1000 229.0000 167.2000 ;
	    RECT 229.4000 167.1000 229.8000 167.2000 ;
	    RECT 228.6000 166.8000 229.8000 167.1000 ;
	    RECT 231.8000 167.1000 232.2000 167.2000 ;
	    RECT 232.6000 167.1000 233.0000 167.2000 ;
	    RECT 231.8000 166.8000 233.0000 167.1000 ;
	    RECT 235.8000 166.8000 236.2000 167.2000 ;
	    RECT 236.6000 166.8000 237.0000 167.2000 ;
	    RECT 239.0000 166.8000 239.4000 167.2000 ;
	    RECT 240.6000 166.8000 241.0000 167.2000 ;
	    RECT 244.6000 167.1000 245.0000 167.2000 ;
	    RECT 245.4000 167.1000 245.8000 167.2000 ;
	    RECT 244.6000 166.8000 245.8000 167.1000 ;
	    RECT 246.2000 167.1000 246.6000 167.2000 ;
	    RECT 246.2000 166.8000 247.3000 167.1000 ;
	    RECT 219.8000 165.8000 220.2000 166.2000 ;
	    RECT 219.8000 163.2000 220.1000 165.8000 ;
	    RECT 219.8000 162.8000 220.2000 163.2000 ;
	    RECT 219.0000 161.8000 219.4000 162.2000 ;
	    RECT 219.8000 161.8000 220.2000 162.2000 ;
	    RECT 210.2000 160.8000 210.6000 161.2000 ;
	    RECT 211.0000 158.1000 211.4000 158.2000 ;
	    RECT 211.8000 158.1000 212.2000 158.2000 ;
	    RECT 205.4000 152.8000 205.8000 153.2000 ;
	    RECT 207.0000 152.8000 207.4000 153.2000 ;
	    RECT 203.8000 147.8000 204.2000 148.2000 ;
	    RECT 203.0000 146.8000 203.4000 147.2000 ;
	    RECT 203.8000 146.3000 204.1000 147.8000 ;
	    RECT 203.8000 145.9000 204.2000 146.3000 ;
	    RECT 204.6000 143.1000 205.0000 148.9000 ;
	    RECT 207.0000 148.2000 207.3000 152.8000 ;
	    RECT 208.6000 152.1000 209.0000 157.9000 ;
	    RECT 211.0000 157.8000 212.2000 158.1000 ;
	    RECT 217.4000 157.1000 217.8000 157.2000 ;
	    RECT 218.2000 157.1000 218.6000 157.2000 ;
	    RECT 217.4000 156.8000 218.6000 157.1000 ;
	    RECT 219.8000 156.2000 220.1000 161.8000 ;
	    RECT 222.2000 159.2000 222.5000 166.8000 ;
	    RECT 223.0000 165.2000 223.3000 166.8000 ;
	    RECT 227.0000 166.2000 227.3000 166.8000 ;
	    RECT 235.8000 166.2000 236.1000 166.8000 ;
	    RECT 236.6000 166.2000 236.9000 166.8000 ;
	    RECT 227.0000 165.8000 227.4000 166.2000 ;
	    RECT 227.8000 165.8000 228.2000 166.2000 ;
	    RECT 229.4000 165.8000 229.8000 166.2000 ;
	    RECT 230.2000 165.8000 230.6000 166.2000 ;
	    RECT 231.0000 165.8000 231.4000 166.2000 ;
	    RECT 233.4000 165.8000 233.8000 166.2000 ;
	    RECT 235.8000 165.8000 236.2000 166.2000 ;
	    RECT 236.6000 165.8000 237.0000 166.2000 ;
	    RECT 239.8000 165.8000 240.2000 166.2000 ;
	    RECT 227.8000 165.2000 228.1000 165.8000 ;
	    RECT 223.0000 164.8000 223.4000 165.2000 ;
	    RECT 224.6000 164.8000 225.0000 165.2000 ;
	    RECT 227.8000 164.8000 228.2000 165.2000 ;
	    RECT 224.6000 162.2000 224.9000 164.8000 ;
	    RECT 229.4000 162.2000 229.7000 165.8000 ;
	    RECT 230.2000 165.2000 230.5000 165.8000 ;
	    RECT 231.0000 165.2000 231.3000 165.8000 ;
	    RECT 230.2000 164.8000 230.6000 165.2000 ;
	    RECT 231.0000 164.8000 231.4000 165.2000 ;
	    RECT 224.6000 161.8000 225.0000 162.2000 ;
	    RECT 229.4000 161.8000 229.8000 162.2000 ;
	    RECT 231.0000 161.8000 231.4000 162.2000 ;
	    RECT 229.4000 160.8000 229.8000 161.2000 ;
	    RECT 223.0000 159.8000 223.4000 160.2000 ;
	    RECT 222.2000 158.8000 222.6000 159.2000 ;
	    RECT 222.2000 156.8000 222.6000 157.2000 ;
	    RECT 215.8000 155.8000 216.2000 156.2000 ;
	    RECT 219.8000 155.8000 220.2000 156.2000 ;
	    RECT 221.4000 155.8000 221.8000 156.2000 ;
	    RECT 214.2000 155.1000 214.6000 155.2000 ;
	    RECT 215.0000 155.1000 215.4000 155.2000 ;
	    RECT 214.2000 154.8000 215.4000 155.1000 ;
	    RECT 213.4000 152.8000 213.8000 153.2000 ;
	    RECT 213.4000 152.2000 213.7000 152.8000 ;
	    RECT 213.4000 151.8000 213.8000 152.2000 ;
	    RECT 214.2000 149.2000 214.5000 154.8000 ;
	    RECT 215.8000 154.2000 216.1000 155.8000 ;
	    RECT 219.8000 155.2000 220.1000 155.8000 ;
	    RECT 221.4000 155.2000 221.7000 155.8000 ;
	    RECT 222.2000 155.2000 222.5000 156.8000 ;
	    RECT 218.2000 154.8000 218.6000 155.2000 ;
	    RECT 219.0000 154.8000 219.4000 155.2000 ;
	    RECT 219.8000 154.8000 220.2000 155.2000 ;
	    RECT 221.4000 154.8000 221.8000 155.2000 ;
	    RECT 222.2000 154.8000 222.6000 155.2000 ;
	    RECT 218.2000 154.2000 218.5000 154.8000 ;
	    RECT 219.0000 154.2000 219.3000 154.8000 ;
	    RECT 215.8000 153.8000 216.2000 154.2000 ;
	    RECT 218.2000 153.8000 218.6000 154.2000 ;
	    RECT 219.0000 153.8000 219.4000 154.2000 ;
	    RECT 220.6000 154.1000 221.0000 154.2000 ;
	    RECT 221.4000 154.1000 221.8000 154.2000 ;
	    RECT 220.6000 153.8000 221.8000 154.1000 ;
	    RECT 222.2000 154.1000 222.6000 154.2000 ;
	    RECT 223.0000 154.1000 223.3000 159.8000 ;
	    RECT 227.8000 155.8000 228.2000 156.2000 ;
	    RECT 227.8000 155.2000 228.1000 155.8000 ;
	    RECT 229.4000 155.2000 229.7000 160.8000 ;
	    RECT 231.0000 159.2000 231.3000 161.8000 ;
	    RECT 233.4000 159.2000 233.7000 165.8000 ;
	    RECT 234.2000 165.1000 234.6000 165.2000 ;
	    RECT 235.0000 165.1000 235.4000 165.2000 ;
	    RECT 234.2000 164.8000 235.4000 165.1000 ;
	    RECT 235.8000 164.2000 236.1000 165.8000 ;
	    RECT 239.8000 165.2000 240.1000 165.8000 ;
	    RECT 236.6000 165.1000 237.0000 165.2000 ;
	    RECT 237.4000 165.1000 237.8000 165.2000 ;
	    RECT 236.6000 164.8000 237.8000 165.1000 ;
	    RECT 238.2000 164.8000 238.6000 165.2000 ;
	    RECT 239.8000 164.8000 240.2000 165.2000 ;
	    RECT 238.2000 164.2000 238.5000 164.8000 ;
	    RECT 235.8000 163.8000 236.2000 164.2000 ;
	    RECT 238.2000 163.8000 238.6000 164.2000 ;
	    RECT 231.0000 158.8000 231.4000 159.2000 ;
	    RECT 233.4000 158.8000 233.8000 159.2000 ;
	    RECT 235.0000 157.8000 235.4000 158.2000 ;
	    RECT 222.2000 153.8000 223.3000 154.1000 ;
	    RECT 227.0000 154.8000 227.4000 155.2000 ;
	    RECT 227.8000 154.8000 228.2000 155.2000 ;
	    RECT 229.4000 154.8000 229.8000 155.2000 ;
	    RECT 234.2000 154.8000 234.6000 155.2000 ;
	    RECT 215.8000 153.1000 216.2000 153.2000 ;
	    RECT 216.6000 153.1000 217.0000 153.2000 ;
	    RECT 226.2000 153.1000 226.6000 153.2000 ;
	    RECT 215.8000 152.8000 217.0000 153.1000 ;
	    RECT 225.4000 152.8000 226.6000 153.1000 ;
	    RECT 224.6000 151.8000 225.0000 152.2000 ;
	    RECT 224.6000 150.2000 224.9000 151.8000 ;
	    RECT 218.2000 149.8000 218.6000 150.2000 ;
	    RECT 224.6000 149.8000 225.0000 150.2000 ;
	    RECT 214.2000 148.8000 214.6000 149.2000 ;
	    RECT 206.2000 145.1000 206.6000 147.9000 ;
	    RECT 207.0000 147.8000 207.4000 148.2000 ;
	    RECT 207.8000 148.1000 208.2000 148.2000 ;
	    RECT 208.6000 148.1000 209.0000 148.2000 ;
	    RECT 207.8000 147.8000 209.0000 148.1000 ;
	    RECT 211.8000 147.8000 212.2000 148.2000 ;
	    RECT 216.6000 147.8000 217.0000 148.2000 ;
	    RECT 211.8000 147.2000 212.1000 147.8000 ;
	    RECT 211.8000 146.8000 212.2000 147.2000 ;
	    RECT 212.6000 147.1000 213.0000 147.2000 ;
	    RECT 213.4000 147.1000 213.8000 147.2000 ;
	    RECT 212.6000 146.8000 213.8000 147.1000 ;
	    RECT 214.2000 146.8000 214.6000 147.2000 ;
	    RECT 214.2000 146.2000 214.5000 146.8000 ;
	    RECT 208.6000 146.1000 209.0000 146.2000 ;
	    RECT 209.4000 146.1000 209.8000 146.2000 ;
	    RECT 208.6000 145.8000 209.8000 146.1000 ;
	    RECT 214.2000 145.8000 214.6000 146.2000 ;
	    RECT 216.6000 145.2000 216.9000 147.8000 ;
	    RECT 218.2000 147.2000 218.5000 149.8000 ;
	    RECT 223.0000 148.8000 223.4000 149.2000 ;
	    RECT 223.0000 147.2000 223.3000 148.8000 ;
	    RECT 225.4000 147.2000 225.7000 152.8000 ;
	    RECT 227.0000 152.2000 227.3000 154.8000 ;
	    RECT 228.6000 153.1000 229.0000 153.2000 ;
	    RECT 229.4000 153.1000 229.8000 153.2000 ;
	    RECT 228.6000 152.8000 229.8000 153.1000 ;
	    RECT 232.6000 152.8000 233.0000 153.2000 ;
	    RECT 227.0000 151.8000 227.4000 152.2000 ;
	    RECT 226.2000 148.8000 226.6000 149.2000 ;
	    RECT 226.2000 148.2000 226.5000 148.8000 ;
	    RECT 226.2000 147.8000 226.6000 148.2000 ;
	    RECT 218.2000 146.8000 218.6000 147.2000 ;
	    RECT 223.0000 146.8000 223.4000 147.2000 ;
	    RECT 225.4000 146.8000 225.8000 147.2000 ;
	    RECT 220.6000 145.8000 221.0000 146.2000 ;
	    RECT 221.4000 145.8000 221.8000 146.2000 ;
	    RECT 222.2000 145.8000 222.6000 146.2000 ;
	    RECT 223.0000 146.1000 223.4000 146.2000 ;
	    RECT 223.8000 146.1000 224.2000 146.2000 ;
	    RECT 223.0000 145.8000 224.2000 146.1000 ;
	    RECT 220.6000 145.2000 220.9000 145.8000 ;
	    RECT 210.2000 144.8000 210.6000 145.2000 ;
	    RECT 216.6000 144.8000 217.0000 145.2000 ;
	    RECT 220.6000 144.8000 221.0000 145.2000 ;
	    RECT 210.2000 143.2000 210.5000 144.8000 ;
	    RECT 216.6000 143.8000 217.0000 144.2000 ;
	    RECT 210.2000 142.8000 210.6000 143.2000 ;
	    RECT 214.2000 141.8000 214.6000 142.2000 ;
	    RECT 201.4000 140.8000 201.8000 141.2000 ;
	    RECT 202.2000 139.8000 202.6000 140.2000 ;
	    RECT 202.2000 139.2000 202.5000 139.8000 ;
	    RECT 202.2000 138.8000 202.6000 139.2000 ;
	    RECT 207.8000 138.8000 208.2000 139.2000 ;
	    RECT 195.0000 138.1000 195.4000 138.2000 ;
	    RECT 195.8000 138.1000 196.2000 138.2000 ;
	    RECT 195.0000 137.8000 196.2000 138.1000 ;
	    RECT 201.4000 137.8000 201.8000 138.2000 ;
	    RECT 194.2000 136.8000 194.6000 137.2000 ;
	    RECT 198.2000 137.1000 198.6000 137.2000 ;
	    RECT 199.0000 137.1000 199.4000 137.2000 ;
	    RECT 198.2000 136.8000 199.4000 137.1000 ;
	    RECT 199.8000 137.1000 200.2000 137.2000 ;
	    RECT 200.6000 137.1000 201.0000 137.2000 ;
	    RECT 199.8000 136.8000 201.0000 137.1000 ;
	    RECT 194.2000 135.2000 194.5000 136.8000 ;
	    RECT 201.4000 136.2000 201.7000 137.8000 ;
	    RECT 206.2000 136.8000 206.6000 137.2000 ;
	    RECT 206.2000 136.2000 206.5000 136.8000 ;
	    RECT 207.8000 136.2000 208.1000 138.8000 ;
	    RECT 210.2000 136.8000 210.6000 137.2000 ;
	    RECT 195.8000 136.1000 196.2000 136.2000 ;
	    RECT 196.6000 136.1000 197.0000 136.2000 ;
	    RECT 195.8000 135.8000 197.0000 136.1000 ;
	    RECT 201.4000 135.8000 201.8000 136.2000 ;
	    RECT 203.8000 135.8000 204.2000 136.2000 ;
	    RECT 206.2000 135.8000 206.6000 136.2000 ;
	    RECT 207.8000 135.8000 208.2000 136.2000 ;
	    RECT 194.2000 134.8000 194.6000 135.2000 ;
	    RECT 195.8000 135.1000 196.2000 135.2000 ;
	    RECT 196.6000 135.1000 197.0000 135.2000 ;
	    RECT 195.8000 134.8000 197.0000 135.1000 ;
	    RECT 197.4000 134.8000 197.8000 135.2000 ;
	    RECT 198.2000 134.8000 198.6000 135.2000 ;
	    RECT 194.2000 134.2000 194.5000 134.8000 ;
	    RECT 197.4000 134.2000 197.7000 134.8000 ;
	    RECT 198.2000 134.2000 198.5000 134.8000 ;
	    RECT 192.6000 134.1000 193.0000 134.2000 ;
	    RECT 193.4000 134.1000 193.8000 134.2000 ;
	    RECT 192.6000 133.8000 193.8000 134.1000 ;
	    RECT 194.2000 133.8000 194.6000 134.2000 ;
	    RECT 197.4000 133.8000 197.8000 134.2000 ;
	    RECT 198.2000 133.8000 198.6000 134.2000 ;
	    RECT 191.0000 130.8000 191.4000 131.2000 ;
	    RECT 191.8000 130.8000 192.2000 131.2000 ;
	    RECT 191.0000 129.2000 191.3000 130.8000 ;
	    RECT 193.4000 129.2000 193.7000 133.8000 ;
	    RECT 194.2000 132.8000 194.6000 133.2000 ;
	    RECT 194.2000 131.2000 194.5000 132.8000 ;
	    RECT 194.2000 130.8000 194.6000 131.2000 ;
	    RECT 191.0000 128.8000 191.4000 129.2000 ;
	    RECT 193.4000 128.8000 193.8000 129.2000 ;
	    RECT 191.8000 127.8000 192.2000 128.2000 ;
	    RECT 195.0000 127.8000 195.4000 128.2000 ;
	    RECT 191.8000 127.2000 192.1000 127.8000 ;
	    RECT 191.8000 126.8000 192.2000 127.2000 ;
	    RECT 193.4000 126.1000 193.8000 126.2000 ;
	    RECT 194.2000 126.1000 194.6000 126.2000 ;
	    RECT 193.4000 125.8000 194.6000 126.1000 ;
	    RECT 195.0000 125.2000 195.3000 127.8000 ;
	    RECT 197.4000 126.2000 197.7000 133.8000 ;
	    RECT 203.8000 133.2000 204.1000 135.8000 ;
	    RECT 206.2000 134.8000 206.6000 135.2000 ;
	    RECT 209.4000 134.8000 209.8000 135.2000 ;
	    RECT 200.6000 133.1000 201.0000 133.2000 ;
	    RECT 201.4000 133.1000 201.8000 133.2000 ;
	    RECT 200.6000 132.8000 201.8000 133.1000 ;
	    RECT 203.8000 132.8000 204.2000 133.2000 ;
	    RECT 205.4000 132.8000 205.8000 133.2000 ;
	    RECT 197.4000 125.8000 197.8000 126.2000 ;
	    RECT 190.2000 124.8000 191.3000 125.1000 ;
	    RECT 195.0000 124.8000 195.4000 125.2000 ;
	    RECT 189.4000 124.1000 189.8000 124.2000 ;
	    RECT 190.2000 124.1000 190.6000 124.2000 ;
	    RECT 189.4000 123.8000 190.6000 124.1000 ;
	    RECT 187.8000 112.1000 188.2000 117.9000 ;
	    RECT 191.0000 117.2000 191.3000 124.8000 ;
	    RECT 192.6000 124.1000 193.0000 124.2000 ;
	    RECT 193.4000 124.1000 193.8000 124.2000 ;
	    RECT 192.6000 123.8000 193.8000 124.1000 ;
	    RECT 198.2000 123.1000 198.6000 128.9000 ;
	    RECT 199.0000 125.8000 199.4000 126.2000 ;
	    RECT 202.2000 125.9000 202.6000 126.3000 ;
	    RECT 194.2000 121.8000 194.6000 122.2000 ;
	    RECT 195.8000 121.8000 196.2000 122.2000 ;
	    RECT 199.0000 122.1000 199.3000 125.8000 ;
	    RECT 202.2000 125.2000 202.5000 125.9000 ;
	    RECT 202.2000 124.8000 202.6000 125.2000 ;
	    RECT 203.0000 123.1000 203.4000 128.9000 ;
	    RECT 198.2000 121.8000 199.3000 122.1000 ;
	    RECT 191.0000 116.8000 191.4000 117.2000 ;
	    RECT 191.0000 113.1000 191.4000 115.9000 ;
	    RECT 191.8000 115.8000 192.2000 116.2000 ;
	    RECT 191.8000 114.2000 192.1000 115.8000 ;
	    RECT 191.8000 113.8000 192.2000 114.2000 ;
	    RECT 191.8000 112.8000 192.2000 113.2000 ;
	    RECT 189.4000 112.1000 189.8000 112.2000 ;
	    RECT 190.2000 112.1000 190.6000 112.2000 ;
	    RECT 189.4000 111.8000 190.6000 112.1000 ;
	    RECT 187.0000 110.8000 187.4000 111.2000 ;
	    RECT 191.8000 109.2000 192.1000 112.8000 ;
	    RECT 192.6000 112.1000 193.0000 117.9000 ;
	    RECT 194.2000 116.2000 194.5000 121.8000 ;
	    RECT 194.2000 115.8000 194.6000 116.2000 ;
	    RECT 193.4000 114.7000 193.8000 115.1000 ;
	    RECT 193.4000 113.2000 193.7000 114.7000 ;
	    RECT 193.4000 112.8000 193.8000 113.2000 ;
	    RECT 191.0000 108.8000 191.4000 109.2000 ;
	    RECT 191.8000 108.8000 192.2000 109.2000 ;
	    RECT 191.0000 108.2000 191.3000 108.8000 ;
	    RECT 186.2000 107.5000 186.6000 107.9000 ;
	    RECT 186.9000 107.5000 189.0000 107.8000 ;
	    RECT 189.5000 107.5000 189.9000 107.9000 ;
	    RECT 191.0000 107.8000 191.4000 108.2000 ;
	    RECT 192.6000 107.8000 193.0000 108.2000 ;
	    RECT 185.4000 106.8000 185.8000 107.2000 ;
	    RECT 186.2000 107.1000 186.5000 107.5000 ;
	    RECT 186.9000 107.4000 187.3000 107.5000 ;
	    RECT 188.6000 107.4000 189.0000 107.5000 ;
	    RECT 186.2000 106.8000 188.6000 107.1000 ;
	    RECT 184.6000 105.8000 185.0000 106.2000 ;
	    RECT 183.8000 93.8000 184.2000 94.2000 ;
	    RECT 181.4000 92.8000 181.8000 93.2000 ;
	    RECT 183.8000 91.2000 184.1000 93.8000 ;
	    RECT 179.8000 90.8000 180.2000 91.2000 ;
	    RECT 183.8000 90.8000 184.2000 91.2000 ;
	    RECT 175.8000 89.8000 176.2000 90.2000 ;
	    RECT 175.0000 87.8000 175.4000 88.2000 ;
	    RECT 175.8000 86.2000 176.1000 89.8000 ;
	    RECT 175.8000 85.8000 176.2000 86.2000 ;
	    RECT 179.0000 83.1000 179.4000 88.9000 ;
	    RECT 179.8000 85.2000 180.1000 90.8000 ;
	    RECT 181.4000 88.8000 181.8000 89.2000 ;
	    RECT 182.2000 88.8000 182.6000 89.2000 ;
	    RECT 183.0000 88.8000 183.4000 89.2000 ;
	    RECT 181.4000 88.2000 181.7000 88.8000 ;
	    RECT 182.2000 88.2000 182.5000 88.8000 ;
	    RECT 183.0000 88.2000 183.3000 88.8000 ;
	    RECT 181.4000 87.8000 181.8000 88.2000 ;
	    RECT 182.2000 87.8000 182.6000 88.2000 ;
	    RECT 183.0000 87.8000 183.4000 88.2000 ;
	    RECT 183.8000 88.1000 184.2000 88.2000 ;
	    RECT 184.6000 88.1000 184.9000 105.8000 ;
	    RECT 186.2000 105.1000 186.5000 106.8000 ;
	    RECT 188.2000 106.7000 188.6000 106.8000 ;
	    RECT 189.6000 105.1000 189.9000 107.5000 ;
	    RECT 192.6000 107.2000 192.9000 107.8000 ;
	    RECT 194.2000 107.2000 194.5000 115.8000 ;
	    RECT 195.8000 115.2000 196.1000 121.8000 ;
	    RECT 195.8000 114.8000 196.2000 115.2000 ;
	    RECT 196.6000 113.8000 197.0000 114.2000 ;
	    RECT 190.2000 107.1000 190.6000 107.2000 ;
	    RECT 191.0000 107.1000 191.4000 107.2000 ;
	    RECT 190.2000 106.8000 191.4000 107.1000 ;
	    RECT 192.6000 106.8000 193.0000 107.2000 ;
	    RECT 194.2000 106.8000 194.6000 107.2000 ;
	    RECT 186.2000 104.7000 186.6000 105.1000 ;
	    RECT 189.5000 104.7000 189.9000 105.1000 ;
	    RECT 193.4000 105.8000 193.8000 106.2000 ;
	    RECT 193.4000 105.2000 193.7000 105.8000 ;
	    RECT 193.4000 104.8000 193.8000 105.2000 ;
	    RECT 187.8000 104.1000 188.2000 104.2000 ;
	    RECT 188.6000 104.1000 189.0000 104.2000 ;
	    RECT 187.8000 103.8000 189.0000 104.1000 ;
	    RECT 186.2000 97.8000 186.6000 98.2000 ;
	    RECT 191.8000 97.8000 192.2000 98.2000 ;
	    RECT 185.4000 96.8000 185.8000 97.2000 ;
	    RECT 185.4000 96.2000 185.7000 96.8000 ;
	    RECT 185.4000 95.8000 185.8000 96.2000 ;
	    RECT 186.2000 94.2000 186.5000 97.8000 ;
	    RECT 187.0000 96.8000 187.4000 97.2000 ;
	    RECT 187.0000 96.2000 187.3000 96.8000 ;
	    RECT 187.0000 95.8000 187.4000 96.2000 ;
	    RECT 187.0000 94.8000 187.4000 95.2000 ;
	    RECT 190.2000 94.8000 190.6000 95.2000 ;
	    RECT 186.2000 93.8000 186.6000 94.2000 ;
	    RECT 186.2000 92.8000 186.6000 93.2000 ;
	    RECT 185.4000 91.8000 185.8000 92.2000 ;
	    RECT 185.4000 91.2000 185.7000 91.8000 ;
	    RECT 185.4000 90.8000 185.8000 91.2000 ;
	    RECT 186.2000 89.2000 186.5000 92.8000 ;
	    RECT 187.0000 90.2000 187.3000 94.8000 ;
	    RECT 189.4000 93.8000 189.8000 94.2000 ;
	    RECT 188.6000 90.8000 189.0000 91.2000 ;
	    RECT 187.0000 89.8000 187.4000 90.2000 ;
	    RECT 186.2000 88.8000 186.6000 89.2000 ;
	    RECT 187.8000 88.8000 188.2000 89.2000 ;
	    RECT 183.8000 87.8000 184.9000 88.1000 ;
	    RECT 181.4000 86.2000 181.7000 87.8000 ;
	    RECT 187.8000 87.2000 188.1000 88.8000 ;
	    RECT 188.6000 88.2000 188.9000 90.8000 ;
	    RECT 189.4000 89.2000 189.7000 93.8000 ;
	    RECT 190.2000 93.2000 190.5000 94.8000 ;
	    RECT 190.2000 92.8000 190.6000 93.2000 ;
	    RECT 191.0000 93.1000 191.4000 95.9000 ;
	    RECT 189.4000 88.8000 189.8000 89.2000 ;
	    RECT 190.2000 88.8000 190.6000 89.2000 ;
	    RECT 188.6000 87.8000 189.0000 88.2000 ;
	    RECT 190.2000 87.2000 190.5000 88.8000 ;
	    RECT 191.8000 87.2000 192.1000 97.8000 ;
	    RECT 192.6000 92.1000 193.0000 97.9000 ;
	    RECT 193.4000 89.8000 193.8000 90.2000 ;
	    RECT 193.4000 88.2000 193.7000 89.8000 ;
	    RECT 193.4000 87.8000 193.8000 88.2000 ;
	    RECT 194.2000 87.2000 194.5000 106.8000 ;
	    RECT 195.0000 106.1000 195.4000 106.2000 ;
	    RECT 195.8000 106.1000 196.2000 106.2000 ;
	    RECT 195.0000 105.8000 196.2000 106.1000 ;
	    RECT 195.0000 105.1000 195.4000 105.2000 ;
	    RECT 195.8000 105.1000 196.2000 105.2000 ;
	    RECT 195.0000 104.8000 196.2000 105.1000 ;
	    RECT 196.6000 95.2000 196.9000 113.8000 ;
	    RECT 197.4000 112.1000 197.8000 117.9000 ;
	    RECT 198.2000 117.2000 198.5000 121.8000 ;
	    RECT 198.2000 116.8000 198.6000 117.2000 ;
	    RECT 200.6000 114.8000 201.0000 115.2000 ;
	    RECT 200.6000 114.2000 200.9000 114.8000 ;
	    RECT 200.6000 113.8000 201.0000 114.2000 ;
	    RECT 203.8000 113.2000 204.1000 132.8000 ;
	    RECT 205.4000 128.2000 205.7000 132.8000 ;
	    RECT 206.2000 129.2000 206.5000 134.8000 ;
	    RECT 208.6000 133.8000 209.0000 134.2000 ;
	    RECT 208.6000 133.2000 208.9000 133.8000 ;
	    RECT 207.0000 133.1000 207.4000 133.2000 ;
	    RECT 207.8000 133.1000 208.2000 133.2000 ;
	    RECT 207.0000 132.8000 208.2000 133.1000 ;
	    RECT 208.6000 132.8000 209.0000 133.2000 ;
	    RECT 206.2000 128.8000 206.6000 129.2000 ;
	    RECT 209.4000 129.1000 209.7000 134.8000 ;
	    RECT 210.2000 134.2000 210.5000 136.8000 ;
	    RECT 214.2000 134.2000 214.5000 141.8000 ;
	    RECT 216.6000 139.2000 216.9000 143.8000 ;
	    RECT 219.8000 141.8000 220.2000 142.2000 ;
	    RECT 216.6000 138.8000 217.0000 139.2000 ;
	    RECT 219.0000 138.8000 219.4000 139.2000 ;
	    RECT 219.0000 138.2000 219.3000 138.8000 ;
	    RECT 219.0000 137.8000 219.4000 138.2000 ;
	    RECT 219.8000 137.2000 220.1000 141.8000 ;
	    RECT 221.4000 139.2000 221.7000 145.8000 ;
	    RECT 222.2000 145.1000 222.5000 145.8000 ;
	    RECT 222.2000 144.8000 223.3000 145.1000 ;
	    RECT 223.0000 139.2000 223.3000 144.8000 ;
	    RECT 223.8000 144.8000 224.2000 145.2000 ;
	    RECT 223.8000 144.2000 224.1000 144.8000 ;
	    RECT 227.0000 144.2000 227.3000 151.8000 ;
	    RECT 228.6000 149.2000 228.9000 152.8000 ;
	    RECT 232.6000 149.2000 232.9000 152.8000 ;
	    RECT 228.6000 148.8000 229.0000 149.2000 ;
	    RECT 230.2000 148.8000 230.6000 149.2000 ;
	    RECT 232.6000 148.8000 233.0000 149.2000 ;
	    RECT 230.2000 148.2000 230.5000 148.8000 ;
	    RECT 230.2000 147.8000 230.6000 148.2000 ;
	    RECT 228.6000 147.1000 229.0000 147.2000 ;
	    RECT 229.4000 147.1000 229.8000 147.2000 ;
	    RECT 228.6000 146.8000 229.8000 147.1000 ;
	    RECT 227.8000 145.8000 228.2000 146.2000 ;
	    RECT 228.6000 145.8000 229.0000 146.2000 ;
	    RECT 230.2000 146.1000 230.5000 147.8000 ;
	    RECT 233.4000 146.8000 233.8000 147.2000 ;
	    RECT 233.4000 146.2000 233.7000 146.8000 ;
	    RECT 229.4000 145.8000 230.5000 146.1000 ;
	    RECT 231.0000 146.1000 231.4000 146.2000 ;
	    RECT 231.8000 146.1000 232.2000 146.2000 ;
	    RECT 231.0000 145.8000 232.2000 146.1000 ;
	    RECT 233.4000 145.8000 233.8000 146.2000 ;
	    RECT 227.8000 145.2000 228.1000 145.8000 ;
	    RECT 228.6000 145.2000 228.9000 145.8000 ;
	    RECT 227.8000 144.8000 228.2000 145.2000 ;
	    RECT 228.6000 144.8000 229.0000 145.2000 ;
	    RECT 223.8000 143.8000 224.2000 144.2000 ;
	    RECT 227.0000 143.8000 227.4000 144.2000 ;
	    RECT 227.8000 143.8000 228.2000 144.2000 ;
	    RECT 227.8000 139.2000 228.1000 143.8000 ;
	    RECT 221.4000 138.8000 221.8000 139.2000 ;
	    RECT 223.0000 138.8000 223.4000 139.2000 ;
	    RECT 227.8000 138.8000 228.2000 139.2000 ;
	    RECT 219.8000 136.8000 220.2000 137.2000 ;
	    RECT 228.6000 136.8000 229.0000 137.2000 ;
	    RECT 228.6000 136.2000 228.9000 136.8000 ;
	    RECT 217.4000 135.8000 217.8000 136.2000 ;
	    RECT 219.8000 135.8000 220.2000 136.2000 ;
	    RECT 222.2000 135.8000 222.6000 136.2000 ;
	    RECT 227.0000 136.1000 227.4000 136.2000 ;
	    RECT 227.0000 135.8000 228.1000 136.1000 ;
	    RECT 217.4000 135.2000 217.7000 135.8000 ;
	    RECT 219.8000 135.2000 220.1000 135.8000 ;
	    RECT 215.0000 134.8000 215.4000 135.2000 ;
	    RECT 217.4000 134.8000 217.8000 135.2000 ;
	    RECT 219.8000 134.8000 220.2000 135.2000 ;
	    RECT 220.6000 134.8000 221.0000 135.2000 ;
	    RECT 210.2000 133.8000 210.6000 134.2000 ;
	    RECT 214.2000 133.8000 214.6000 134.2000 ;
	    RECT 215.0000 133.2000 215.3000 134.8000 ;
	    RECT 219.8000 134.2000 220.1000 134.8000 ;
	    RECT 215.8000 133.8000 216.2000 134.2000 ;
	    RECT 218.2000 133.8000 218.6000 134.2000 ;
	    RECT 219.8000 133.8000 220.2000 134.2000 ;
	    RECT 211.8000 133.1000 212.2000 133.2000 ;
	    RECT 212.6000 133.1000 213.0000 133.2000 ;
	    RECT 211.8000 132.8000 213.0000 133.1000 ;
	    RECT 213.4000 132.8000 213.8000 133.2000 ;
	    RECT 215.0000 132.8000 215.4000 133.2000 ;
	    RECT 213.4000 132.2000 213.7000 132.8000 ;
	    RECT 213.4000 131.8000 213.8000 132.2000 ;
	    RECT 209.4000 128.8000 210.5000 129.1000 ;
	    RECT 204.6000 125.1000 205.0000 127.9000 ;
	    RECT 205.4000 127.8000 205.8000 128.2000 ;
	    RECT 207.8000 127.8000 208.2000 128.2000 ;
	    RECT 207.8000 127.2000 208.1000 127.8000 ;
	    RECT 207.8000 126.8000 208.2000 127.2000 ;
	    RECT 208.6000 127.1000 209.0000 127.2000 ;
	    RECT 209.4000 127.1000 209.8000 127.2000 ;
	    RECT 208.6000 126.8000 209.8000 127.1000 ;
	    RECT 207.0000 125.8000 207.4000 126.2000 ;
	    RECT 208.6000 125.8000 209.0000 126.2000 ;
	    RECT 207.0000 124.2000 207.3000 125.8000 ;
	    RECT 208.6000 125.2000 208.9000 125.8000 ;
	    RECT 208.6000 124.8000 209.0000 125.2000 ;
	    RECT 207.0000 123.8000 207.4000 124.2000 ;
	    RECT 210.2000 121.2000 210.5000 128.8000 ;
	    RECT 211.0000 127.8000 211.4000 128.2000 ;
	    RECT 214.2000 128.1000 214.6000 128.2000 ;
	    RECT 215.0000 128.1000 215.4000 128.2000 ;
	    RECT 214.2000 127.8000 215.4000 128.1000 ;
	    RECT 211.0000 127.2000 211.3000 127.8000 ;
	    RECT 211.0000 126.8000 211.4000 127.2000 ;
	    RECT 215.0000 127.1000 215.4000 127.2000 ;
	    RECT 215.8000 127.1000 216.1000 133.8000 ;
	    RECT 218.2000 131.2000 218.5000 133.8000 ;
	    RECT 219.0000 132.8000 219.4000 133.2000 ;
	    RECT 218.2000 130.8000 218.6000 131.2000 ;
	    RECT 216.6000 128.1000 217.0000 128.2000 ;
	    RECT 217.4000 128.1000 217.8000 128.2000 ;
	    RECT 216.6000 127.8000 217.8000 128.1000 ;
	    RECT 215.0000 126.8000 216.1000 127.1000 ;
	    RECT 217.4000 127.1000 217.8000 127.2000 ;
	    RECT 218.2000 127.1000 218.5000 130.8000 ;
	    RECT 217.4000 126.8000 218.5000 127.1000 ;
	    RECT 211.8000 126.1000 212.2000 126.2000 ;
	    RECT 212.6000 126.1000 213.0000 126.2000 ;
	    RECT 211.8000 125.8000 213.0000 126.1000 ;
	    RECT 214.2000 125.8000 214.6000 126.2000 ;
	    RECT 215.8000 126.1000 216.2000 126.2000 ;
	    RECT 216.6000 126.1000 217.0000 126.2000 ;
	    RECT 215.8000 125.8000 217.0000 126.1000 ;
	    RECT 218.2000 126.1000 218.6000 126.2000 ;
	    RECT 219.0000 126.1000 219.3000 132.8000 ;
	    RECT 220.6000 128.2000 220.9000 134.8000 ;
	    RECT 222.2000 133.2000 222.5000 135.8000 ;
	    RECT 224.6000 134.8000 225.0000 135.2000 ;
	    RECT 224.6000 134.2000 224.9000 134.8000 ;
	    RECT 224.6000 133.8000 225.0000 134.2000 ;
	    RECT 226.2000 134.1000 226.6000 134.2000 ;
	    RECT 227.0000 134.1000 227.4000 134.2000 ;
	    RECT 226.2000 133.8000 227.4000 134.1000 ;
	    RECT 222.2000 132.8000 222.6000 133.2000 ;
	    RECT 223.8000 132.8000 224.2000 133.2000 ;
	    RECT 220.6000 127.8000 221.0000 128.2000 ;
	    RECT 222.2000 127.2000 222.5000 132.8000 ;
	    RECT 223.8000 128.2000 224.1000 132.8000 ;
	    RECT 225.4000 132.1000 225.8000 132.2000 ;
	    RECT 226.2000 132.1000 226.6000 132.2000 ;
	    RECT 225.4000 131.8000 226.6000 132.1000 ;
	    RECT 223.0000 127.8000 223.4000 128.2000 ;
	    RECT 223.8000 127.8000 224.2000 128.2000 ;
	    RECT 222.2000 126.8000 222.6000 127.2000 ;
	    RECT 223.0000 126.2000 223.3000 127.8000 ;
	    RECT 227.0000 127.2000 227.3000 133.8000 ;
	    RECT 227.8000 133.1000 228.1000 135.8000 ;
	    RECT 228.6000 135.8000 229.0000 136.2000 ;
	    RECT 228.6000 134.2000 228.9000 135.8000 ;
	    RECT 228.6000 133.8000 229.0000 134.2000 ;
	    RECT 228.6000 133.1000 229.0000 133.2000 ;
	    RECT 227.8000 132.8000 229.0000 133.1000 ;
	    RECT 227.8000 131.8000 228.2000 132.2000 ;
	    RECT 225.4000 126.8000 225.8000 127.2000 ;
	    RECT 227.0000 126.8000 227.4000 127.2000 ;
	    RECT 225.4000 126.2000 225.7000 126.8000 ;
	    RECT 227.8000 126.2000 228.1000 131.8000 ;
	    RECT 228.6000 129.2000 228.9000 132.8000 ;
	    RECT 228.6000 128.8000 229.0000 129.2000 ;
	    RECT 228.6000 126.8000 229.0000 127.2000 ;
	    RECT 218.2000 125.8000 219.3000 126.1000 ;
	    RECT 219.8000 125.8000 220.2000 126.2000 ;
	    RECT 222.2000 125.8000 222.6000 126.2000 ;
	    RECT 223.0000 125.8000 223.4000 126.2000 ;
	    RECT 224.6000 125.8000 225.0000 126.2000 ;
	    RECT 225.4000 125.8000 225.8000 126.2000 ;
	    RECT 227.8000 125.8000 228.2000 126.2000 ;
	    RECT 214.2000 125.2000 214.5000 125.8000 ;
	    RECT 214.2000 124.8000 214.6000 125.2000 ;
	    RECT 219.8000 124.2000 220.1000 125.8000 ;
	    RECT 222.2000 124.2000 222.5000 125.8000 ;
	    RECT 224.6000 125.2000 224.9000 125.8000 ;
	    RECT 224.6000 124.8000 225.0000 125.2000 ;
	    RECT 226.2000 125.1000 226.6000 125.2000 ;
	    RECT 227.0000 125.1000 227.4000 125.2000 ;
	    RECT 226.2000 124.8000 227.4000 125.1000 ;
	    RECT 216.6000 123.8000 217.0000 124.2000 ;
	    RECT 219.8000 123.8000 220.2000 124.2000 ;
	    RECT 222.2000 123.8000 222.6000 124.2000 ;
	    RECT 213.4000 121.8000 213.8000 122.2000 ;
	    RECT 210.2000 120.8000 210.6000 121.2000 ;
	    RECT 213.4000 119.2000 213.7000 121.8000 ;
	    RECT 216.6000 119.2000 216.9000 123.8000 ;
	    RECT 223.8000 120.8000 224.2000 121.2000 ;
	    RECT 223.8000 119.2000 224.1000 120.8000 ;
	    RECT 213.4000 118.8000 213.8000 119.2000 ;
	    RECT 216.6000 118.8000 217.0000 119.2000 ;
	    RECT 223.8000 118.8000 224.2000 119.2000 ;
	    RECT 222.2000 116.8000 222.6000 117.2000 ;
	    RECT 222.2000 116.2000 222.5000 116.8000 ;
	    RECT 204.6000 115.8000 205.0000 116.2000 ;
	    RECT 215.0000 116.1000 215.4000 116.2000 ;
	    RECT 214.2000 115.8000 215.4000 116.1000 ;
	    RECT 218.2000 115.8000 218.6000 116.2000 ;
	    RECT 222.2000 115.8000 222.6000 116.2000 ;
	    RECT 204.6000 115.2000 204.9000 115.8000 ;
	    RECT 204.6000 114.8000 205.0000 115.2000 ;
	    RECT 207.8000 114.8000 208.2000 115.2000 ;
	    RECT 211.8000 115.1000 212.2000 115.2000 ;
	    RECT 212.6000 115.1000 213.0000 115.2000 ;
	    RECT 211.8000 114.8000 213.0000 115.1000 ;
	    RECT 203.8000 112.8000 204.2000 113.2000 ;
	    RECT 206.2000 112.8000 206.6000 113.2000 ;
	    RECT 199.8000 111.8000 200.2000 112.2000 ;
	    RECT 201.4000 111.8000 201.8000 112.2000 ;
	    RECT 204.6000 111.8000 205.0000 112.2000 ;
	    RECT 199.8000 111.2000 200.1000 111.8000 ;
	    RECT 197.4000 110.8000 197.8000 111.2000 ;
	    RECT 199.8000 110.8000 200.2000 111.2000 ;
	    RECT 197.4000 107.2000 197.7000 110.8000 ;
	    RECT 201.4000 109.2000 201.7000 111.8000 ;
	    RECT 204.6000 109.2000 204.9000 111.8000 ;
	    RECT 201.4000 108.8000 201.8000 109.2000 ;
	    RECT 204.6000 108.8000 205.0000 109.2000 ;
	    RECT 198.2000 107.5000 198.6000 107.9000 ;
	    RECT 198.9000 107.5000 201.0000 107.8000 ;
	    RECT 201.5000 107.5000 201.9000 107.9000 ;
	    RECT 197.4000 106.8000 197.8000 107.2000 ;
	    RECT 198.2000 107.1000 198.5000 107.5000 ;
	    RECT 198.9000 107.4000 199.3000 107.5000 ;
	    RECT 200.6000 107.4000 201.0000 107.5000 ;
	    RECT 198.2000 106.8000 200.6000 107.1000 ;
	    RECT 198.2000 105.1000 198.5000 106.8000 ;
	    RECT 200.2000 106.7000 200.6000 106.8000 ;
	    RECT 198.2000 104.7000 198.6000 105.1000 ;
	    RECT 200.6000 104.8000 201.0000 105.2000 ;
	    RECT 201.6000 105.1000 201.9000 107.5000 ;
	    RECT 202.2000 107.8000 202.6000 108.2000 ;
	    RECT 203.0000 107.8000 203.4000 108.2000 ;
	    RECT 203.8000 107.8000 204.2000 108.2000 ;
	    RECT 205.4000 107.8000 205.8000 108.2000 ;
	    RECT 202.2000 107.2000 202.5000 107.8000 ;
	    RECT 203.0000 107.2000 203.3000 107.8000 ;
	    RECT 202.2000 106.8000 202.6000 107.2000 ;
	    RECT 203.0000 106.8000 203.4000 107.2000 ;
	    RECT 200.6000 104.2000 200.9000 104.8000 ;
	    RECT 201.5000 104.7000 201.9000 105.1000 ;
	    RECT 200.6000 103.8000 201.0000 104.2000 ;
	    RECT 203.8000 99.2000 204.1000 107.8000 ;
	    RECT 205.4000 107.2000 205.7000 107.8000 ;
	    RECT 204.6000 106.8000 205.0000 107.2000 ;
	    RECT 205.4000 106.8000 205.8000 107.2000 ;
	    RECT 204.6000 105.2000 204.9000 106.8000 ;
	    RECT 206.2000 106.2000 206.5000 112.8000 ;
	    RECT 207.0000 111.8000 207.4000 112.2000 ;
	    RECT 207.0000 110.2000 207.3000 111.8000 ;
	    RECT 207.0000 109.8000 207.4000 110.2000 ;
	    RECT 207.8000 109.2000 208.1000 114.8000 ;
	    RECT 209.4000 114.1000 209.8000 114.2000 ;
	    RECT 209.4000 113.8000 210.5000 114.1000 ;
	    RECT 209.4000 112.8000 209.8000 113.2000 ;
	    RECT 209.4000 112.2000 209.7000 112.8000 ;
	    RECT 210.2000 112.2000 210.5000 113.8000 ;
	    RECT 209.4000 111.8000 209.8000 112.2000 ;
	    RECT 210.2000 111.8000 210.6000 112.2000 ;
	    RECT 207.8000 108.8000 208.2000 109.2000 ;
	    RECT 208.6000 108.8000 209.0000 109.2000 ;
	    RECT 208.6000 108.2000 208.9000 108.8000 ;
	    RECT 208.6000 107.8000 209.0000 108.2000 ;
	    RECT 207.0000 106.8000 207.4000 107.2000 ;
	    RECT 206.2000 105.8000 206.6000 106.2000 ;
	    RECT 204.6000 104.8000 205.0000 105.2000 ;
	    RECT 199.8000 99.1000 200.2000 99.2000 ;
	    RECT 200.6000 99.1000 201.0000 99.2000 ;
	    RECT 199.8000 98.8000 201.0000 99.1000 ;
	    RECT 203.8000 98.8000 204.2000 99.2000 ;
	    RECT 195.0000 94.8000 195.4000 95.2000 ;
	    RECT 196.6000 94.8000 197.0000 95.2000 ;
	    RECT 195.0000 92.2000 195.3000 94.8000 ;
	    RECT 195.0000 91.8000 195.4000 92.2000 ;
	    RECT 196.6000 91.2000 196.9000 94.8000 ;
	    RECT 197.4000 92.1000 197.8000 97.9000 ;
	    RECT 203.8000 96.2000 204.1000 98.8000 ;
	    RECT 204.6000 96.2000 204.9000 104.8000 ;
	    RECT 206.2000 97.2000 206.5000 105.8000 ;
	    RECT 207.0000 104.2000 207.3000 106.8000 ;
	    RECT 207.8000 105.1000 208.2000 105.2000 ;
	    RECT 208.6000 105.1000 208.9000 107.8000 ;
	    RECT 214.2000 107.2000 214.5000 115.8000 ;
	    RECT 218.2000 115.2000 218.5000 115.8000 ;
	    RECT 218.2000 114.8000 218.6000 115.2000 ;
	    RECT 221.4000 114.8000 221.8000 115.2000 ;
	    RECT 223.8000 114.8000 224.2000 115.2000 ;
	    RECT 224.6000 114.8000 225.0000 115.2000 ;
	    RECT 225.4000 114.8000 225.8000 115.2000 ;
	    RECT 221.4000 114.2000 221.7000 114.8000 ;
	    RECT 215.8000 113.8000 216.2000 114.2000 ;
	    RECT 221.4000 113.8000 221.8000 114.2000 ;
	    RECT 223.0000 113.8000 223.4000 114.2000 ;
	    RECT 215.8000 113.2000 216.1000 113.8000 ;
	    RECT 215.8000 112.8000 216.2000 113.2000 ;
	    RECT 218.2000 113.1000 218.6000 113.2000 ;
	    RECT 219.0000 113.1000 219.4000 113.2000 ;
	    RECT 218.2000 112.8000 219.4000 113.1000 ;
	    RECT 220.6000 113.1000 221.0000 113.2000 ;
	    RECT 221.4000 113.1000 221.8000 113.2000 ;
	    RECT 220.6000 112.8000 221.8000 113.1000 ;
	    RECT 222.2000 110.8000 222.6000 111.2000 ;
	    RECT 221.4000 108.8000 221.8000 109.2000 ;
	    RECT 221.4000 108.2000 221.7000 108.8000 ;
	    RECT 222.2000 108.2000 222.5000 110.8000 ;
	    RECT 223.0000 109.2000 223.3000 113.8000 ;
	    RECT 223.8000 109.2000 224.1000 114.8000 ;
	    RECT 224.6000 114.2000 224.9000 114.8000 ;
	    RECT 225.4000 114.2000 225.7000 114.8000 ;
	    RECT 224.6000 113.8000 225.0000 114.2000 ;
	    RECT 225.4000 113.8000 225.8000 114.2000 ;
	    RECT 226.2000 114.0000 226.6000 114.4000 ;
	    RECT 228.6000 114.2000 228.9000 126.8000 ;
	    RECT 229.4000 118.2000 229.7000 145.8000 ;
	    RECT 234.2000 145.2000 234.5000 154.8000 ;
	    RECT 235.0000 154.2000 235.3000 157.8000 ;
	    RECT 235.8000 155.9000 236.2000 156.3000 ;
	    RECT 235.8000 154.2000 236.1000 155.9000 ;
	    RECT 236.6000 155.8000 237.0000 156.2000 ;
	    RECT 239.1000 155.9000 239.5000 156.3000 ;
	    RECT 240.6000 156.1000 240.9000 166.8000 ;
	    RECT 247.0000 166.2000 247.3000 166.8000 ;
	    RECT 249.4000 166.8000 249.8000 167.2000 ;
	    RECT 251.8000 167.1000 252.1000 171.8000 ;
	    RECT 252.6000 171.2000 252.9000 174.8000 ;
	    RECT 254.2000 173.2000 254.5000 175.8000 ;
	    RECT 255.0000 174.8000 255.4000 175.2000 ;
	    RECT 255.0000 174.2000 255.3000 174.8000 ;
	    RECT 255.0000 173.8000 255.4000 174.2000 ;
	    RECT 254.2000 172.8000 254.6000 173.2000 ;
	    RECT 256.6000 173.1000 257.0000 175.9000 ;
	    RECT 257.4000 173.8000 257.8000 174.2000 ;
	    RECT 255.8000 171.8000 256.2000 172.2000 ;
	    RECT 252.6000 170.8000 253.0000 171.2000 ;
	    RECT 255.8000 169.2000 256.1000 171.8000 ;
	    RECT 253.4000 168.8000 253.8000 169.2000 ;
	    RECT 255.8000 168.8000 256.2000 169.2000 ;
	    RECT 252.6000 167.1000 253.0000 167.2000 ;
	    RECT 251.8000 166.8000 253.0000 167.1000 ;
	    RECT 249.4000 166.2000 249.7000 166.8000 ;
	    RECT 253.4000 166.2000 253.7000 168.8000 ;
	    RECT 257.4000 168.2000 257.7000 173.8000 ;
	    RECT 258.2000 172.1000 258.6000 177.9000 ;
	    RECT 259.0000 174.7000 259.4000 175.1000 ;
	    RECT 259.0000 174.2000 259.3000 174.7000 ;
	    RECT 259.0000 173.8000 259.4000 174.2000 ;
	    RECT 260.6000 171.8000 261.0000 172.2000 ;
	    RECT 263.0000 172.1000 263.4000 177.9000 ;
	    RECT 266.2000 176.1000 266.6000 176.2000 ;
	    RECT 267.0000 176.1000 267.4000 176.2000 ;
	    RECT 266.2000 175.8000 267.4000 176.1000 ;
	    RECT 267.0000 174.8000 267.4000 175.2000 ;
	    RECT 267.0000 173.2000 267.3000 174.8000 ;
	    RECT 265.4000 172.8000 265.8000 173.2000 ;
	    RECT 267.0000 172.8000 267.4000 173.2000 ;
	    RECT 265.4000 172.2000 265.7000 172.8000 ;
	    RECT 265.4000 171.8000 265.8000 172.2000 ;
	    RECT 255.8000 167.8000 256.2000 168.2000 ;
	    RECT 257.4000 167.8000 257.8000 168.2000 ;
	    RECT 259.0000 167.8000 259.4000 168.2000 ;
	    RECT 241.4000 165.8000 241.8000 166.2000 ;
	    RECT 244.6000 166.1000 245.0000 166.2000 ;
	    RECT 245.4000 166.1000 245.8000 166.2000 ;
	    RECT 244.6000 165.8000 245.8000 166.1000 ;
	    RECT 246.2000 165.8000 246.6000 166.2000 ;
	    RECT 247.0000 165.8000 247.4000 166.2000 ;
	    RECT 247.8000 166.1000 248.2000 166.2000 ;
	    RECT 248.6000 166.1000 249.0000 166.2000 ;
	    RECT 247.8000 165.8000 249.0000 166.1000 ;
	    RECT 249.4000 165.8000 249.8000 166.2000 ;
	    RECT 251.8000 165.8000 252.2000 166.2000 ;
	    RECT 253.4000 165.8000 253.8000 166.2000 ;
	    RECT 254.2000 165.8000 254.6000 166.2000 ;
	    RECT 241.4000 165.2000 241.7000 165.8000 ;
	    RECT 241.4000 164.8000 241.8000 165.2000 ;
	    RECT 241.4000 163.8000 241.8000 164.2000 ;
	    RECT 241.4000 159.2000 241.7000 163.8000 ;
	    RECT 246.2000 162.2000 246.5000 165.8000 ;
	    RECT 248.6000 165.1000 249.0000 165.2000 ;
	    RECT 247.8000 164.8000 249.0000 165.1000 ;
	    RECT 243.8000 161.8000 244.2000 162.2000 ;
	    RECT 246.2000 161.8000 246.6000 162.2000 ;
	    RECT 243.8000 159.2000 244.1000 161.8000 ;
	    RECT 247.8000 159.2000 248.1000 164.8000 ;
	    RECT 251.8000 161.2000 252.1000 165.8000 ;
	    RECT 251.8000 160.8000 252.2000 161.2000 ;
	    RECT 241.4000 158.8000 241.8000 159.2000 ;
	    RECT 243.8000 158.8000 244.2000 159.2000 ;
	    RECT 247.8000 158.8000 248.2000 159.2000 ;
	    RECT 236.6000 155.2000 236.9000 155.8000 ;
	    RECT 236.6000 154.8000 237.0000 155.2000 ;
	    RECT 237.8000 154.2000 238.2000 154.3000 ;
	    RECT 235.0000 153.8000 235.4000 154.2000 ;
	    RECT 235.8000 153.9000 238.2000 154.2000 ;
	    RECT 235.8000 153.5000 236.1000 153.9000 ;
	    RECT 236.5000 153.5000 236.9000 153.6000 ;
	    RECT 238.2000 153.5000 238.6000 153.6000 ;
	    RECT 239.2000 153.5000 239.5000 155.9000 ;
	    RECT 239.8000 155.8000 240.9000 156.1000 ;
	    RECT 247.8000 157.8000 248.2000 158.2000 ;
	    RECT 239.8000 154.2000 240.1000 155.8000 ;
	    RECT 240.6000 154.8000 241.0000 155.2000 ;
	    RECT 243.0000 154.8000 243.4000 155.2000 ;
	    RECT 246.2000 154.8000 246.6000 155.2000 ;
	    RECT 239.8000 153.8000 240.2000 154.2000 ;
	    RECT 235.8000 153.1000 236.2000 153.5000 ;
	    RECT 236.5000 153.2000 238.6000 153.5000 ;
	    RECT 239.1000 153.1000 239.5000 153.5000 ;
	    RECT 239.0000 151.1000 239.4000 151.2000 ;
	    RECT 238.2000 150.8000 239.4000 151.1000 ;
	    RECT 235.8000 149.8000 236.2000 150.2000 ;
	    RECT 235.8000 149.2000 236.1000 149.8000 ;
	    RECT 238.2000 149.2000 238.5000 150.8000 ;
	    RECT 239.0000 149.8000 239.4000 150.2000 ;
	    RECT 235.8000 148.8000 236.2000 149.2000 ;
	    RECT 238.2000 148.8000 238.6000 149.2000 ;
	    RECT 239.0000 148.2000 239.3000 149.8000 ;
	    RECT 239.0000 147.8000 239.4000 148.2000 ;
	    RECT 239.8000 147.8000 240.2000 148.2000 ;
	    RECT 239.8000 147.2000 240.1000 147.8000 ;
	    RECT 239.8000 146.8000 240.2000 147.2000 ;
	    RECT 240.6000 146.2000 240.9000 154.8000 ;
	    RECT 243.0000 153.2000 243.3000 154.8000 ;
	    RECT 246.2000 154.2000 246.5000 154.8000 ;
	    RECT 246.2000 153.8000 246.6000 154.2000 ;
	    RECT 247.8000 153.2000 248.1000 157.8000 ;
	    RECT 249.4000 156.8000 249.8000 157.2000 ;
	    RECT 249.4000 156.2000 249.7000 156.8000 ;
	    RECT 254.2000 156.2000 254.5000 165.8000 ;
	    RECT 255.0000 164.8000 255.4000 165.2000 ;
	    RECT 255.0000 164.2000 255.3000 164.8000 ;
	    RECT 255.0000 163.8000 255.4000 164.2000 ;
	    RECT 255.8000 163.1000 256.1000 167.8000 ;
	    RECT 257.4000 166.8000 257.8000 167.2000 ;
	    RECT 257.4000 166.2000 257.7000 166.8000 ;
	    RECT 257.4000 165.8000 257.8000 166.2000 ;
	    RECT 259.0000 164.2000 259.3000 167.8000 ;
	    RECT 260.6000 167.2000 260.9000 171.8000 ;
	    RECT 263.8000 169.8000 264.2000 170.2000 ;
	    RECT 263.8000 169.2000 264.1000 169.8000 ;
	    RECT 263.8000 168.8000 264.2000 169.2000 ;
	    RECT 263.0000 167.5000 263.4000 167.9000 ;
	    RECT 266.1000 167.8000 266.5000 167.9000 ;
	    RECT 263.7000 167.5000 266.5000 167.8000 ;
	    RECT 260.6000 166.8000 261.0000 167.2000 ;
	    RECT 262.2000 166.8000 262.6000 167.2000 ;
	    RECT 263.0000 167.1000 263.3000 167.5000 ;
	    RECT 263.7000 167.4000 264.1000 167.5000 ;
	    RECT 265.4000 167.4000 265.8000 167.5000 ;
	    RECT 263.0000 166.8000 265.8000 167.1000 ;
	    RECT 261.4000 165.8000 261.8000 166.2000 ;
	    RECT 259.0000 163.8000 259.4000 164.2000 ;
	    RECT 255.0000 162.8000 256.1000 163.1000 ;
	    RECT 255.0000 159.2000 255.3000 162.8000 ;
	    RECT 255.8000 161.8000 256.2000 162.2000 ;
	    RECT 255.8000 160.2000 256.1000 161.8000 ;
	    RECT 255.8000 159.8000 256.2000 160.2000 ;
	    RECT 255.0000 158.8000 255.4000 159.2000 ;
	    RECT 259.0000 158.8000 259.4000 159.2000 ;
	    RECT 249.4000 155.8000 249.8000 156.2000 ;
	    RECT 253.4000 155.8000 253.8000 156.2000 ;
	    RECT 254.2000 155.8000 254.6000 156.2000 ;
	    RECT 255.8000 156.1000 256.2000 156.2000 ;
	    RECT 256.6000 156.1000 257.0000 156.2000 ;
	    RECT 255.8000 155.8000 257.0000 156.1000 ;
	    RECT 257.4000 155.8000 257.8000 156.2000 ;
	    RECT 253.4000 155.2000 253.7000 155.8000 ;
	    RECT 257.4000 155.2000 257.7000 155.8000 ;
	    RECT 250.2000 154.8000 250.6000 155.2000 ;
	    RECT 253.4000 154.8000 253.8000 155.2000 ;
	    RECT 254.2000 155.1000 254.6000 155.2000 ;
	    RECT 255.0000 155.1000 255.4000 155.2000 ;
	    RECT 254.2000 154.8000 255.4000 155.1000 ;
	    RECT 257.4000 154.8000 257.8000 155.2000 ;
	    RECT 242.2000 152.8000 242.6000 153.2000 ;
	    RECT 243.0000 152.8000 243.4000 153.2000 ;
	    RECT 244.6000 152.8000 245.0000 153.2000 ;
	    RECT 247.8000 152.8000 248.2000 153.2000 ;
	    RECT 248.6000 152.8000 249.0000 153.2000 ;
	    RECT 242.2000 150.2000 242.5000 152.8000 ;
	    RECT 244.6000 150.2000 244.9000 152.8000 ;
	    RECT 242.2000 149.8000 242.6000 150.2000 ;
	    RECT 244.6000 149.8000 245.0000 150.2000 ;
	    RECT 247.8000 149.2000 248.1000 152.8000 ;
	    RECT 248.6000 149.2000 248.9000 152.8000 ;
	    RECT 250.2000 152.2000 250.5000 154.8000 ;
	    RECT 252.6000 153.8000 253.0000 154.2000 ;
	    RECT 252.6000 153.2000 252.9000 153.8000 ;
	    RECT 251.0000 152.8000 251.4000 153.2000 ;
	    RECT 252.6000 152.8000 253.0000 153.2000 ;
	    RECT 251.0000 152.2000 251.3000 152.8000 ;
	    RECT 250.2000 151.8000 250.6000 152.2000 ;
	    RECT 251.0000 151.8000 251.4000 152.2000 ;
	    RECT 251.8000 151.8000 252.2000 152.2000 ;
	    RECT 251.8000 151.2000 252.1000 151.8000 ;
	    RECT 250.2000 150.8000 250.6000 151.2000 ;
	    RECT 251.8000 150.8000 252.2000 151.2000 ;
	    RECT 249.4000 149.8000 249.8000 150.2000 ;
	    RECT 247.8000 148.8000 248.2000 149.2000 ;
	    RECT 248.6000 148.8000 249.0000 149.2000 ;
	    RECT 243.0000 147.8000 243.4000 148.2000 ;
	    RECT 248.6000 148.1000 249.0000 148.2000 ;
	    RECT 249.4000 148.1000 249.7000 149.8000 ;
	    RECT 248.6000 147.8000 249.7000 148.1000 ;
	    RECT 243.0000 147.2000 243.3000 147.8000 ;
	    RECT 243.0000 146.8000 243.4000 147.2000 ;
	    RECT 244.6000 146.8000 245.0000 147.2000 ;
	    RECT 244.6000 146.2000 244.9000 146.8000 ;
	    RECT 237.4000 145.8000 237.8000 146.2000 ;
	    RECT 239.0000 145.8000 239.4000 146.2000 ;
	    RECT 240.6000 145.8000 241.0000 146.2000 ;
	    RECT 241.4000 145.8000 241.8000 146.2000 ;
	    RECT 242.2000 146.1000 242.6000 146.2000 ;
	    RECT 243.0000 146.1000 243.4000 146.2000 ;
	    RECT 242.2000 145.8000 243.4000 146.1000 ;
	    RECT 244.6000 145.8000 245.0000 146.2000 ;
	    RECT 247.0000 145.8000 247.4000 146.2000 ;
	    RECT 230.2000 144.8000 230.6000 145.2000 ;
	    RECT 234.2000 144.8000 234.6000 145.2000 ;
	    RECT 230.2000 139.2000 230.5000 144.8000 ;
	    RECT 237.4000 144.2000 237.7000 145.8000 ;
	    RECT 237.4000 143.8000 237.8000 144.2000 ;
	    RECT 230.2000 138.8000 230.6000 139.2000 ;
	    RECT 237.4000 138.1000 237.8000 138.2000 ;
	    RECT 238.2000 138.1000 238.6000 138.2000 ;
	    RECT 237.4000 137.8000 238.6000 138.1000 ;
	    RECT 233.4000 136.8000 233.8000 137.2000 ;
	    RECT 234.2000 137.1000 234.6000 137.2000 ;
	    RECT 235.0000 137.1000 235.4000 137.2000 ;
	    RECT 234.2000 136.8000 235.4000 137.1000 ;
	    RECT 233.4000 136.2000 233.7000 136.8000 ;
	    RECT 231.0000 135.8000 231.4000 136.2000 ;
	    RECT 231.8000 136.1000 232.2000 136.2000 ;
	    RECT 232.6000 136.1000 233.0000 136.2000 ;
	    RECT 231.8000 135.8000 233.0000 136.1000 ;
	    RECT 233.4000 135.8000 233.8000 136.2000 ;
	    RECT 235.8000 135.8000 236.2000 136.2000 ;
	    RECT 231.0000 133.2000 231.3000 135.8000 ;
	    RECT 233.4000 134.2000 233.7000 135.8000 ;
	    RECT 235.8000 135.2000 236.1000 135.8000 ;
	    RECT 235.8000 134.8000 236.2000 135.2000 ;
	    RECT 238.2000 135.1000 238.6000 135.2000 ;
	    RECT 239.0000 135.1000 239.3000 145.8000 ;
	    RECT 239.8000 145.1000 240.2000 145.2000 ;
	    RECT 240.6000 145.1000 241.0000 145.2000 ;
	    RECT 239.8000 144.8000 241.0000 145.1000 ;
	    RECT 241.4000 139.2000 241.7000 145.8000 ;
	    RECT 243.0000 145.1000 243.4000 145.2000 ;
	    RECT 243.8000 145.1000 244.2000 145.2000 ;
	    RECT 243.0000 144.8000 244.2000 145.1000 ;
	    RECT 245.4000 144.1000 245.8000 144.2000 ;
	    RECT 246.2000 144.1000 246.6000 144.2000 ;
	    RECT 245.4000 143.8000 246.6000 144.1000 ;
	    RECT 244.6000 142.8000 245.0000 143.2000 ;
	    RECT 244.6000 142.2000 244.9000 142.8000 ;
	    RECT 244.6000 141.8000 245.0000 142.2000 ;
	    RECT 242.2000 140.8000 242.6000 141.2000 ;
	    RECT 242.2000 139.2000 242.5000 140.8000 ;
	    RECT 241.4000 138.8000 241.8000 139.2000 ;
	    RECT 242.2000 138.8000 242.6000 139.2000 ;
	    RECT 241.4000 136.8000 241.8000 137.2000 ;
	    RECT 238.2000 134.8000 239.3000 135.1000 ;
	    RECT 240.6000 135.8000 241.0000 136.2000 ;
	    RECT 240.6000 135.2000 240.9000 135.8000 ;
	    RECT 241.4000 135.2000 241.7000 136.8000 ;
	    RECT 240.6000 134.8000 241.0000 135.2000 ;
	    RECT 241.4000 134.8000 241.8000 135.2000 ;
	    RECT 231.8000 134.1000 232.2000 134.2000 ;
	    RECT 232.6000 134.1000 233.0000 134.2000 ;
	    RECT 231.8000 133.8000 233.0000 134.1000 ;
	    RECT 233.4000 133.8000 233.8000 134.2000 ;
	    RECT 231.0000 132.8000 231.4000 133.2000 ;
	    RECT 236.6000 133.1000 237.0000 133.2000 ;
	    RECT 237.4000 133.1000 237.8000 133.2000 ;
	    RECT 236.6000 132.8000 237.8000 133.1000 ;
	    RECT 230.2000 131.8000 230.6000 132.2000 ;
	    RECT 230.2000 127.2000 230.5000 131.8000 ;
	    RECT 230.2000 126.8000 230.6000 127.2000 ;
	    RECT 229.4000 117.8000 229.8000 118.2000 ;
	    RECT 231.0000 116.2000 231.3000 132.8000 ;
	    RECT 238.2000 132.2000 238.5000 134.8000 ;
	    RECT 239.0000 132.8000 239.4000 133.2000 ;
	    RECT 238.2000 131.8000 238.6000 132.2000 ;
	    RECT 231.8000 129.8000 232.2000 130.2000 ;
	    RECT 231.8000 129.2000 232.1000 129.8000 ;
	    RECT 231.8000 128.8000 232.2000 129.2000 ;
	    RECT 232.6000 128.8000 233.0000 129.2000 ;
	    RECT 235.0000 128.8000 235.4000 129.2000 ;
	    RECT 232.6000 127.2000 232.9000 128.8000 ;
	    RECT 235.0000 128.2000 235.3000 128.8000 ;
	    RECT 235.0000 127.8000 235.4000 128.2000 ;
	    RECT 235.8000 127.8000 236.2000 128.2000 ;
	    RECT 232.6000 126.8000 233.0000 127.2000 ;
	    RECT 233.4000 126.8000 233.8000 127.2000 ;
	    RECT 233.4000 126.2000 233.7000 126.8000 ;
	    RECT 233.4000 125.8000 233.8000 126.2000 ;
	    RECT 234.2000 121.8000 234.6000 122.2000 ;
	    RECT 234.2000 121.2000 234.5000 121.8000 ;
	    RECT 234.2000 120.8000 234.6000 121.2000 ;
	    RECT 235.0000 117.2000 235.3000 127.8000 ;
	    RECT 235.8000 124.2000 236.1000 127.8000 ;
	    RECT 236.6000 126.1000 237.0000 126.2000 ;
	    RECT 237.4000 126.1000 237.8000 126.2000 ;
	    RECT 236.6000 125.8000 237.8000 126.1000 ;
	    RECT 238.2000 124.8000 238.6000 125.2000 ;
	    RECT 238.2000 124.2000 238.5000 124.8000 ;
	    RECT 235.8000 123.8000 236.2000 124.2000 ;
	    RECT 238.2000 123.8000 238.6000 124.2000 ;
	    RECT 239.0000 123.2000 239.3000 132.8000 ;
	    RECT 239.8000 131.8000 240.2000 132.2000 ;
	    RECT 239.8000 131.2000 240.1000 131.8000 ;
	    RECT 239.8000 130.8000 240.2000 131.2000 ;
	    RECT 239.8000 126.1000 240.2000 126.2000 ;
	    RECT 240.6000 126.1000 241.0000 126.2000 ;
	    RECT 239.8000 125.8000 241.0000 126.1000 ;
	    RECT 240.6000 123.8000 241.0000 124.2000 ;
	    RECT 240.6000 123.2000 240.9000 123.8000 ;
	    RECT 238.2000 122.8000 238.6000 123.2000 ;
	    RECT 239.0000 122.8000 239.4000 123.2000 ;
	    RECT 240.6000 122.8000 241.0000 123.2000 ;
	    RECT 235.0000 116.8000 235.4000 117.2000 ;
	    RECT 229.4000 116.1000 229.8000 116.2000 ;
	    RECT 230.2000 116.1000 230.6000 116.2000 ;
	    RECT 229.4000 115.8000 230.6000 116.1000 ;
	    RECT 231.0000 115.8000 231.4000 116.2000 ;
	    RECT 236.6000 116.1000 237.0000 116.2000 ;
	    RECT 237.4000 116.1000 237.8000 116.2000 ;
	    RECT 236.6000 115.8000 237.8000 116.1000 ;
	    RECT 230.2000 115.2000 230.5000 115.8000 ;
	    RECT 230.2000 114.8000 230.6000 115.2000 ;
	    RECT 231.0000 114.8000 231.4000 115.2000 ;
	    RECT 235.0000 114.8000 235.4000 115.2000 ;
	    RECT 235.8000 114.8000 236.2000 115.2000 ;
	    RECT 231.0000 114.2000 231.3000 114.8000 ;
	    RECT 235.0000 114.2000 235.3000 114.8000 ;
	    RECT 235.8000 114.2000 236.1000 114.8000 ;
	    RECT 237.4000 114.2000 237.7000 115.8000 ;
	    RECT 226.2000 113.2000 226.5000 114.0000 ;
	    RECT 228.6000 113.8000 229.0000 114.2000 ;
	    RECT 231.0000 113.8000 231.4000 114.2000 ;
	    RECT 235.0000 113.8000 235.4000 114.2000 ;
	    RECT 235.8000 113.8000 236.2000 114.2000 ;
	    RECT 237.4000 113.8000 237.8000 114.2000 ;
	    RECT 226.2000 112.8000 226.6000 113.2000 ;
	    RECT 232.6000 112.8000 233.0000 113.2000 ;
	    RECT 227.8000 111.8000 228.2000 112.2000 ;
	    RECT 231.8000 111.8000 232.2000 112.2000 ;
	    RECT 223.0000 108.8000 223.4000 109.2000 ;
	    RECT 223.8000 108.8000 224.2000 109.2000 ;
	    RECT 215.8000 107.8000 216.2000 108.2000 ;
	    RECT 216.6000 107.8000 217.0000 108.2000 ;
	    RECT 218.2000 107.8000 218.6000 108.2000 ;
	    RECT 221.4000 107.8000 221.8000 108.2000 ;
	    RECT 222.2000 107.8000 222.6000 108.2000 ;
	    RECT 215.8000 107.2000 216.1000 107.8000 ;
	    RECT 209.4000 107.1000 209.8000 107.2000 ;
	    RECT 210.2000 107.1000 210.6000 107.2000 ;
	    RECT 209.4000 106.8000 210.6000 107.1000 ;
	    RECT 214.2000 106.8000 214.6000 107.2000 ;
	    RECT 215.8000 106.8000 216.2000 107.2000 ;
	    RECT 216.6000 106.2000 216.9000 107.8000 ;
	    RECT 218.2000 107.2000 218.5000 107.8000 ;
	    RECT 218.2000 106.8000 218.6000 107.2000 ;
	    RECT 224.6000 107.1000 225.0000 107.2000 ;
	    RECT 225.4000 107.1000 225.8000 107.2000 ;
	    RECT 224.6000 106.8000 225.8000 107.1000 ;
	    RECT 226.2000 106.8000 226.6000 107.2000 ;
	    RECT 227.0000 106.8000 227.4000 107.2000 ;
	    RECT 207.8000 104.8000 208.9000 105.1000 ;
	    RECT 209.4000 105.8000 209.8000 106.2000 ;
	    RECT 211.0000 106.1000 211.4000 106.2000 ;
	    RECT 211.8000 106.1000 212.2000 106.2000 ;
	    RECT 211.0000 105.8000 212.2000 106.1000 ;
	    RECT 215.0000 106.1000 215.4000 106.2000 ;
	    RECT 215.8000 106.1000 216.2000 106.2000 ;
	    RECT 215.0000 105.8000 216.2000 106.1000 ;
	    RECT 216.6000 105.8000 217.0000 106.2000 ;
	    RECT 217.4000 105.8000 217.8000 106.2000 ;
	    RECT 219.8000 106.1000 220.2000 106.2000 ;
	    RECT 220.6000 106.1000 221.0000 106.2000 ;
	    RECT 219.8000 105.8000 221.0000 106.1000 ;
	    RECT 222.2000 105.8000 222.6000 106.2000 ;
	    RECT 225.4000 106.1000 225.8000 106.2000 ;
	    RECT 226.2000 106.1000 226.5000 106.8000 ;
	    RECT 225.4000 105.8000 226.5000 106.1000 ;
	    RECT 227.0000 106.2000 227.3000 106.8000 ;
	    RECT 227.0000 105.8000 227.4000 106.2000 ;
	    RECT 209.4000 105.1000 209.7000 105.8000 ;
	    RECT 217.4000 105.2000 217.7000 105.8000 ;
	    RECT 211.8000 105.1000 212.2000 105.2000 ;
	    RECT 209.4000 104.8000 212.2000 105.1000 ;
	    RECT 217.4000 104.8000 217.8000 105.2000 ;
	    RECT 207.0000 103.8000 207.4000 104.2000 ;
	    RECT 222.2000 99.2000 222.5000 105.8000 ;
	    RECT 223.0000 104.8000 223.4000 105.2000 ;
	    RECT 223.0000 104.2000 223.3000 104.8000 ;
	    RECT 223.0000 103.8000 223.4000 104.2000 ;
	    RECT 225.4000 99.2000 225.7000 105.8000 ;
	    RECT 222.2000 98.8000 222.6000 99.2000 ;
	    RECT 225.4000 98.8000 225.8000 99.2000 ;
	    RECT 223.8000 97.8000 224.2000 98.2000 ;
	    RECT 205.4000 96.8000 205.8000 97.2000 ;
	    RECT 206.2000 96.8000 206.6000 97.2000 ;
	    RECT 211.0000 96.8000 211.4000 97.2000 ;
	    RECT 203.8000 95.8000 204.2000 96.2000 ;
	    RECT 204.6000 95.8000 205.0000 96.2000 ;
	    RECT 205.4000 95.2000 205.7000 96.8000 ;
	    RECT 208.6000 96.1000 209.0000 96.2000 ;
	    RECT 209.4000 96.1000 209.8000 96.2000 ;
	    RECT 208.6000 95.8000 209.8000 96.1000 ;
	    RECT 205.4000 94.8000 205.8000 95.2000 ;
	    RECT 207.0000 94.8000 207.4000 95.2000 ;
	    RECT 209.4000 94.8000 209.8000 95.2000 ;
	    RECT 200.6000 93.8000 201.0000 94.2000 ;
	    RECT 202.2000 93.8000 202.6000 94.2000 ;
	    RECT 200.6000 93.2000 200.9000 93.8000 ;
	    RECT 202.2000 93.2000 202.5000 93.8000 ;
	    RECT 200.6000 92.8000 201.0000 93.2000 ;
	    RECT 201.4000 92.8000 201.8000 93.2000 ;
	    RECT 202.2000 92.8000 202.6000 93.2000 ;
	    RECT 201.4000 92.2000 201.7000 92.8000 ;
	    RECT 201.4000 91.8000 201.8000 92.2000 ;
	    RECT 196.6000 90.8000 197.0000 91.2000 ;
	    RECT 200.6000 89.8000 201.0000 90.2000 ;
	    RECT 198.2000 88.8000 198.6000 89.2000 ;
	    RECT 198.2000 88.2000 198.5000 88.8000 ;
	    RECT 200.6000 88.2000 200.9000 89.8000 ;
	    RECT 197.4000 87.8000 197.8000 88.2000 ;
	    RECT 198.2000 87.8000 198.6000 88.2000 ;
	    RECT 199.0000 87.8000 199.4000 88.2000 ;
	    RECT 200.6000 87.8000 201.0000 88.2000 ;
	    RECT 197.4000 87.2000 197.7000 87.8000 ;
	    RECT 184.6000 86.8000 185.0000 87.2000 ;
	    RECT 185.4000 86.8000 185.8000 87.2000 ;
	    RECT 187.8000 86.8000 188.2000 87.2000 ;
	    RECT 190.2000 86.8000 190.6000 87.2000 ;
	    RECT 191.8000 86.8000 192.2000 87.2000 ;
	    RECT 194.2000 86.8000 194.6000 87.2000 ;
	    RECT 197.4000 86.8000 197.8000 87.2000 ;
	    RECT 181.4000 85.8000 181.8000 86.2000 ;
	    RECT 184.6000 85.2000 184.9000 86.8000 ;
	    RECT 185.4000 86.2000 185.7000 86.8000 ;
	    RECT 191.8000 86.2000 192.1000 86.8000 ;
	    RECT 199.0000 86.2000 199.3000 87.8000 ;
	    RECT 200.6000 86.2000 200.9000 87.8000 ;
	    RECT 201.4000 87.1000 201.8000 87.2000 ;
	    RECT 202.2000 87.1000 202.6000 87.2000 ;
	    RECT 201.4000 86.8000 202.6000 87.1000 ;
	    RECT 185.4000 85.8000 185.8000 86.2000 ;
	    RECT 191.8000 85.8000 192.2000 86.2000 ;
	    RECT 195.0000 86.1000 195.4000 86.2000 ;
	    RECT 195.8000 86.1000 196.2000 86.2000 ;
	    RECT 195.0000 85.8000 196.2000 86.1000 ;
	    RECT 199.0000 85.8000 199.4000 86.2000 ;
	    RECT 200.6000 85.8000 201.0000 86.2000 ;
	    RECT 179.8000 84.8000 180.2000 85.2000 ;
	    RECT 184.6000 84.8000 185.0000 85.2000 ;
	    RECT 195.8000 85.1000 196.2000 85.2000 ;
	    RECT 196.6000 85.1000 197.0000 85.2000 ;
	    RECT 195.8000 84.8000 197.0000 85.1000 ;
	    RECT 179.8000 80.2000 180.1000 84.8000 ;
	    RECT 181.4000 81.8000 181.8000 82.2000 ;
	    RECT 179.8000 79.8000 180.2000 80.2000 ;
	    RECT 171.0000 74.8000 171.4000 75.2000 ;
	    RECT 173.4000 74.8000 173.8000 75.2000 ;
	    RECT 171.0000 73.2000 171.3000 74.8000 ;
	    RECT 173.4000 73.8000 173.8000 74.2000 ;
	    RECT 171.0000 72.8000 171.4000 73.2000 ;
	    RECT 173.4000 68.2000 173.7000 73.8000 ;
	    RECT 174.2000 72.1000 174.6000 77.9000 ;
	    RECT 177.4000 75.8000 177.8000 76.2000 ;
	    RECT 177.4000 72.2000 177.7000 75.8000 ;
	    RECT 179.8000 74.2000 180.1000 79.8000 ;
	    RECT 181.4000 77.2000 181.7000 81.8000 ;
	    RECT 181.4000 76.8000 181.8000 77.2000 ;
	    RECT 183.0000 77.1000 183.4000 77.2000 ;
	    RECT 183.8000 77.1000 184.2000 77.2000 ;
	    RECT 183.0000 76.8000 184.2000 77.1000 ;
	    RECT 184.6000 75.2000 184.9000 84.8000 ;
	    RECT 199.0000 84.2000 199.3000 85.8000 ;
	    RECT 199.8000 84.8000 200.2000 85.2000 ;
	    RECT 199.8000 84.2000 200.1000 84.8000 ;
	    RECT 194.2000 84.1000 194.6000 84.2000 ;
	    RECT 195.0000 84.1000 195.4000 84.2000 ;
	    RECT 194.2000 83.8000 195.4000 84.1000 ;
	    RECT 195.8000 83.8000 196.2000 84.2000 ;
	    RECT 199.0000 83.8000 199.4000 84.2000 ;
	    RECT 199.8000 83.8000 200.2000 84.2000 ;
	    RECT 195.0000 82.2000 195.3000 83.8000 ;
	    RECT 195.8000 83.2000 196.1000 83.8000 ;
	    RECT 195.8000 82.8000 196.2000 83.2000 ;
	    RECT 195.0000 81.8000 195.4000 82.2000 ;
	    RECT 188.6000 80.8000 189.0000 81.2000 ;
	    RECT 199.0000 80.8000 199.4000 81.2000 ;
	    RECT 185.4000 76.8000 185.8000 77.2000 ;
	    RECT 185.4000 76.2000 185.7000 76.8000 ;
	    RECT 188.6000 76.2000 188.9000 80.8000 ;
	    RECT 191.0000 76.8000 191.4000 77.2000 ;
	    RECT 194.2000 76.8000 194.6000 77.2000 ;
	    RECT 185.4000 75.8000 185.8000 76.2000 ;
	    RECT 188.6000 75.8000 189.0000 76.2000 ;
	    RECT 181.4000 74.8000 181.8000 75.2000 ;
	    RECT 182.2000 74.8000 182.6000 75.2000 ;
	    RECT 184.6000 74.8000 185.0000 75.2000 ;
	    RECT 186.2000 74.8000 186.6000 75.2000 ;
	    RECT 181.4000 74.2000 181.7000 74.8000 ;
	    RECT 178.2000 73.8000 178.6000 74.2000 ;
	    RECT 179.8000 73.8000 180.2000 74.2000 ;
	    RECT 181.4000 73.8000 181.8000 74.2000 ;
	    RECT 178.2000 73.2000 178.5000 73.8000 ;
	    RECT 178.2000 72.8000 178.6000 73.2000 ;
	    RECT 179.0000 73.1000 179.4000 73.2000 ;
	    RECT 179.8000 73.1000 180.2000 73.2000 ;
	    RECT 179.0000 72.8000 180.2000 73.1000 ;
	    RECT 175.0000 71.8000 175.4000 72.2000 ;
	    RECT 175.8000 72.1000 176.2000 72.2000 ;
	    RECT 176.6000 72.1000 177.0000 72.2000 ;
	    RECT 175.8000 71.8000 177.0000 72.1000 ;
	    RECT 177.4000 71.8000 177.8000 72.2000 ;
	    RECT 180.6000 71.8000 181.0000 72.2000 ;
	    RECT 175.0000 68.2000 175.3000 71.8000 ;
	    RECT 173.4000 68.1000 173.8000 68.2000 ;
	    RECT 174.2000 68.1000 174.6000 68.2000 ;
	    RECT 173.4000 67.8000 174.6000 68.1000 ;
	    RECT 175.0000 67.8000 175.4000 68.2000 ;
	    RECT 176.6000 67.8000 177.0000 68.2000 ;
	    RECT 176.6000 67.2000 176.9000 67.8000 ;
	    RECT 175.0000 67.1000 175.4000 67.2000 ;
	    RECT 175.8000 67.1000 176.2000 67.2000 ;
	    RECT 175.0000 66.8000 176.2000 67.1000 ;
	    RECT 176.6000 66.8000 177.0000 67.2000 ;
	    RECT 172.6000 65.8000 173.0000 66.2000 ;
	    RECT 167.8000 61.8000 168.2000 62.2000 ;
	    RECT 171.8000 61.8000 172.2000 62.2000 ;
	    RECT 167.8000 59.2000 168.1000 61.8000 ;
	    RECT 167.8000 58.8000 168.2000 59.2000 ;
	    RECT 167.0000 54.8000 167.4000 55.2000 ;
	    RECT 166.2000 53.8000 166.6000 54.2000 ;
	    RECT 166.2000 49.2000 166.5000 53.8000 ;
	    RECT 167.8000 52.1000 168.2000 57.9000 ;
	    RECT 170.2000 54.1000 170.6000 54.2000 ;
	    RECT 171.0000 54.1000 171.4000 54.2000 ;
	    RECT 170.2000 53.8000 171.4000 54.1000 ;
	    RECT 170.2000 51.8000 170.6000 52.2000 ;
	    RECT 170.2000 51.2000 170.5000 51.8000 ;
	    RECT 170.2000 50.8000 170.6000 51.2000 ;
	    RECT 166.2000 48.8000 166.6000 49.2000 ;
	    RECT 165.4000 47.8000 165.8000 48.2000 ;
	    RECT 168.6000 43.1000 169.0000 48.9000 ;
	    RECT 171.8000 48.2000 172.1000 61.8000 ;
	    RECT 172.6000 56.2000 172.9000 65.8000 ;
	    RECT 176.6000 65.1000 177.0000 65.2000 ;
	    RECT 177.4000 65.1000 177.7000 71.8000 ;
	    RECT 178.2000 67.1000 178.6000 67.2000 ;
	    RECT 179.0000 67.1000 179.4000 67.2000 ;
	    RECT 178.2000 66.8000 179.4000 67.1000 ;
	    RECT 180.6000 67.1000 180.9000 71.8000 ;
	    RECT 182.2000 71.2000 182.5000 74.8000 ;
	    RECT 186.2000 74.2000 186.5000 74.8000 ;
	    RECT 184.6000 73.8000 185.0000 74.2000 ;
	    RECT 186.2000 73.8000 186.6000 74.2000 ;
	    RECT 189.4000 74.1000 189.8000 74.2000 ;
	    RECT 190.2000 74.1000 190.6000 74.2000 ;
	    RECT 189.4000 73.8000 190.6000 74.1000 ;
	    RECT 184.6000 73.2000 184.9000 73.8000 ;
	    RECT 184.6000 72.8000 185.0000 73.2000 ;
	    RECT 182.2000 70.8000 182.6000 71.2000 ;
	    RECT 186.2000 68.2000 186.5000 73.8000 ;
	    RECT 191.0000 73.2000 191.3000 76.8000 ;
	    RECT 194.2000 76.2000 194.5000 76.8000 ;
	    RECT 194.2000 75.8000 194.6000 76.2000 ;
	    RECT 191.8000 74.8000 192.2000 75.2000 ;
	    RECT 193.4000 74.8000 193.8000 75.2000 ;
	    RECT 195.8000 74.8000 196.2000 75.2000 ;
	    RECT 191.8000 74.2000 192.1000 74.8000 ;
	    RECT 193.4000 74.2000 193.7000 74.8000 ;
	    RECT 195.8000 74.2000 196.1000 74.8000 ;
	    RECT 199.0000 74.2000 199.3000 80.8000 ;
	    RECT 201.4000 78.1000 201.7000 86.8000 ;
	    RECT 200.6000 77.8000 201.7000 78.1000 ;
	    RECT 202.2000 85.8000 202.6000 86.2000 ;
	    RECT 203.0000 85.8000 203.4000 86.2000 ;
	    RECT 200.6000 75.2000 200.9000 77.8000 ;
	    RECT 201.4000 76.8000 201.8000 77.2000 ;
	    RECT 201.4000 76.2000 201.7000 76.8000 ;
	    RECT 201.4000 75.8000 201.8000 76.2000 ;
	    RECT 199.8000 74.8000 200.2000 75.2000 ;
	    RECT 200.6000 74.8000 201.0000 75.2000 ;
	    RECT 191.8000 73.8000 192.2000 74.2000 ;
	    RECT 193.4000 73.8000 193.8000 74.2000 ;
	    RECT 195.8000 73.8000 196.2000 74.2000 ;
	    RECT 199.0000 73.8000 199.4000 74.2000 ;
	    RECT 187.0000 72.8000 187.4000 73.2000 ;
	    RECT 187.8000 72.8000 188.2000 73.2000 ;
	    RECT 191.0000 72.8000 191.4000 73.2000 ;
	    RECT 187.0000 72.2000 187.3000 72.8000 ;
	    RECT 187.0000 71.8000 187.4000 72.2000 ;
	    RECT 183.8000 67.8000 184.2000 68.2000 ;
	    RECT 186.2000 67.8000 186.6000 68.2000 ;
	    RECT 183.8000 67.2000 184.1000 67.8000 ;
	    RECT 180.6000 66.8000 181.7000 67.1000 ;
	    RECT 183.8000 66.8000 184.2000 67.2000 ;
	    RECT 185.4000 67.1000 185.8000 67.2000 ;
	    RECT 186.2000 67.1000 186.6000 67.2000 ;
	    RECT 185.4000 66.8000 186.6000 67.1000 ;
	    RECT 187.0000 67.1000 187.4000 67.2000 ;
	    RECT 187.8000 67.1000 188.1000 72.8000 ;
	    RECT 191.0000 70.2000 191.3000 72.8000 ;
	    RECT 191.0000 69.8000 191.4000 70.2000 ;
	    RECT 191.8000 67.2000 192.1000 73.8000 ;
	    RECT 199.8000 73.2000 200.1000 74.8000 ;
	    RECT 202.2000 74.2000 202.5000 85.8000 ;
	    RECT 203.0000 76.2000 203.3000 85.8000 ;
	    RECT 205.4000 85.2000 205.7000 94.8000 ;
	    RECT 207.0000 94.2000 207.3000 94.8000 ;
	    RECT 209.4000 94.2000 209.7000 94.8000 ;
	    RECT 206.2000 93.8000 206.6000 94.2000 ;
	    RECT 207.0000 93.8000 207.4000 94.2000 ;
	    RECT 209.4000 93.8000 209.8000 94.2000 ;
	    RECT 206.2000 88.2000 206.5000 93.8000 ;
	    RECT 207.0000 88.2000 207.3000 93.8000 ;
	    RECT 211.0000 93.2000 211.3000 96.8000 ;
	    RECT 216.7000 95.9000 217.1000 96.3000 ;
	    RECT 219.8000 95.9000 220.2000 96.3000 ;
	    RECT 215.8000 94.8000 216.2000 95.2000 ;
	    RECT 215.8000 94.2000 216.1000 94.8000 ;
	    RECT 215.0000 93.8000 215.4000 94.2000 ;
	    RECT 215.8000 93.8000 216.2000 94.2000 ;
	    RECT 211.0000 92.8000 211.4000 93.2000 ;
	    RECT 212.6000 93.1000 213.0000 93.2000 ;
	    RECT 213.4000 93.1000 213.8000 93.2000 ;
	    RECT 212.6000 92.8000 213.8000 93.1000 ;
	    RECT 215.0000 92.2000 215.3000 93.8000 ;
	    RECT 208.6000 91.8000 209.0000 92.2000 ;
	    RECT 215.0000 91.8000 215.4000 92.2000 ;
	    RECT 208.6000 88.2000 208.9000 91.8000 ;
	    RECT 215.0000 89.8000 215.4000 90.2000 ;
	    RECT 206.2000 87.8000 206.6000 88.2000 ;
	    RECT 207.0000 87.8000 207.4000 88.2000 ;
	    RECT 208.6000 87.8000 209.0000 88.2000 ;
	    RECT 206.2000 87.1000 206.6000 87.2000 ;
	    RECT 207.0000 87.1000 207.4000 87.2000 ;
	    RECT 206.2000 86.8000 207.4000 87.1000 ;
	    RECT 207.0000 86.1000 207.4000 86.2000 ;
	    RECT 207.8000 86.1000 208.2000 86.2000 ;
	    RECT 207.0000 85.8000 208.2000 86.1000 ;
	    RECT 209.4000 85.8000 209.8000 86.2000 ;
	    RECT 212.6000 86.1000 213.0000 86.2000 ;
	    RECT 213.4000 86.1000 213.8000 86.2000 ;
	    RECT 212.6000 85.8000 213.8000 86.1000 ;
	    RECT 203.8000 84.8000 204.2000 85.2000 ;
	    RECT 204.6000 84.8000 205.0000 85.2000 ;
	    RECT 205.4000 84.8000 205.8000 85.2000 ;
	    RECT 208.6000 84.8000 209.0000 85.2000 ;
	    RECT 203.8000 83.2000 204.1000 84.8000 ;
	    RECT 204.6000 84.2000 204.9000 84.8000 ;
	    RECT 204.6000 83.8000 205.0000 84.2000 ;
	    RECT 203.8000 82.8000 204.2000 83.2000 ;
	    RECT 205.4000 81.8000 205.8000 82.2000 ;
	    RECT 204.6000 79.8000 205.0000 80.2000 ;
	    RECT 203.0000 75.8000 203.4000 76.2000 ;
	    RECT 204.6000 74.2000 204.9000 79.8000 ;
	    RECT 205.4000 77.2000 205.7000 81.8000 ;
	    RECT 208.6000 81.2000 208.9000 84.8000 ;
	    RECT 208.6000 80.8000 209.0000 81.2000 ;
	    RECT 205.4000 76.8000 205.8000 77.2000 ;
	    RECT 207.8000 75.8000 208.2000 76.2000 ;
	    RECT 207.8000 75.2000 208.1000 75.8000 ;
	    RECT 205.4000 75.1000 205.8000 75.2000 ;
	    RECT 206.2000 75.1000 206.6000 75.2000 ;
	    RECT 205.4000 74.8000 206.6000 75.1000 ;
	    RECT 207.8000 74.8000 208.2000 75.2000 ;
	    RECT 202.2000 73.8000 202.6000 74.2000 ;
	    RECT 204.6000 73.8000 205.0000 74.2000 ;
	    RECT 206.2000 73.8000 206.6000 74.2000 ;
	    RECT 207.0000 74.1000 207.4000 74.2000 ;
	    RECT 207.8000 74.1000 208.2000 74.2000 ;
	    RECT 207.0000 73.8000 208.2000 74.1000 ;
	    RECT 202.2000 73.2000 202.5000 73.8000 ;
	    RECT 199.8000 72.8000 200.2000 73.2000 ;
	    RECT 202.2000 72.8000 202.6000 73.2000 ;
	    RECT 203.0000 73.1000 203.4000 73.2000 ;
	    RECT 203.8000 73.1000 204.2000 73.2000 ;
	    RECT 203.0000 72.8000 204.2000 73.1000 ;
	    RECT 204.6000 73.1000 205.0000 73.2000 ;
	    RECT 205.4000 73.1000 205.8000 73.2000 ;
	    RECT 204.6000 72.8000 205.8000 73.1000 ;
	    RECT 194.2000 71.8000 194.6000 72.2000 ;
	    RECT 194.2000 69.2000 194.5000 71.8000 ;
	    RECT 195.8000 70.8000 196.2000 71.2000 ;
	    RECT 195.8000 69.2000 196.1000 70.8000 ;
	    RECT 199.8000 70.1000 200.1000 72.8000 ;
	    RECT 199.0000 69.8000 200.1000 70.1000 ;
	    RECT 202.2000 71.8000 202.6000 72.2000 ;
	    RECT 202.2000 70.2000 202.5000 71.8000 ;
	    RECT 203.8000 70.8000 204.2000 71.2000 ;
	    RECT 202.2000 69.8000 202.6000 70.2000 ;
	    RECT 194.2000 68.8000 194.6000 69.2000 ;
	    RECT 195.8000 68.8000 196.2000 69.2000 ;
	    RECT 195.0000 67.5000 195.4000 67.9000 ;
	    RECT 195.7000 67.5000 197.8000 67.8000 ;
	    RECT 198.3000 67.5000 198.7000 67.9000 ;
	    RECT 187.0000 66.8000 188.1000 67.1000 ;
	    RECT 190.2000 66.8000 190.6000 67.2000 ;
	    RECT 191.8000 66.8000 192.2000 67.2000 ;
	    RECT 193.4000 67.1000 193.8000 67.2000 ;
	    RECT 194.2000 67.1000 194.6000 67.2000 ;
	    RECT 193.4000 66.8000 194.6000 67.1000 ;
	    RECT 195.0000 67.1000 195.3000 67.5000 ;
	    RECT 195.7000 67.4000 196.1000 67.5000 ;
	    RECT 197.4000 67.4000 197.8000 67.5000 ;
	    RECT 195.0000 66.8000 197.4000 67.1000 ;
	    RECT 176.6000 64.8000 177.7000 65.1000 ;
	    RECT 178.2000 65.8000 178.6000 66.2000 ;
	    RECT 179.8000 66.1000 180.2000 66.2000 ;
	    RECT 180.6000 66.1000 181.0000 66.2000 ;
	    RECT 179.8000 65.8000 181.0000 66.1000 ;
	    RECT 178.2000 64.1000 178.5000 65.8000 ;
	    RECT 177.4000 63.8000 178.5000 64.1000 ;
	    RECT 177.4000 59.2000 177.7000 63.8000 ;
	    RECT 180.6000 61.8000 181.0000 62.2000 ;
	    RECT 177.4000 58.8000 177.8000 59.2000 ;
	    RECT 180.6000 57.2000 180.9000 61.8000 ;
	    RECT 175.8000 56.8000 176.2000 57.2000 ;
	    RECT 180.6000 56.8000 181.0000 57.2000 ;
	    RECT 172.6000 55.8000 173.0000 56.2000 ;
	    RECT 175.8000 55.2000 176.1000 56.8000 ;
	    RECT 179.0000 56.1000 179.4000 56.2000 ;
	    RECT 179.8000 56.1000 180.2000 56.2000 ;
	    RECT 179.0000 55.8000 180.2000 56.1000 ;
	    RECT 181.4000 55.2000 181.7000 66.8000 ;
	    RECT 190.2000 66.2000 190.5000 66.8000 ;
	    RECT 185.4000 66.1000 185.8000 66.2000 ;
	    RECT 186.2000 66.1000 186.6000 66.2000 ;
	    RECT 185.4000 65.8000 186.6000 66.1000 ;
	    RECT 188.6000 66.1000 189.0000 66.2000 ;
	    RECT 189.4000 66.1000 189.8000 66.2000 ;
	    RECT 188.6000 65.8000 189.8000 66.1000 ;
	    RECT 190.2000 65.8000 190.6000 66.2000 ;
	    RECT 191.8000 66.1000 192.2000 66.2000 ;
	    RECT 192.6000 66.1000 193.0000 66.2000 ;
	    RECT 191.8000 65.8000 193.0000 66.1000 ;
	    RECT 193.4000 65.8000 193.8000 66.2000 ;
	    RECT 191.0000 61.8000 191.4000 62.2000 ;
	    RECT 183.0000 56.8000 183.4000 57.2000 ;
	    RECT 183.0000 55.2000 183.3000 56.8000 ;
	    RECT 175.8000 54.8000 176.2000 55.2000 ;
	    RECT 177.4000 54.8000 177.8000 55.2000 ;
	    RECT 178.2000 54.8000 178.6000 55.2000 ;
	    RECT 181.4000 54.8000 181.8000 55.2000 ;
	    RECT 183.0000 54.8000 183.4000 55.2000 ;
	    RECT 172.6000 54.1000 173.0000 54.2000 ;
	    RECT 173.4000 54.1000 173.8000 54.2000 ;
	    RECT 172.6000 53.8000 173.8000 54.1000 ;
	    RECT 174.2000 54.1000 174.6000 54.2000 ;
	    RECT 175.0000 54.1000 175.4000 54.2000 ;
	    RECT 174.2000 53.8000 175.4000 54.1000 ;
	    RECT 173.4000 52.8000 173.8000 53.2000 ;
	    RECT 175.8000 53.1000 176.2000 53.2000 ;
	    RECT 176.6000 53.1000 177.0000 53.2000 ;
	    RECT 175.8000 52.8000 177.0000 53.1000 ;
	    RECT 173.4000 52.2000 173.7000 52.8000 ;
	    RECT 173.4000 51.8000 173.8000 52.2000 ;
	    RECT 174.2000 51.8000 174.6000 52.2000 ;
	    RECT 176.6000 51.8000 177.0000 52.2000 ;
	    RECT 171.8000 47.8000 172.2000 48.2000 ;
	    RECT 171.8000 46.2000 172.2000 46.3000 ;
	    RECT 172.6000 46.2000 173.0000 46.3000 ;
	    RECT 169.4000 45.8000 169.8000 46.2000 ;
	    RECT 171.8000 45.9000 173.0000 46.2000 ;
	    RECT 169.4000 42.1000 169.7000 45.8000 ;
	    RECT 173.4000 43.1000 173.8000 48.9000 ;
	    RECT 174.2000 46.2000 174.5000 51.8000 ;
	    RECT 176.6000 49.2000 176.9000 51.8000 ;
	    RECT 177.4000 49.2000 177.7000 54.8000 ;
	    RECT 178.2000 54.2000 178.5000 54.8000 ;
	    RECT 178.2000 53.8000 178.6000 54.2000 ;
	    RECT 179.8000 54.1000 180.2000 54.2000 ;
	    RECT 180.6000 54.1000 181.0000 54.2000 ;
	    RECT 179.8000 53.8000 181.0000 54.1000 ;
	    RECT 181.4000 54.1000 181.8000 54.2000 ;
	    RECT 182.2000 54.1000 182.6000 54.2000 ;
	    RECT 181.4000 53.8000 182.6000 54.1000 ;
	    RECT 183.0000 53.8000 183.4000 54.2000 ;
	    RECT 180.6000 52.8000 181.0000 53.2000 ;
	    RECT 180.6000 52.2000 180.9000 52.8000 ;
	    RECT 180.6000 51.8000 181.0000 52.2000 ;
	    RECT 181.4000 51.8000 181.8000 52.2000 ;
	    RECT 175.8000 48.8000 176.2000 49.2000 ;
	    RECT 176.6000 48.8000 177.0000 49.2000 ;
	    RECT 177.4000 48.8000 177.8000 49.2000 ;
	    RECT 175.8000 48.2000 176.1000 48.8000 ;
	    RECT 174.2000 45.8000 174.6000 46.2000 ;
	    RECT 175.0000 45.1000 175.4000 47.9000 ;
	    RECT 175.8000 47.8000 176.2000 48.2000 ;
	    RECT 174.2000 43.8000 174.6000 44.2000 ;
	    RECT 168.6000 41.8000 169.7000 42.1000 ;
	    RECT 164.6000 36.8000 165.0000 37.2000 ;
	    RECT 163.8000 34.8000 164.2000 35.2000 ;
	    RECT 163.8000 34.2000 164.1000 34.8000 ;
	    RECT 167.0000 34.7000 167.4000 35.1000 ;
	    RECT 167.0000 34.2000 167.3000 34.7000 ;
	    RECT 163.8000 33.8000 164.2000 34.2000 ;
	    RECT 167.0000 33.8000 167.4000 34.2000 ;
	    RECT 167.8000 32.1000 168.2000 37.9000 ;
	    RECT 168.6000 34.2000 168.9000 41.8000 ;
	    RECT 174.2000 39.2000 174.5000 43.8000 ;
	    RECT 179.8000 43.1000 180.2000 48.9000 ;
	    RECT 181.4000 46.2000 181.7000 51.8000 ;
	    RECT 183.0000 47.2000 183.3000 53.8000 ;
	    RECT 183.8000 53.1000 184.2000 55.9000 ;
	    RECT 185.4000 52.1000 185.8000 57.9000 ;
	    RECT 186.2000 55.8000 186.6000 56.2000 ;
	    RECT 186.2000 55.1000 186.5000 55.8000 ;
	    RECT 186.2000 54.7000 186.6000 55.1000 ;
	    RECT 189.4000 54.8000 189.8000 55.2000 ;
	    RECT 189.4000 51.2000 189.7000 54.8000 ;
	    RECT 190.2000 52.1000 190.6000 57.9000 ;
	    RECT 191.0000 57.2000 191.3000 61.8000 ;
	    RECT 192.6000 59.8000 193.0000 60.2000 ;
	    RECT 192.6000 59.2000 192.9000 59.8000 ;
	    RECT 193.4000 59.2000 193.7000 65.8000 ;
	    RECT 194.2000 59.2000 194.5000 66.8000 ;
	    RECT 195.0000 65.1000 195.3000 66.8000 ;
	    RECT 197.0000 66.7000 197.4000 66.8000 ;
	    RECT 198.4000 65.1000 198.7000 67.5000 ;
	    RECT 199.0000 67.2000 199.3000 69.8000 ;
	    RECT 202.2000 67.2000 202.5000 69.8000 ;
	    RECT 203.8000 69.2000 204.1000 70.8000 ;
	    RECT 206.2000 70.2000 206.5000 73.8000 ;
	    RECT 206.2000 69.8000 206.6000 70.2000 ;
	    RECT 203.8000 68.8000 204.2000 69.2000 ;
	    RECT 205.4000 68.8000 205.8000 69.2000 ;
	    RECT 205.4000 68.2000 205.7000 68.8000 ;
	    RECT 205.4000 67.8000 205.8000 68.2000 ;
	    RECT 206.2000 67.2000 206.5000 69.8000 ;
	    RECT 208.6000 69.2000 208.9000 80.8000 ;
	    RECT 209.4000 76.2000 209.7000 85.8000 ;
	    RECT 215.0000 85.2000 215.3000 89.8000 ;
	    RECT 215.0000 84.8000 215.4000 85.2000 ;
	    RECT 209.4000 75.8000 209.8000 76.2000 ;
	    RECT 210.2000 73.1000 210.6000 75.9000 ;
	    RECT 211.0000 73.8000 211.4000 74.2000 ;
	    RECT 211.0000 73.2000 211.3000 73.8000 ;
	    RECT 211.0000 72.8000 211.4000 73.2000 ;
	    RECT 209.4000 71.8000 209.8000 72.2000 ;
	    RECT 211.8000 72.1000 212.2000 77.9000 ;
	    RECT 212.6000 75.0000 213.0000 75.1000 ;
	    RECT 213.4000 75.0000 213.8000 75.1000 ;
	    RECT 212.6000 74.7000 213.8000 75.0000 ;
	    RECT 215.8000 73.2000 216.1000 93.8000 ;
	    RECT 216.7000 93.5000 217.0000 95.9000 ;
	    RECT 217.3000 94.9000 217.7000 95.3000 ;
	    RECT 217.4000 94.2000 217.7000 94.9000 ;
	    RECT 219.9000 94.2000 220.2000 95.9000 ;
	    RECT 223.8000 95.2000 224.1000 97.8000 ;
	    RECT 225.4000 96.2000 225.7000 98.8000 ;
	    RECT 227.8000 96.2000 228.1000 111.8000 ;
	    RECT 231.8000 111.2000 232.1000 111.8000 ;
	    RECT 231.8000 110.8000 232.2000 111.2000 ;
	    RECT 228.6000 109.1000 229.0000 109.2000 ;
	    RECT 229.4000 109.1000 229.8000 109.2000 ;
	    RECT 228.6000 108.8000 229.8000 109.1000 ;
	    RECT 230.2000 108.8000 230.6000 109.2000 ;
	    RECT 230.2000 108.2000 230.5000 108.8000 ;
	    RECT 232.6000 108.2000 232.9000 112.8000 ;
	    RECT 234.2000 111.8000 234.6000 112.2000 ;
	    RECT 236.6000 111.8000 237.0000 112.2000 ;
	    RECT 234.2000 110.2000 234.5000 111.8000 ;
	    RECT 234.2000 109.8000 234.6000 110.2000 ;
	    RECT 230.2000 107.8000 230.6000 108.2000 ;
	    RECT 231.8000 108.1000 232.2000 108.2000 ;
	    RECT 232.6000 108.1000 233.0000 108.2000 ;
	    RECT 231.8000 107.8000 233.0000 108.1000 ;
	    RECT 234.2000 108.1000 234.6000 108.2000 ;
	    RECT 235.0000 108.1000 235.4000 108.2000 ;
	    RECT 234.2000 107.8000 235.4000 108.1000 ;
	    RECT 236.6000 106.2000 236.9000 111.8000 ;
	    RECT 238.2000 110.1000 238.5000 122.8000 ;
	    RECT 239.0000 114.8000 239.4000 115.2000 ;
	    RECT 241.4000 114.8000 241.8000 115.2000 ;
	    RECT 239.0000 113.2000 239.3000 114.8000 ;
	    RECT 241.4000 114.2000 241.7000 114.8000 ;
	    RECT 241.4000 113.8000 241.8000 114.2000 ;
	    RECT 239.0000 112.8000 239.4000 113.2000 ;
	    RECT 242.2000 113.1000 242.5000 138.8000 ;
	    RECT 247.0000 137.2000 247.3000 145.8000 ;
	    RECT 249.4000 145.1000 249.8000 145.2000 ;
	    RECT 250.2000 145.1000 250.5000 150.8000 ;
	    RECT 253.4000 149.2000 253.7000 154.8000 ;
	    RECT 259.0000 154.2000 259.3000 158.8000 ;
	    RECT 261.4000 158.2000 261.7000 165.8000 ;
	    RECT 261.4000 157.8000 261.8000 158.2000 ;
	    RECT 254.2000 153.8000 254.6000 154.2000 ;
	    RECT 259.0000 153.8000 259.4000 154.2000 ;
	    RECT 254.2000 150.2000 254.5000 153.8000 ;
	    RECT 259.0000 153.2000 259.3000 153.8000 ;
	    RECT 259.0000 152.8000 259.4000 153.2000 ;
	    RECT 260.6000 153.1000 261.0000 153.2000 ;
	    RECT 261.4000 153.1000 261.8000 153.2000 ;
	    RECT 260.6000 152.8000 261.8000 153.1000 ;
	    RECT 262.2000 152.2000 262.5000 166.8000 ;
	    RECT 263.0000 165.1000 263.3000 166.8000 ;
	    RECT 265.5000 166.1000 265.8000 166.8000 ;
	    RECT 265.5000 165.7000 265.9000 166.1000 ;
	    RECT 266.2000 165.1000 266.5000 167.5000 ;
	    RECT 263.0000 164.7000 263.4000 165.1000 ;
	    RECT 266.1000 164.7000 266.5000 165.1000 ;
	    RECT 267.8000 165.8000 268.2000 166.2000 ;
	    RECT 267.8000 161.2000 268.1000 165.8000 ;
	    RECT 269.4000 161.8000 269.8000 162.2000 ;
	    RECT 267.8000 160.8000 268.2000 161.2000 ;
	    RECT 269.4000 156.2000 269.7000 161.8000 ;
	    RECT 263.8000 156.1000 264.2000 156.2000 ;
	    RECT 264.6000 156.1000 265.0000 156.2000 ;
	    RECT 263.8000 155.8000 265.0000 156.1000 ;
	    RECT 269.4000 155.8000 269.8000 156.2000 ;
	    RECT 262.2000 151.8000 262.6000 152.2000 ;
	    RECT 263.8000 150.2000 264.1000 155.8000 ;
	    RECT 264.6000 154.1000 265.0000 154.2000 ;
	    RECT 265.4000 154.1000 265.8000 154.2000 ;
	    RECT 264.6000 153.8000 265.8000 154.1000 ;
	    RECT 268.6000 153.1000 269.0000 153.2000 ;
	    RECT 267.8000 152.8000 269.0000 153.1000 ;
	    RECT 266.2000 151.8000 266.6000 152.2000 ;
	    RECT 254.2000 149.8000 254.6000 150.2000 ;
	    RECT 261.4000 149.8000 261.8000 150.2000 ;
	    RECT 263.8000 149.8000 264.2000 150.2000 ;
	    RECT 251.0000 148.8000 251.4000 149.2000 ;
	    RECT 253.4000 148.8000 253.8000 149.2000 ;
	    RECT 251.0000 146.2000 251.3000 148.8000 ;
	    RECT 257.4000 147.8000 257.8000 148.2000 ;
	    RECT 258.2000 148.1000 258.6000 148.2000 ;
	    RECT 259.0000 148.1000 259.4000 148.2000 ;
	    RECT 258.2000 147.8000 259.4000 148.1000 ;
	    RECT 251.8000 146.8000 252.2000 147.2000 ;
	    RECT 252.6000 147.1000 253.0000 147.2000 ;
	    RECT 253.4000 147.1000 253.8000 147.2000 ;
	    RECT 252.6000 146.8000 253.8000 147.1000 ;
	    RECT 254.2000 146.8000 254.6000 147.2000 ;
	    RECT 257.4000 147.0000 257.7000 147.8000 ;
	    RECT 251.0000 145.8000 251.4000 146.2000 ;
	    RECT 251.8000 145.2000 252.1000 146.8000 ;
	    RECT 254.2000 146.2000 254.5000 146.8000 ;
	    RECT 257.4000 146.6000 257.8000 147.0000 ;
	    RECT 258.2000 146.8000 258.6000 147.2000 ;
	    RECT 259.0000 146.8000 259.4000 147.2000 ;
	    RECT 258.2000 146.2000 258.5000 146.8000 ;
	    RECT 259.0000 146.2000 259.3000 146.8000 ;
	    RECT 261.4000 146.2000 261.7000 149.8000 ;
	    RECT 263.8000 148.8000 264.2000 149.2000 ;
	    RECT 263.8000 147.2000 264.1000 148.8000 ;
	    RECT 264.6000 147.8000 265.0000 148.2000 ;
	    RECT 266.2000 148.1000 266.5000 151.8000 ;
	    RECT 266.2000 147.8000 267.3000 148.1000 ;
	    RECT 264.6000 147.2000 264.9000 147.8000 ;
	    RECT 263.0000 146.8000 263.4000 147.2000 ;
	    RECT 263.8000 146.8000 264.2000 147.2000 ;
	    RECT 264.6000 146.8000 265.0000 147.2000 ;
	    RECT 266.2000 146.8000 266.6000 147.2000 ;
	    RECT 263.0000 146.2000 263.3000 146.8000 ;
	    RECT 252.6000 145.8000 253.0000 146.2000 ;
	    RECT 254.2000 145.8000 254.6000 146.2000 ;
	    RECT 258.2000 145.8000 258.6000 146.2000 ;
	    RECT 259.0000 145.8000 259.4000 146.2000 ;
	    RECT 261.4000 145.8000 261.8000 146.2000 ;
	    RECT 262.2000 145.8000 262.6000 146.2000 ;
	    RECT 263.0000 145.8000 263.4000 146.2000 ;
	    RECT 264.6000 146.1000 265.0000 146.2000 ;
	    RECT 265.4000 146.1000 265.8000 146.2000 ;
	    RECT 264.6000 145.8000 265.8000 146.1000 ;
	    RECT 252.6000 145.2000 252.9000 145.8000 ;
	    RECT 249.4000 144.8000 250.5000 145.1000 ;
	    RECT 251.0000 144.8000 251.4000 145.2000 ;
	    RECT 251.8000 144.8000 252.2000 145.2000 ;
	    RECT 252.6000 144.8000 253.0000 145.2000 ;
	    RECT 255.0000 144.8000 255.4000 145.2000 ;
	    RECT 251.0000 144.2000 251.3000 144.8000 ;
	    RECT 251.0000 143.8000 251.4000 144.2000 ;
	    RECT 255.0000 139.2000 255.3000 144.8000 ;
	    RECT 256.6000 139.8000 257.0000 140.2000 ;
	    RECT 255.0000 138.8000 255.4000 139.2000 ;
	    RECT 255.0000 137.8000 255.4000 138.2000 ;
	    RECT 247.0000 136.8000 247.4000 137.2000 ;
	    RECT 247.8000 136.8000 248.2000 137.2000 ;
	    RECT 249.4000 136.8000 249.8000 137.2000 ;
	    RECT 245.4000 136.1000 245.8000 136.2000 ;
	    RECT 246.2000 136.1000 246.6000 136.2000 ;
	    RECT 245.4000 135.8000 246.6000 136.1000 ;
	    RECT 247.8000 135.2000 248.1000 136.8000 ;
	    RECT 249.4000 136.2000 249.7000 136.8000 ;
	    RECT 249.4000 135.8000 249.8000 136.2000 ;
	    RECT 251.0000 135.8000 251.4000 136.2000 ;
	    RECT 251.0000 135.2000 251.3000 135.8000 ;
	    RECT 255.0000 135.2000 255.3000 137.8000 ;
	    RECT 256.6000 136.2000 256.9000 139.8000 ;
	    RECT 258.2000 136.2000 258.5000 145.8000 ;
	    RECT 261.4000 144.8000 261.8000 145.2000 ;
	    RECT 261.4000 142.2000 261.7000 144.8000 ;
	    RECT 261.4000 141.8000 261.8000 142.2000 ;
	    RECT 262.2000 140.2000 262.5000 145.8000 ;
	    RECT 262.2000 139.8000 262.6000 140.2000 ;
	    RECT 266.2000 139.2000 266.5000 146.8000 ;
	    RECT 266.2000 138.8000 266.6000 139.2000 ;
	    RECT 259.0000 137.8000 259.4000 138.2000 ;
	    RECT 259.0000 137.2000 259.3000 137.8000 ;
	    RECT 259.0000 136.8000 259.4000 137.2000 ;
	    RECT 256.6000 135.8000 257.0000 136.2000 ;
	    RECT 257.4000 135.8000 257.8000 136.2000 ;
	    RECT 258.2000 135.8000 258.6000 136.2000 ;
	    RECT 260.6000 135.8000 261.0000 136.2000 ;
	    RECT 266.2000 135.8000 266.6000 136.2000 ;
	    RECT 245.4000 135.1000 245.8000 135.2000 ;
	    RECT 246.2000 135.1000 246.6000 135.2000 ;
	    RECT 245.4000 134.8000 246.6000 135.1000 ;
	    RECT 247.8000 134.8000 248.2000 135.2000 ;
	    RECT 248.6000 134.8000 249.0000 135.2000 ;
	    RECT 249.4000 135.1000 249.8000 135.2000 ;
	    RECT 250.2000 135.1000 250.6000 135.2000 ;
	    RECT 249.4000 134.8000 250.6000 135.1000 ;
	    RECT 251.0000 134.8000 251.4000 135.2000 ;
	    RECT 251.8000 135.1000 252.2000 135.2000 ;
	    RECT 252.6000 135.1000 253.0000 135.2000 ;
	    RECT 251.8000 134.8000 253.0000 135.1000 ;
	    RECT 253.4000 134.8000 253.8000 135.2000 ;
	    RECT 255.0000 134.8000 255.4000 135.2000 ;
	    RECT 247.0000 133.8000 247.4000 134.2000 ;
	    RECT 243.0000 132.8000 243.4000 133.2000 ;
	    RECT 243.0000 129.2000 243.3000 132.8000 ;
	    RECT 245.4000 131.8000 245.8000 132.2000 ;
	    RECT 245.4000 129.2000 245.7000 131.8000 ;
	    RECT 243.0000 128.8000 243.4000 129.2000 ;
	    RECT 245.4000 128.8000 245.8000 129.2000 ;
	    RECT 247.0000 128.2000 247.3000 133.8000 ;
	    RECT 243.0000 127.8000 243.4000 128.2000 ;
	    RECT 247.0000 127.8000 247.4000 128.2000 ;
	    RECT 243.0000 125.2000 243.3000 127.8000 ;
	    RECT 248.6000 126.2000 248.9000 134.8000 ;
	    RECT 253.4000 134.2000 253.7000 134.8000 ;
	    RECT 250.2000 133.8000 250.6000 134.2000 ;
	    RECT 253.4000 133.8000 253.8000 134.2000 ;
	    RECT 254.2000 133.8000 254.6000 134.2000 ;
	    RECT 256.6000 133.8000 257.0000 134.2000 ;
	    RECT 250.2000 132.2000 250.5000 133.8000 ;
	    RECT 254.2000 133.2000 254.5000 133.8000 ;
	    RECT 252.6000 132.8000 253.0000 133.2000 ;
	    RECT 254.2000 132.8000 254.6000 133.2000 ;
	    RECT 252.6000 132.2000 252.9000 132.8000 ;
	    RECT 250.2000 131.8000 250.6000 132.2000 ;
	    RECT 252.6000 131.8000 253.0000 132.2000 ;
	    RECT 255.0000 130.8000 255.4000 131.2000 ;
	    RECT 253.4000 128.8000 253.8000 129.2000 ;
	    RECT 253.4000 128.2000 253.7000 128.8000 ;
	    RECT 255.0000 128.2000 255.3000 130.8000 ;
	    RECT 256.6000 129.2000 256.9000 133.8000 ;
	    RECT 257.4000 131.2000 257.7000 135.8000 ;
	    RECT 260.6000 135.2000 260.9000 135.8000 ;
	    RECT 266.2000 135.2000 266.5000 135.8000 ;
	    RECT 259.0000 134.8000 259.4000 135.2000 ;
	    RECT 259.8000 134.8000 260.2000 135.2000 ;
	    RECT 260.6000 134.8000 261.0000 135.2000 ;
	    RECT 262.2000 134.8000 262.6000 135.2000 ;
	    RECT 266.2000 134.8000 266.6000 135.2000 ;
	    RECT 259.0000 133.2000 259.3000 134.8000 ;
	    RECT 259.8000 134.2000 260.1000 134.8000 ;
	    RECT 262.2000 134.2000 262.5000 134.8000 ;
	    RECT 259.8000 133.8000 260.2000 134.2000 ;
	    RECT 260.6000 133.8000 261.0000 134.2000 ;
	    RECT 262.2000 133.8000 262.6000 134.2000 ;
	    RECT 265.4000 134.1000 265.8000 134.2000 ;
	    RECT 266.2000 134.1000 266.6000 134.2000 ;
	    RECT 265.4000 133.8000 266.6000 134.1000 ;
	    RECT 260.6000 133.2000 260.9000 133.8000 ;
	    RECT 259.0000 132.8000 259.4000 133.2000 ;
	    RECT 260.6000 132.8000 261.0000 133.2000 ;
	    RECT 257.4000 130.8000 257.8000 131.2000 ;
	    RECT 257.4000 129.8000 257.8000 130.2000 ;
	    RECT 262.2000 129.8000 262.6000 130.2000 ;
	    RECT 255.8000 128.8000 256.2000 129.2000 ;
	    RECT 256.6000 128.8000 257.0000 129.2000 ;
	    RECT 255.8000 128.2000 256.1000 128.8000 ;
	    RECT 253.4000 127.8000 253.8000 128.2000 ;
	    RECT 255.0000 127.8000 255.4000 128.2000 ;
	    RECT 255.8000 127.8000 256.2000 128.2000 ;
	    RECT 257.4000 127.2000 257.7000 129.8000 ;
	    RECT 262.2000 129.2000 262.5000 129.8000 ;
	    RECT 259.8000 128.8000 260.2000 129.2000 ;
	    RECT 262.2000 128.8000 262.6000 129.2000 ;
	    RECT 259.8000 128.2000 260.1000 128.8000 ;
	    RECT 259.0000 127.8000 259.4000 128.2000 ;
	    RECT 259.8000 127.8000 260.2000 128.2000 ;
	    RECT 263.0000 128.1000 263.4000 128.2000 ;
	    RECT 263.8000 128.1000 264.2000 128.2000 ;
	    RECT 263.0000 127.8000 264.2000 128.1000 ;
	    RECT 251.0000 126.8000 251.4000 127.2000 ;
	    RECT 257.4000 126.8000 257.8000 127.2000 ;
	    RECT 244.6000 126.1000 245.0000 126.2000 ;
	    RECT 245.4000 126.1000 245.8000 126.2000 ;
	    RECT 244.6000 125.8000 245.8000 126.1000 ;
	    RECT 248.6000 126.1000 249.0000 126.2000 ;
	    RECT 249.4000 126.1000 249.8000 126.2000 ;
	    RECT 248.6000 125.8000 249.8000 126.1000 ;
	    RECT 243.0000 124.8000 243.4000 125.2000 ;
	    RECT 243.8000 124.8000 244.2000 125.2000 ;
	    RECT 243.0000 124.2000 243.3000 124.8000 ;
	    RECT 243.8000 124.2000 244.1000 124.8000 ;
	    RECT 243.0000 123.8000 243.4000 124.2000 ;
	    RECT 243.8000 123.8000 244.2000 124.2000 ;
	    RECT 251.0000 123.2000 251.3000 126.8000 ;
	    RECT 258.2000 125.8000 258.6000 126.2000 ;
	    RECT 258.2000 125.2000 258.5000 125.8000 ;
	    RECT 258.2000 124.8000 258.6000 125.2000 ;
	    RECT 251.0000 122.8000 251.4000 123.2000 ;
	    RECT 259.0000 121.2000 259.3000 127.8000 ;
	    RECT 261.4000 127.1000 261.8000 127.2000 ;
	    RECT 262.2000 127.1000 262.6000 127.2000 ;
	    RECT 261.4000 126.8000 262.6000 127.1000 ;
	    RECT 264.6000 126.8000 265.0000 127.2000 ;
	    RECT 259.0000 120.8000 259.4000 121.2000 ;
	    RECT 243.0000 119.8000 243.4000 120.2000 ;
	    RECT 243.0000 116.2000 243.3000 119.8000 ;
	    RECT 264.6000 119.2000 264.9000 126.8000 ;
	    RECT 266.2000 126.2000 266.5000 133.8000 ;
	    RECT 267.0000 127.2000 267.3000 147.8000 ;
	    RECT 267.8000 139.2000 268.1000 152.8000 ;
	    RECT 268.6000 149.1000 269.0000 149.2000 ;
	    RECT 269.4000 149.1000 269.8000 149.2000 ;
	    RECT 268.6000 148.8000 269.8000 149.1000 ;
	    RECT 270.2000 148.8000 270.6000 149.2000 ;
	    RECT 270.2000 148.2000 270.5000 148.8000 ;
	    RECT 268.6000 147.8000 269.0000 148.2000 ;
	    RECT 270.2000 147.8000 270.6000 148.2000 ;
	    RECT 268.6000 147.2000 268.9000 147.8000 ;
	    RECT 268.6000 146.8000 269.0000 147.2000 ;
	    RECT 268.6000 145.8000 269.0000 146.2000 ;
	    RECT 268.6000 145.2000 268.9000 145.8000 ;
	    RECT 268.6000 144.8000 269.0000 145.2000 ;
	    RECT 267.8000 138.8000 268.2000 139.2000 ;
	    RECT 267.8000 134.1000 268.2000 134.2000 ;
	    RECT 268.6000 134.1000 269.0000 134.2000 ;
	    RECT 267.8000 133.8000 269.0000 134.1000 ;
	    RECT 267.0000 126.8000 267.4000 127.2000 ;
	    RECT 266.2000 125.8000 266.6000 126.2000 ;
	    RECT 266.2000 125.1000 266.5000 125.8000 ;
	    RECT 267.0000 125.1000 267.4000 125.2000 ;
	    RECT 266.2000 124.8000 267.4000 125.1000 ;
	    RECT 255.0000 118.8000 255.4000 119.2000 ;
	    RECT 264.6000 118.8000 265.0000 119.2000 ;
	    RECT 252.6000 117.8000 253.0000 118.2000 ;
	    RECT 243.0000 115.8000 243.4000 116.2000 ;
	    RECT 247.0000 116.1000 247.4000 116.2000 ;
	    RECT 247.8000 116.1000 248.2000 116.2000 ;
	    RECT 247.0000 115.8000 248.2000 116.1000 ;
	    RECT 246.2000 114.8000 246.6000 115.2000 ;
	    RECT 247.8000 115.1000 248.2000 115.2000 ;
	    RECT 248.6000 115.1000 249.0000 115.2000 ;
	    RECT 247.8000 114.8000 249.0000 115.1000 ;
	    RECT 251.0000 114.8000 251.4000 115.2000 ;
	    RECT 246.2000 114.2000 246.5000 114.8000 ;
	    RECT 247.8000 114.2000 248.1000 114.8000 ;
	    RECT 251.0000 114.2000 251.3000 114.8000 ;
	    RECT 241.4000 112.8000 242.5000 113.1000 ;
	    RECT 245.4000 113.8000 245.8000 114.2000 ;
	    RECT 246.2000 113.8000 246.6000 114.2000 ;
	    RECT 247.8000 113.8000 248.2000 114.2000 ;
	    RECT 250.2000 113.8000 250.6000 114.2000 ;
	    RECT 251.0000 113.8000 251.4000 114.2000 ;
	    RECT 245.4000 113.2000 245.7000 113.8000 ;
	    RECT 250.2000 113.2000 250.5000 113.8000 ;
	    RECT 252.6000 113.2000 252.9000 117.8000 ;
	    RECT 253.4000 115.8000 253.8000 116.2000 ;
	    RECT 254.2000 115.8000 254.6000 116.2000 ;
	    RECT 253.4000 115.2000 253.7000 115.8000 ;
	    RECT 254.2000 115.2000 254.5000 115.8000 ;
	    RECT 253.4000 114.8000 253.8000 115.2000 ;
	    RECT 254.2000 114.8000 254.6000 115.2000 ;
	    RECT 255.0000 113.2000 255.3000 118.8000 ;
	    RECT 255.8000 116.8000 256.2000 117.2000 ;
	    RECT 255.8000 115.2000 256.1000 116.8000 ;
	    RECT 267.0000 116.2000 267.3000 124.8000 ;
	    RECT 258.2000 115.8000 258.6000 116.2000 ;
	    RECT 263.0000 115.8000 263.4000 116.2000 ;
	    RECT 266.2000 115.8000 266.6000 116.2000 ;
	    RECT 267.0000 115.8000 267.4000 116.2000 ;
	    RECT 258.2000 115.2000 258.5000 115.8000 ;
	    RECT 263.0000 115.2000 263.3000 115.8000 ;
	    RECT 255.8000 114.8000 256.2000 115.2000 ;
	    RECT 258.2000 114.8000 258.6000 115.2000 ;
	    RECT 263.0000 114.8000 263.4000 115.2000 ;
	    RECT 266.2000 114.2000 266.5000 115.8000 ;
	    RECT 257.4000 114.1000 257.8000 114.2000 ;
	    RECT 258.2000 114.1000 258.6000 114.2000 ;
	    RECT 257.4000 113.8000 258.6000 114.1000 ;
	    RECT 259.8000 114.1000 260.2000 114.2000 ;
	    RECT 260.6000 114.1000 261.0000 114.2000 ;
	    RECT 259.8000 113.8000 261.0000 114.1000 ;
	    RECT 262.2000 114.1000 262.6000 114.2000 ;
	    RECT 263.0000 114.1000 263.4000 114.2000 ;
	    RECT 262.2000 113.8000 263.4000 114.1000 ;
	    RECT 263.8000 114.1000 264.2000 114.2000 ;
	    RECT 263.8000 113.8000 264.9000 114.1000 ;
	    RECT 266.2000 113.8000 266.6000 114.2000 ;
	    RECT 245.4000 112.8000 245.8000 113.2000 ;
	    RECT 250.2000 112.8000 250.6000 113.2000 ;
	    RECT 252.6000 112.8000 253.0000 113.2000 ;
	    RECT 255.0000 112.8000 255.4000 113.2000 ;
	    RECT 256.6000 113.1000 257.0000 113.2000 ;
	    RECT 257.4000 113.1000 257.8000 113.2000 ;
	    RECT 256.6000 112.8000 257.8000 113.1000 ;
	    RECT 240.6000 111.8000 241.0000 112.2000 ;
	    RECT 238.2000 109.8000 239.3000 110.1000 ;
	    RECT 239.0000 108.2000 239.3000 109.8000 ;
	    RECT 239.0000 107.8000 239.4000 108.2000 ;
	    RECT 231.0000 106.1000 231.4000 106.2000 ;
	    RECT 231.8000 106.1000 232.2000 106.2000 ;
	    RECT 231.0000 105.8000 232.9000 106.1000 ;
	    RECT 230.2000 99.8000 230.6000 100.2000 ;
	    RECT 225.4000 95.8000 225.8000 96.2000 ;
	    RECT 227.8000 95.8000 228.2000 96.2000 ;
	    RECT 217.4000 93.9000 220.2000 94.2000 ;
	    RECT 217.4000 93.5000 217.8000 93.6000 ;
	    RECT 219.1000 93.5000 219.5000 93.6000 ;
	    RECT 219.9000 93.5000 220.2000 93.9000 ;
	    RECT 216.7000 93.2000 219.5000 93.5000 ;
	    RECT 216.7000 93.1000 217.1000 93.2000 ;
	    RECT 219.8000 93.1000 220.2000 93.5000 ;
	    RECT 221.4000 95.1000 221.8000 95.2000 ;
	    RECT 222.2000 95.1000 222.6000 95.2000 ;
	    RECT 221.4000 94.8000 222.6000 95.1000 ;
	    RECT 223.8000 94.8000 224.2000 95.2000 ;
	    RECT 217.4000 92.1000 217.8000 92.2000 ;
	    RECT 218.2000 92.1000 218.6000 92.2000 ;
	    RECT 217.4000 91.8000 218.6000 92.1000 ;
	    RECT 219.0000 88.1000 219.4000 88.2000 ;
	    RECT 219.8000 88.1000 220.2000 88.2000 ;
	    RECT 219.0000 87.8000 220.2000 88.1000 ;
	    RECT 221.4000 87.2000 221.7000 94.8000 ;
	    RECT 230.2000 94.2000 230.5000 99.8000 ;
	    RECT 231.0000 96.8000 231.4000 97.2000 ;
	    RECT 231.0000 96.2000 231.3000 96.8000 ;
	    RECT 231.0000 95.8000 231.4000 96.2000 ;
	    RECT 232.6000 95.2000 232.9000 105.8000 ;
	    RECT 233.4000 105.8000 233.8000 106.2000 ;
	    RECT 234.2000 106.1000 234.6000 106.2000 ;
	    RECT 235.0000 106.1000 235.4000 106.2000 ;
	    RECT 234.2000 105.8000 235.4000 106.1000 ;
	    RECT 236.6000 105.8000 237.0000 106.2000 ;
	    RECT 233.4000 105.2000 233.7000 105.8000 ;
	    RECT 233.4000 104.8000 233.8000 105.2000 ;
	    RECT 239.8000 103.8000 240.2000 104.2000 ;
	    RECT 239.8000 103.1000 240.1000 103.8000 ;
	    RECT 240.6000 103.1000 240.9000 111.8000 ;
	    RECT 239.8000 102.8000 240.9000 103.1000 ;
	    RECT 241.4000 107.2000 241.7000 112.8000 ;
	    RECT 242.2000 112.1000 242.6000 112.2000 ;
	    RECT 243.0000 112.1000 243.4000 112.2000 ;
	    RECT 242.2000 111.8000 243.4000 112.1000 ;
	    RECT 243.8000 111.8000 244.2000 112.2000 ;
	    RECT 247.0000 111.8000 247.4000 112.2000 ;
	    RECT 249.4000 111.8000 249.8000 112.2000 ;
	    RECT 251.8000 111.8000 252.2000 112.2000 ;
	    RECT 243.8000 111.2000 244.1000 111.8000 ;
	    RECT 243.0000 110.8000 243.4000 111.2000 ;
	    RECT 243.8000 110.8000 244.2000 111.2000 ;
	    RECT 243.0000 109.2000 243.3000 110.8000 ;
	    RECT 243.0000 108.8000 243.4000 109.2000 ;
	    RECT 242.3000 107.8000 242.7000 107.9000 ;
	    RECT 242.3000 107.5000 245.1000 107.8000 ;
	    RECT 245.4000 107.5000 245.8000 107.9000 ;
	    RECT 241.4000 106.8000 241.8000 107.2000 ;
	    RECT 235.8000 101.8000 236.2000 102.2000 ;
	    RECT 235.8000 96.2000 236.1000 101.8000 ;
	    RECT 239.8000 96.2000 240.1000 102.8000 ;
	    RECT 240.6000 101.8000 241.0000 102.2000 ;
	    RECT 240.6000 96.2000 240.9000 101.8000 ;
	    RECT 235.8000 95.8000 236.2000 96.2000 ;
	    RECT 239.8000 95.8000 240.2000 96.2000 ;
	    RECT 240.6000 95.8000 241.0000 96.2000 ;
	    RECT 241.4000 95.2000 241.7000 106.8000 ;
	    RECT 242.3000 105.1000 242.6000 107.5000 ;
	    RECT 243.0000 107.4000 243.4000 107.5000 ;
	    RECT 244.7000 107.4000 245.1000 107.5000 ;
	    RECT 245.5000 107.1000 245.8000 107.5000 ;
	    RECT 243.0000 106.8000 245.8000 107.1000 ;
	    RECT 243.0000 106.1000 243.3000 106.8000 ;
	    RECT 242.9000 105.7000 243.3000 106.1000 ;
	    RECT 245.5000 105.1000 245.8000 106.8000 ;
	    RECT 247.0000 106.2000 247.3000 111.8000 ;
	    RECT 248.6000 108.8000 249.0000 109.2000 ;
	    RECT 248.6000 108.2000 248.9000 108.8000 ;
	    RECT 248.6000 107.8000 249.0000 108.2000 ;
	    RECT 247.0000 105.8000 247.4000 106.2000 ;
	    RECT 247.8000 105.8000 248.2000 106.2000 ;
	    RECT 242.3000 104.7000 242.7000 105.1000 ;
	    RECT 245.4000 104.7000 245.8000 105.1000 ;
	    RECT 247.8000 105.2000 248.1000 105.8000 ;
	    RECT 247.8000 104.8000 248.2000 105.2000 ;
	    RECT 249.4000 105.1000 249.7000 111.8000 ;
	    RECT 248.6000 104.8000 249.7000 105.1000 ;
	    RECT 251.0000 106.8000 251.4000 107.2000 ;
	    RECT 243.8000 100.8000 244.2000 101.2000 ;
	    RECT 243.8000 95.2000 244.1000 100.8000 ;
	    RECT 247.0000 99.8000 247.4000 100.2000 ;
	    RECT 246.2000 96.8000 246.6000 97.2000 ;
	    RECT 232.6000 94.8000 233.0000 95.2000 ;
	    RECT 239.8000 94.8000 240.2000 95.2000 ;
	    RECT 241.4000 94.8000 241.8000 95.2000 ;
	    RECT 243.8000 94.8000 244.2000 95.2000 ;
	    RECT 230.2000 93.8000 230.6000 94.2000 ;
	    RECT 232.6000 94.1000 233.0000 94.2000 ;
	    RECT 233.4000 94.1000 233.8000 94.2000 ;
	    RECT 232.6000 93.8000 233.8000 94.1000 ;
	    RECT 235.0000 94.1000 235.4000 94.2000 ;
	    RECT 235.8000 94.1000 236.2000 94.2000 ;
	    RECT 235.0000 93.8000 236.2000 94.1000 ;
	    RECT 237.4000 94.1000 237.8000 94.2000 ;
	    RECT 238.2000 94.1000 238.6000 94.2000 ;
	    RECT 237.4000 93.8000 238.6000 94.1000 ;
	    RECT 239.0000 93.8000 239.4000 94.2000 ;
	    RECT 238.2000 93.2000 238.5000 93.8000 ;
	    RECT 239.0000 93.2000 239.3000 93.8000 ;
	    RECT 223.0000 93.1000 223.4000 93.2000 ;
	    RECT 223.0000 92.8000 224.1000 93.1000 ;
	    RECT 221.4000 86.8000 221.8000 87.2000 ;
	    RECT 222.2000 86.8000 222.6000 87.2000 ;
	    RECT 223.0000 86.8000 223.4000 87.2000 ;
	    RECT 222.2000 86.2000 222.5000 86.8000 ;
	    RECT 223.0000 86.2000 223.3000 86.8000 ;
	    RECT 217.4000 86.1000 217.8000 86.2000 ;
	    RECT 218.2000 86.1000 218.6000 86.2000 ;
	    RECT 217.4000 85.8000 218.6000 86.1000 ;
	    RECT 222.2000 85.8000 222.6000 86.2000 ;
	    RECT 223.0000 85.8000 223.4000 86.2000 ;
	    RECT 219.8000 82.8000 220.2000 83.2000 ;
	    RECT 217.4000 81.8000 217.8000 82.2000 ;
	    RECT 218.2000 81.8000 218.6000 82.2000 ;
	    RECT 215.8000 72.8000 216.2000 73.2000 ;
	    RECT 216.6000 72.1000 217.0000 77.9000 ;
	    RECT 217.4000 74.2000 217.7000 81.8000 ;
	    RECT 217.4000 73.8000 217.8000 74.2000 ;
	    RECT 208.6000 68.8000 209.0000 69.2000 ;
	    RECT 208.6000 68.2000 208.9000 68.8000 ;
	    RECT 208.6000 67.8000 209.0000 68.2000 ;
	    RECT 199.0000 66.8000 199.4000 67.2000 ;
	    RECT 202.2000 66.8000 202.6000 67.2000 ;
	    RECT 206.2000 66.8000 206.6000 67.2000 ;
	    RECT 199.0000 66.2000 199.3000 66.8000 ;
	    RECT 199.0000 65.8000 199.4000 66.2000 ;
	    RECT 209.4000 66.1000 209.7000 71.8000 ;
	    RECT 214.2000 67.8000 214.6000 68.2000 ;
	    RECT 214.2000 67.2000 214.5000 67.8000 ;
	    RECT 218.2000 67.2000 218.5000 81.8000 ;
	    RECT 219.8000 79.2000 220.1000 82.8000 ;
	    RECT 222.2000 79.2000 222.5000 85.8000 ;
	    RECT 219.8000 78.8000 220.2000 79.2000 ;
	    RECT 222.2000 78.8000 222.6000 79.2000 ;
	    RECT 223.8000 77.2000 224.1000 92.8000 ;
	    RECT 236.6000 92.8000 237.0000 93.2000 ;
	    RECT 238.2000 92.8000 238.6000 93.2000 ;
	    RECT 239.0000 92.8000 239.4000 93.2000 ;
	    RECT 236.6000 92.2000 236.9000 92.8000 ;
	    RECT 227.0000 91.8000 227.4000 92.2000 ;
	    RECT 231.0000 91.8000 231.4000 92.2000 ;
	    RECT 231.8000 91.8000 232.2000 92.2000 ;
	    RECT 236.6000 91.8000 237.0000 92.2000 ;
	    RECT 226.2000 88.8000 226.6000 89.2000 ;
	    RECT 224.6000 87.8000 225.0000 88.2000 ;
	    RECT 225.4000 87.8000 225.8000 88.2000 ;
	    RECT 224.6000 87.2000 224.9000 87.8000 ;
	    RECT 225.4000 87.2000 225.7000 87.8000 ;
	    RECT 224.6000 86.8000 225.0000 87.2000 ;
	    RECT 225.4000 86.8000 225.8000 87.2000 ;
	    RECT 226.2000 86.2000 226.5000 88.8000 ;
	    RECT 227.0000 88.2000 227.3000 91.8000 ;
	    RECT 229.4000 89.8000 229.8000 90.2000 ;
	    RECT 229.4000 88.2000 229.7000 89.8000 ;
	    RECT 231.0000 88.2000 231.3000 91.8000 ;
	    RECT 231.8000 91.2000 232.1000 91.8000 ;
	    RECT 231.8000 90.8000 232.2000 91.2000 ;
	    RECT 237.4000 90.8000 237.8000 91.2000 ;
	    RECT 237.4000 88.2000 237.7000 90.8000 ;
	    RECT 239.8000 89.2000 240.1000 94.8000 ;
	    RECT 241.4000 93.8000 241.8000 94.2000 ;
	    RECT 241.4000 93.2000 241.7000 93.8000 ;
	    RECT 246.2000 93.2000 246.5000 96.8000 ;
	    RECT 247.0000 93.2000 247.3000 99.8000 ;
	    RECT 248.6000 95.2000 248.9000 104.8000 ;
	    RECT 249.4000 103.8000 249.8000 104.2000 ;
	    RECT 249.4000 103.2000 249.7000 103.8000 ;
	    RECT 249.4000 102.8000 249.8000 103.2000 ;
	    RECT 250.2000 96.8000 250.6000 97.2000 ;
	    RECT 249.4000 95.8000 249.8000 96.2000 ;
	    RECT 249.4000 95.2000 249.7000 95.8000 ;
	    RECT 250.2000 95.2000 250.5000 96.8000 ;
	    RECT 248.6000 94.8000 249.0000 95.2000 ;
	    RECT 249.4000 94.8000 249.8000 95.2000 ;
	    RECT 250.2000 94.8000 250.6000 95.2000 ;
	    RECT 248.6000 94.2000 248.9000 94.8000 ;
	    RECT 248.6000 93.8000 249.0000 94.2000 ;
	    RECT 241.4000 93.1000 241.8000 93.2000 ;
	    RECT 242.2000 93.1000 242.6000 93.2000 ;
	    RECT 241.4000 92.8000 242.6000 93.1000 ;
	    RECT 246.2000 92.8000 246.6000 93.2000 ;
	    RECT 247.0000 92.8000 247.4000 93.2000 ;
	    RECT 240.6000 91.8000 241.0000 92.2000 ;
	    RECT 243.0000 91.8000 243.4000 92.2000 ;
	    RECT 245.4000 91.8000 245.8000 92.2000 ;
	    RECT 247.8000 91.8000 248.2000 92.2000 ;
	    RECT 239.8000 88.8000 240.2000 89.2000 ;
	    RECT 227.0000 87.8000 227.4000 88.2000 ;
	    RECT 229.4000 87.8000 229.8000 88.2000 ;
	    RECT 231.0000 87.8000 231.4000 88.2000 ;
	    RECT 231.8000 87.8000 232.2000 88.2000 ;
	    RECT 232.7000 87.8000 233.1000 87.9000 ;
	    RECT 231.8000 87.2000 232.1000 87.8000 ;
	    RECT 232.7000 87.5000 235.5000 87.8000 ;
	    RECT 235.8000 87.5000 236.2000 87.9000 ;
	    RECT 237.4000 87.8000 237.8000 88.2000 ;
	    RECT 240.6000 88.1000 240.9000 91.8000 ;
	    RECT 243.0000 90.2000 243.3000 91.8000 ;
	    RECT 243.0000 89.8000 243.4000 90.2000 ;
	    RECT 245.4000 89.2000 245.7000 91.8000 ;
	    RECT 243.0000 88.8000 243.4000 89.2000 ;
	    RECT 245.4000 88.8000 245.8000 89.2000 ;
	    RECT 241.4000 88.1000 241.8000 88.2000 ;
	    RECT 240.6000 87.8000 241.8000 88.1000 ;
	    RECT 227.0000 87.1000 227.4000 87.2000 ;
	    RECT 227.8000 87.1000 228.2000 87.2000 ;
	    RECT 227.0000 86.8000 228.2000 87.1000 ;
	    RECT 231.8000 86.8000 232.2000 87.2000 ;
	    RECT 226.2000 85.8000 226.6000 86.2000 ;
	    RECT 231.8000 84.8000 232.2000 85.2000 ;
	    RECT 232.7000 85.1000 233.0000 87.5000 ;
	    RECT 233.4000 87.4000 233.8000 87.5000 ;
	    RECT 235.1000 87.4000 235.5000 87.5000 ;
	    RECT 235.9000 87.1000 236.2000 87.5000 ;
	    RECT 243.0000 87.2000 243.3000 88.8000 ;
	    RECT 233.4000 86.8000 236.2000 87.1000 ;
	    RECT 233.4000 86.1000 233.7000 86.8000 ;
	    RECT 233.3000 85.7000 233.7000 86.1000 ;
	    RECT 234.2000 86.1000 234.6000 86.2000 ;
	    RECT 235.0000 86.1000 235.4000 86.2000 ;
	    RECT 234.2000 85.8000 235.4000 86.1000 ;
	    RECT 235.9000 85.1000 236.2000 86.8000 ;
	    RECT 239.0000 86.8000 239.4000 87.2000 ;
	    RECT 240.6000 86.8000 241.0000 87.2000 ;
	    RECT 243.0000 86.8000 243.4000 87.2000 ;
	    RECT 239.0000 86.2000 239.3000 86.8000 ;
	    RECT 239.0000 85.8000 239.4000 86.2000 ;
	    RECT 229.4000 83.8000 229.8000 84.2000 ;
	    RECT 229.4000 77.2000 229.7000 83.8000 ;
	    RECT 231.8000 79.2000 232.1000 84.8000 ;
	    RECT 232.7000 84.7000 233.1000 85.1000 ;
	    RECT 235.8000 84.7000 236.2000 85.1000 ;
	    RECT 234.2000 83.8000 234.6000 84.2000 ;
	    RECT 231.8000 78.8000 232.2000 79.2000 ;
	    RECT 222.2000 76.8000 222.6000 77.2000 ;
	    RECT 223.8000 76.8000 224.2000 77.2000 ;
	    RECT 229.4000 76.8000 229.8000 77.2000 ;
	    RECT 220.6000 72.8000 221.0000 73.2000 ;
	    RECT 220.6000 72.2000 220.9000 72.8000 ;
	    RECT 219.0000 72.1000 219.4000 72.2000 ;
	    RECT 219.8000 72.1000 220.2000 72.2000 ;
	    RECT 219.0000 71.8000 220.2000 72.1000 ;
	    RECT 220.6000 71.8000 221.0000 72.2000 ;
	    RECT 219.8000 69.8000 220.2000 70.2000 ;
	    RECT 219.8000 69.2000 220.1000 69.8000 ;
	    RECT 219.8000 68.8000 220.2000 69.2000 ;
	    RECT 219.8000 68.1000 220.2000 68.2000 ;
	    RECT 220.6000 68.1000 221.0000 68.2000 ;
	    RECT 219.8000 67.8000 221.0000 68.1000 ;
	    RECT 222.2000 67.2000 222.5000 76.8000 ;
	    RECT 227.8000 75.8000 228.2000 76.2000 ;
	    RECT 225.4000 75.1000 225.8000 75.2000 ;
	    RECT 226.2000 75.1000 226.6000 75.2000 ;
	    RECT 225.4000 74.8000 226.6000 75.1000 ;
	    RECT 227.0000 74.8000 227.4000 75.2000 ;
	    RECT 227.0000 74.2000 227.3000 74.8000 ;
	    RECT 223.0000 74.1000 223.4000 74.2000 ;
	    RECT 223.8000 74.1000 224.2000 74.2000 ;
	    RECT 223.0000 73.8000 224.2000 74.1000 ;
	    RECT 227.0000 73.8000 227.4000 74.2000 ;
	    RECT 223.8000 72.8000 224.2000 73.2000 ;
	    RECT 223.8000 71.2000 224.1000 72.8000 ;
	    RECT 223.8000 70.8000 224.2000 71.2000 ;
	    RECT 227.8000 69.2000 228.1000 75.8000 ;
	    RECT 229.4000 75.2000 229.7000 76.8000 ;
	    RECT 234.2000 76.2000 234.5000 83.8000 ;
	    RECT 240.6000 76.2000 240.9000 86.8000 ;
	    RECT 244.6000 86.1000 245.0000 86.2000 ;
	    RECT 245.4000 86.1000 245.8000 86.2000 ;
	    RECT 244.6000 85.8000 245.8000 86.1000 ;
	    RECT 242.2000 81.8000 242.6000 82.2000 ;
	    RECT 242.2000 79.2000 242.5000 81.8000 ;
	    RECT 242.2000 78.8000 242.6000 79.2000 ;
	    RECT 244.6000 78.2000 244.9000 85.8000 ;
	    RECT 245.4000 84.8000 245.8000 85.2000 ;
	    RECT 245.4000 84.2000 245.7000 84.8000 ;
	    RECT 245.4000 83.8000 245.8000 84.2000 ;
	    RECT 244.6000 77.8000 245.0000 78.2000 ;
	    RECT 247.8000 77.2000 248.1000 91.8000 ;
	    RECT 251.0000 91.2000 251.3000 106.8000 ;
	    RECT 251.8000 106.2000 252.1000 111.8000 ;
	    RECT 252.6000 109.2000 252.9000 112.8000 ;
	    RECT 264.6000 109.2000 264.9000 113.8000 ;
	    RECT 267.8000 111.8000 268.2000 112.2000 ;
	    RECT 252.6000 108.8000 253.0000 109.2000 ;
	    RECT 264.6000 108.8000 265.0000 109.2000 ;
	    RECT 267.8000 108.1000 268.1000 111.8000 ;
	    RECT 268.6000 108.1000 269.0000 108.2000 ;
	    RECT 256.7000 107.8000 257.1000 107.9000 ;
	    RECT 256.7000 107.5000 259.5000 107.8000 ;
	    RECT 259.8000 107.5000 260.2000 107.9000 ;
	    RECT 267.8000 107.8000 269.0000 108.1000 ;
	    RECT 252.6000 106.8000 253.0000 107.2000 ;
	    RECT 251.8000 105.8000 252.2000 106.2000 ;
	    RECT 252.6000 105.1000 252.9000 106.8000 ;
	    RECT 255.0000 106.1000 255.4000 106.2000 ;
	    RECT 255.8000 106.1000 256.2000 106.2000 ;
	    RECT 255.0000 105.8000 256.2000 106.1000 ;
	    RECT 251.8000 104.8000 252.9000 105.1000 ;
	    RECT 255.0000 104.8000 255.4000 105.2000 ;
	    RECT 256.7000 105.1000 257.0000 107.5000 ;
	    RECT 257.4000 107.4000 257.8000 107.5000 ;
	    RECT 259.1000 107.4000 259.5000 107.5000 ;
	    RECT 259.9000 107.1000 260.2000 107.5000 ;
	    RECT 257.4000 106.8000 260.2000 107.1000 ;
	    RECT 261.4000 107.1000 261.8000 107.2000 ;
	    RECT 262.2000 107.1000 262.6000 107.2000 ;
	    RECT 261.4000 106.8000 262.6000 107.1000 ;
	    RECT 266.2000 106.8000 266.6000 107.2000 ;
	    RECT 257.4000 106.1000 257.7000 106.8000 ;
	    RECT 257.3000 105.7000 257.7000 106.1000 ;
	    RECT 259.9000 105.1000 260.2000 106.8000 ;
	    RECT 266.2000 106.2000 266.5000 106.8000 ;
	    RECT 263.0000 105.8000 263.4000 106.2000 ;
	    RECT 264.6000 105.8000 265.0000 106.2000 ;
	    RECT 266.2000 105.8000 266.6000 106.2000 ;
	    RECT 251.8000 99.2000 252.1000 104.8000 ;
	    RECT 255.0000 104.2000 255.3000 104.8000 ;
	    RECT 256.7000 104.7000 257.1000 105.1000 ;
	    RECT 259.8000 104.7000 260.2000 105.1000 ;
	    RECT 260.6000 105.1000 261.0000 105.2000 ;
	    RECT 261.4000 105.1000 261.8000 105.2000 ;
	    RECT 260.6000 104.8000 261.8000 105.1000 ;
	    RECT 263.0000 104.2000 263.3000 105.8000 ;
	    RECT 264.6000 105.2000 264.9000 105.8000 ;
	    RECT 264.6000 104.8000 265.0000 105.2000 ;
	    RECT 255.0000 103.8000 255.4000 104.2000 ;
	    RECT 263.0000 103.8000 263.4000 104.2000 ;
	    RECT 267.0000 103.8000 267.4000 104.2000 ;
	    RECT 257.4000 102.1000 257.8000 102.2000 ;
	    RECT 258.2000 102.1000 258.6000 102.2000 ;
	    RECT 257.4000 101.8000 258.6000 102.1000 ;
	    RECT 251.8000 98.8000 252.2000 99.2000 ;
	    RECT 263.8000 97.1000 264.2000 97.2000 ;
	    RECT 264.6000 97.1000 265.0000 97.2000 ;
	    RECT 263.8000 96.8000 265.0000 97.1000 ;
	    RECT 257.5000 95.9000 257.9000 96.3000 ;
	    RECT 260.6000 95.9000 261.0000 96.3000 ;
	    RECT 253.4000 94.8000 253.8000 95.2000 ;
	    RECT 251.0000 90.8000 251.4000 91.2000 ;
	    RECT 251.0000 88.8000 251.4000 89.2000 ;
	    RECT 251.0000 88.2000 251.3000 88.8000 ;
	    RECT 251.0000 87.8000 251.4000 88.2000 ;
	    RECT 253.4000 87.2000 253.7000 94.8000 ;
	    RECT 257.5000 93.5000 257.8000 95.9000 ;
	    RECT 258.1000 94.9000 258.5000 95.3000 ;
	    RECT 258.2000 94.2000 258.5000 94.9000 ;
	    RECT 260.7000 94.2000 261.0000 95.9000 ;
	    RECT 258.2000 93.9000 261.0000 94.2000 ;
	    RECT 258.2000 93.5000 258.6000 93.6000 ;
	    RECT 259.9000 93.5000 260.3000 93.6000 ;
	    RECT 260.7000 93.5000 261.0000 93.9000 ;
	    RECT 257.5000 93.2000 260.3000 93.5000 ;
	    RECT 254.2000 93.1000 254.6000 93.2000 ;
	    RECT 255.0000 93.1000 255.4000 93.2000 ;
	    RECT 257.5000 93.1000 257.9000 93.2000 ;
	    RECT 260.6000 93.1000 261.0000 93.5000 ;
	    RECT 263.0000 95.9000 263.4000 96.3000 ;
	    RECT 266.3000 95.9000 266.7000 96.3000 ;
	    RECT 263.0000 94.2000 263.3000 95.9000 ;
	    RECT 265.0000 94.2000 265.4000 94.3000 ;
	    RECT 263.0000 93.9000 265.4000 94.2000 ;
	    RECT 263.0000 93.5000 263.3000 93.9000 ;
	    RECT 263.7000 93.5000 264.1000 93.6000 ;
	    RECT 265.4000 93.5000 265.8000 93.6000 ;
	    RECT 266.4000 93.5000 266.7000 95.9000 ;
	    RECT 263.0000 93.1000 263.4000 93.5000 ;
	    RECT 263.7000 93.2000 265.8000 93.5000 ;
	    RECT 266.3000 93.1000 266.7000 93.5000 ;
	    RECT 267.0000 94.2000 267.3000 103.8000 ;
	    RECT 267.0000 93.8000 267.4000 94.2000 ;
	    RECT 254.2000 92.8000 255.4000 93.1000 ;
	    RECT 258.2000 92.1000 258.6000 92.2000 ;
	    RECT 259.0000 92.1000 259.4000 92.2000 ;
	    RECT 258.2000 91.8000 259.4000 92.1000 ;
	    RECT 265.4000 90.8000 265.8000 91.2000 ;
	    RECT 265.4000 89.2000 265.7000 90.8000 ;
	    RECT 259.8000 89.1000 260.2000 89.2000 ;
	    RECT 260.6000 89.1000 261.0000 89.2000 ;
	    RECT 259.8000 88.8000 261.0000 89.1000 ;
	    RECT 265.4000 88.8000 265.8000 89.2000 ;
	    RECT 259.1000 87.8000 259.5000 87.9000 ;
	    RECT 259.1000 87.5000 261.9000 87.8000 ;
	    RECT 262.2000 87.5000 262.6000 87.9000 ;
	    RECT 253.4000 86.8000 253.8000 87.2000 ;
	    RECT 255.0000 87.1000 255.4000 87.2000 ;
	    RECT 255.8000 87.1000 256.2000 87.2000 ;
	    RECT 255.0000 86.8000 256.2000 87.1000 ;
	    RECT 252.6000 86.1000 253.0000 86.2000 ;
	    RECT 253.4000 86.1000 253.8000 86.2000 ;
	    RECT 252.6000 85.8000 253.8000 86.1000 ;
	    RECT 255.8000 85.8000 256.2000 86.2000 ;
	    RECT 256.6000 86.1000 257.0000 86.2000 ;
	    RECT 257.4000 86.1000 257.8000 86.2000 ;
	    RECT 256.6000 85.8000 257.8000 86.1000 ;
	    RECT 248.6000 84.8000 249.0000 85.2000 ;
	    RECT 251.8000 84.8000 252.2000 85.2000 ;
	    RECT 254.2000 84.8000 254.6000 85.2000 ;
	    RECT 248.6000 80.2000 248.9000 84.8000 ;
	    RECT 248.6000 79.8000 249.0000 80.2000 ;
	    RECT 251.8000 79.2000 252.1000 84.8000 ;
	    RECT 254.2000 83.2000 254.5000 84.8000 ;
	    RECT 254.2000 82.8000 254.6000 83.2000 ;
	    RECT 251.8000 78.8000 252.2000 79.2000 ;
	    RECT 252.6000 78.8000 253.0000 79.2000 ;
	    RECT 252.6000 77.2000 252.9000 78.8000 ;
	    RECT 247.8000 76.8000 248.2000 77.2000 ;
	    RECT 252.6000 76.8000 253.0000 77.2000 ;
	    RECT 234.2000 75.8000 234.6000 76.2000 ;
	    RECT 238.2000 75.8000 238.6000 76.2000 ;
	    RECT 240.6000 75.8000 241.0000 76.2000 ;
	    RECT 243.0000 76.1000 243.4000 76.2000 ;
	    RECT 243.8000 76.1000 244.2000 76.2000 ;
	    RECT 243.0000 75.8000 244.2000 76.1000 ;
	    RECT 247.1000 75.9000 247.5000 76.3000 ;
	    RECT 250.2000 75.9000 250.6000 76.3000 ;
	    RECT 234.2000 75.2000 234.5000 75.8000 ;
	    RECT 228.6000 74.8000 229.0000 75.2000 ;
	    RECT 229.4000 74.8000 229.8000 75.2000 ;
	    RECT 231.8000 75.1000 232.2000 75.2000 ;
	    RECT 232.6000 75.1000 233.0000 75.2000 ;
	    RECT 231.8000 74.8000 233.0000 75.1000 ;
	    RECT 234.2000 74.8000 234.6000 75.2000 ;
	    RECT 236.6000 74.8000 237.0000 75.2000 ;
	    RECT 228.6000 71.2000 228.9000 74.8000 ;
	    RECT 236.6000 74.2000 236.9000 74.8000 ;
	    RECT 230.2000 74.1000 230.6000 74.2000 ;
	    RECT 231.0000 74.1000 231.4000 74.2000 ;
	    RECT 230.2000 73.8000 231.4000 74.1000 ;
	    RECT 236.6000 73.8000 237.0000 74.2000 ;
	    RECT 237.4000 73.8000 237.8000 74.2000 ;
	    RECT 238.2000 74.1000 238.5000 75.8000 ;
	    RECT 239.0000 75.1000 239.4000 75.2000 ;
	    RECT 239.8000 75.1000 240.2000 75.2000 ;
	    RECT 239.0000 74.8000 240.2000 75.1000 ;
	    RECT 240.6000 74.8000 241.0000 75.2000 ;
	    RECT 240.6000 74.2000 240.9000 74.8000 ;
	    RECT 239.0000 74.1000 239.4000 74.2000 ;
	    RECT 238.2000 73.8000 239.4000 74.1000 ;
	    RECT 239.8000 73.8000 240.2000 74.2000 ;
	    RECT 240.6000 73.8000 241.0000 74.2000 ;
	    RECT 237.4000 73.2000 237.7000 73.8000 ;
	    RECT 237.4000 72.8000 237.8000 73.2000 ;
	    RECT 229.4000 71.8000 229.8000 72.2000 ;
	    RECT 239.0000 71.8000 239.4000 72.2000 ;
	    RECT 228.6000 70.8000 229.0000 71.2000 ;
	    RECT 229.4000 69.2000 229.7000 71.8000 ;
	    RECT 234.2000 70.8000 234.6000 71.2000 ;
	    RECT 234.2000 69.2000 234.5000 70.8000 ;
	    RECT 237.4000 69.8000 237.8000 70.2000 ;
	    RECT 224.6000 68.8000 225.0000 69.2000 ;
	    RECT 227.0000 68.8000 227.4000 69.2000 ;
	    RECT 227.8000 68.8000 228.2000 69.2000 ;
	    RECT 229.4000 68.8000 229.8000 69.2000 ;
	    RECT 232.6000 68.8000 233.0000 69.2000 ;
	    RECT 234.2000 68.8000 234.6000 69.2000 ;
	    RECT 214.2000 66.8000 214.6000 67.2000 ;
	    RECT 218.2000 66.8000 218.6000 67.2000 ;
	    RECT 222.2000 66.8000 222.6000 67.2000 ;
	    RECT 223.0000 67.1000 223.4000 67.2000 ;
	    RECT 223.8000 67.1000 224.2000 67.2000 ;
	    RECT 223.0000 66.8000 224.2000 67.1000 ;
	    RECT 210.2000 66.1000 210.6000 66.2000 ;
	    RECT 209.4000 65.8000 210.6000 66.1000 ;
	    RECT 211.8000 66.1000 212.2000 66.2000 ;
	    RECT 212.6000 66.1000 213.0000 66.2000 ;
	    RECT 211.8000 65.8000 213.0000 66.1000 ;
	    RECT 213.4000 66.1000 213.8000 66.2000 ;
	    RECT 214.2000 66.1000 214.6000 66.2000 ;
	    RECT 213.4000 65.8000 214.6000 66.1000 ;
	    RECT 215.8000 66.1000 216.2000 66.2000 ;
	    RECT 216.6000 66.1000 217.0000 66.2000 ;
	    RECT 215.8000 65.8000 217.0000 66.1000 ;
	    RECT 195.0000 64.7000 195.4000 65.1000 ;
	    RECT 198.3000 64.7000 198.7000 65.1000 ;
	    RECT 218.2000 65.2000 218.5000 66.8000 ;
	    RECT 224.6000 66.2000 224.9000 68.8000 ;
	    RECT 227.0000 67.2000 227.3000 68.8000 ;
	    RECT 232.6000 68.2000 232.9000 68.8000 ;
	    RECT 232.6000 67.8000 233.0000 68.2000 ;
	    RECT 237.4000 67.2000 237.7000 69.8000 ;
	    RECT 227.0000 66.8000 227.4000 67.2000 ;
	    RECT 232.6000 67.1000 233.0000 67.2000 ;
	    RECT 233.4000 67.1000 233.8000 67.2000 ;
	    RECT 232.6000 66.8000 233.8000 67.1000 ;
	    RECT 235.8000 67.1000 236.2000 67.2000 ;
	    RECT 236.6000 67.1000 237.0000 67.2000 ;
	    RECT 235.8000 66.8000 237.0000 67.1000 ;
	    RECT 237.4000 66.8000 237.8000 67.2000 ;
	    RECT 219.8000 65.8000 220.2000 66.2000 ;
	    RECT 221.4000 65.8000 221.8000 66.2000 ;
	    RECT 223.8000 65.8000 224.2000 66.2000 ;
	    RECT 224.6000 65.8000 225.0000 66.2000 ;
	    RECT 219.8000 65.2000 220.1000 65.8000 ;
	    RECT 218.2000 64.8000 218.6000 65.2000 ;
	    RECT 219.8000 64.8000 220.2000 65.2000 ;
	    RECT 211.0000 64.1000 211.4000 64.2000 ;
	    RECT 211.8000 64.1000 212.2000 64.2000 ;
	    RECT 211.0000 63.8000 212.2000 64.1000 ;
	    RECT 215.0000 64.1000 215.4000 64.2000 ;
	    RECT 215.8000 64.1000 216.2000 64.2000 ;
	    RECT 215.0000 63.8000 216.2000 64.1000 ;
	    RECT 216.6000 61.8000 217.0000 62.2000 ;
	    RECT 192.6000 58.8000 193.0000 59.2000 ;
	    RECT 193.4000 58.8000 193.8000 59.2000 ;
	    RECT 194.2000 58.8000 194.6000 59.2000 ;
	    RECT 191.0000 56.8000 191.4000 57.2000 ;
	    RECT 197.4000 52.1000 197.8000 57.9000 ;
	    RECT 198.2000 54.8000 198.6000 55.2000 ;
	    RECT 198.2000 51.2000 198.5000 54.8000 ;
	    RECT 202.2000 52.1000 202.6000 57.9000 ;
	    RECT 203.8000 53.1000 204.2000 55.9000 ;
	    RECT 206.2000 54.8000 206.6000 55.2000 ;
	    RECT 207.0000 54.8000 207.4000 55.2000 ;
	    RECT 206.2000 54.2000 206.5000 54.8000 ;
	    RECT 204.6000 54.1000 205.0000 54.2000 ;
	    RECT 205.4000 54.1000 205.8000 54.2000 ;
	    RECT 204.6000 53.8000 205.8000 54.1000 ;
	    RECT 206.2000 53.8000 206.6000 54.2000 ;
	    RECT 204.6000 52.8000 205.0000 53.2000 ;
	    RECT 205.4000 52.8000 205.8000 53.2000 ;
	    RECT 187.8000 50.8000 188.2000 51.2000 ;
	    RECT 189.4000 50.8000 189.8000 51.2000 ;
	    RECT 195.8000 50.8000 196.2000 51.2000 ;
	    RECT 198.2000 50.8000 198.6000 51.2000 ;
	    RECT 199.8000 50.8000 200.2000 51.2000 ;
	    RECT 183.0000 46.8000 183.4000 47.2000 ;
	    RECT 181.4000 45.8000 181.8000 46.2000 ;
	    RECT 184.6000 43.1000 185.0000 48.9000 ;
	    RECT 186.2000 45.1000 186.6000 47.9000 ;
	    RECT 187.0000 47.8000 187.4000 48.2000 ;
	    RECT 187.0000 47.2000 187.3000 47.8000 ;
	    RECT 187.0000 46.8000 187.4000 47.2000 ;
	    RECT 187.8000 46.2000 188.1000 50.8000 ;
	    RECT 187.8000 45.8000 188.2000 46.2000 ;
	    RECT 189.4000 45.8000 189.8000 46.2000 ;
	    RECT 189.4000 45.2000 189.7000 45.8000 ;
	    RECT 189.4000 44.8000 189.8000 45.2000 ;
	    RECT 190.2000 45.1000 190.6000 47.9000 ;
	    RECT 191.8000 43.1000 192.2000 48.9000 ;
	    RECT 194.2000 47.8000 194.6000 48.2000 ;
	    RECT 192.6000 45.9000 193.0000 46.3000 ;
	    RECT 192.6000 45.2000 192.9000 45.9000 ;
	    RECT 192.6000 44.8000 193.0000 45.2000 ;
	    RECT 175.8000 41.8000 176.2000 42.2000 ;
	    RECT 174.2000 38.8000 174.6000 39.2000 ;
	    RECT 168.6000 33.8000 169.0000 34.2000 ;
	    RECT 169.4000 33.1000 169.8000 35.9000 ;
	    RECT 173.4000 35.8000 173.8000 36.2000 ;
	    RECT 173.4000 35.2000 173.7000 35.8000 ;
	    RECT 175.8000 35.2000 176.1000 41.8000 ;
	    RECT 171.8000 34.8000 172.2000 35.2000 ;
	    RECT 173.4000 35.1000 173.8000 35.2000 ;
	    RECT 174.2000 35.1000 174.6000 35.2000 ;
	    RECT 173.4000 34.8000 174.6000 35.1000 ;
	    RECT 175.8000 34.8000 176.2000 35.2000 ;
	    RECT 177.4000 34.8000 177.8000 35.2000 ;
	    RECT 171.8000 34.2000 172.1000 34.8000 ;
	    RECT 177.4000 34.2000 177.7000 34.8000 ;
	    RECT 171.8000 33.8000 172.2000 34.2000 ;
	    RECT 177.4000 33.8000 177.8000 34.2000 ;
	    RECT 170.2000 32.8000 170.6000 33.2000 ;
	    RECT 175.0000 32.8000 175.4000 33.2000 ;
	    RECT 177.4000 32.8000 177.8000 33.2000 ;
	    RECT 179.0000 33.1000 179.4000 35.9000 ;
	    RECT 179.8000 34.8000 180.2000 35.2000 ;
	    RECT 179.8000 34.2000 180.1000 34.8000 ;
	    RECT 179.8000 33.8000 180.2000 34.2000 ;
	    RECT 170.2000 32.2000 170.5000 32.8000 ;
	    RECT 160.6000 31.8000 161.8000 32.1000 ;
	    RECT 170.2000 31.8000 170.6000 32.2000 ;
	    RECT 156.6000 25.2000 156.9000 25.9000 ;
	    RECT 159.0000 25.8000 159.4000 26.2000 ;
	    RECT 156.6000 24.8000 157.0000 25.2000 ;
	    RECT 143.0000 21.8000 143.4000 22.2000 ;
	    RECT 131.0000 15.8000 131.4000 16.2000 ;
	    RECT 131.0000 15.1000 131.3000 15.8000 ;
	    RECT 131.0000 14.7000 131.4000 15.1000 ;
	    RECT 130.2000 13.8000 130.6000 14.2000 ;
	    RECT 131.8000 12.1000 132.2000 17.9000 ;
	    RECT 136.6000 16.1000 137.0000 16.2000 ;
	    RECT 137.4000 16.1000 137.8000 16.2000 ;
	    RECT 133.4000 13.1000 133.8000 15.9000 ;
	    RECT 136.6000 15.8000 137.8000 16.1000 ;
	    RECT 139.0000 15.9000 139.4000 16.3000 ;
	    RECT 142.3000 15.9000 142.7000 16.3000 ;
	    RECT 137.4000 14.8000 137.8000 15.2000 ;
	    RECT 138.2000 14.8000 138.6000 15.2000 ;
	    RECT 137.4000 14.2000 137.7000 14.8000 ;
	    RECT 138.2000 14.2000 138.5000 14.8000 ;
	    RECT 139.0000 14.2000 139.3000 15.9000 ;
	    RECT 141.0000 14.2000 141.4000 14.3000 ;
	    RECT 137.4000 13.8000 137.8000 14.2000 ;
	    RECT 138.2000 13.8000 138.6000 14.2000 ;
	    RECT 139.0000 13.9000 141.4000 14.2000 ;
	    RECT 139.0000 13.5000 139.3000 13.9000 ;
	    RECT 139.7000 13.5000 140.1000 13.6000 ;
	    RECT 141.4000 13.5000 141.8000 13.6000 ;
	    RECT 142.4000 13.5000 142.7000 15.9000 ;
	    RECT 143.0000 14.2000 143.3000 21.8000 ;
	    RECT 157.4000 15.8000 157.8000 16.2000 ;
	    RECT 157.4000 15.2000 157.7000 15.8000 ;
	    RECT 147.0000 15.1000 147.4000 15.2000 ;
	    RECT 147.8000 15.1000 148.2000 15.2000 ;
	    RECT 147.0000 14.8000 148.2000 15.1000 ;
	    RECT 155.0000 14.8000 155.4000 15.2000 ;
	    RECT 157.4000 14.8000 157.8000 15.2000 ;
	    RECT 147.0000 14.2000 147.3000 14.8000 ;
	    RECT 155.0000 14.2000 155.3000 14.8000 ;
	    RECT 143.0000 13.8000 143.4000 14.2000 ;
	    RECT 147.0000 13.8000 147.4000 14.2000 ;
	    RECT 155.0000 13.8000 155.4000 14.2000 ;
	    RECT 134.2000 12.8000 134.6000 13.2000 ;
	    RECT 136.6000 12.8000 137.0000 13.2000 ;
	    RECT 139.0000 13.1000 139.4000 13.5000 ;
	    RECT 139.7000 13.2000 141.8000 13.5000 ;
	    RECT 142.3000 13.1000 142.7000 13.5000 ;
	    RECT 155.0000 13.2000 155.3000 13.8000 ;
	    RECT 143.8000 12.8000 144.2000 13.2000 ;
	    RECT 147.0000 12.8000 147.4000 13.2000 ;
	    RECT 155.0000 12.8000 155.4000 13.2000 ;
	    RECT 158.2000 12.8000 158.6000 13.2000 ;
	    RECT 124.6000 11.8000 125.7000 12.1000 ;
	    RECT 124.6000 9.8000 125.0000 10.2000 ;
	    RECT 115.8000 8.8000 116.2000 9.2000 ;
	    RECT 117.4000 8.8000 117.8000 9.2000 ;
	    RECT 123.0000 8.8000 123.4000 9.2000 ;
	    RECT 112.5000 7.5000 114.6000 7.8000 ;
	    RECT 115.1000 7.5000 115.5000 7.9000 ;
	    RECT 104.6000 7.1000 105.0000 7.2000 ;
	    RECT 103.8000 6.8000 105.0000 7.1000 ;
	    RECT 105.4000 6.8000 105.8000 7.2000 ;
	    RECT 111.0000 6.8000 111.4000 7.2000 ;
	    RECT 111.8000 7.1000 112.1000 7.5000 ;
	    RECT 112.5000 7.4000 112.9000 7.5000 ;
	    RECT 114.2000 7.4000 114.6000 7.5000 ;
	    RECT 111.8000 6.8000 114.2000 7.1000 ;
	    RECT 96.6000 6.2000 96.9000 6.8000 ;
	    RECT 99.8000 6.2000 100.1000 6.8000 ;
	    RECT 105.4000 6.2000 105.7000 6.8000 ;
	    RECT 96.6000 5.8000 97.0000 6.2000 ;
	    RECT 99.8000 5.8000 100.2000 6.2000 ;
	    RECT 100.6000 6.1000 101.0000 6.2000 ;
	    RECT 101.4000 6.1000 101.8000 6.2000 ;
	    RECT 100.6000 5.8000 101.8000 6.1000 ;
	    RECT 103.0000 5.8000 103.4000 6.2000 ;
	    RECT 105.4000 5.8000 105.8000 6.2000 ;
	    RECT 103.0000 5.2000 103.3000 5.8000 ;
	    RECT 83.0000 4.8000 83.4000 5.2000 ;
	    RECT 86.2000 4.8000 86.6000 5.2000 ;
	    RECT 87.0000 4.8000 87.4000 5.2000 ;
	    RECT 89.4000 4.8000 89.8000 5.2000 ;
	    RECT 93.4000 4.8000 93.8000 5.2000 ;
	    RECT 95.8000 4.8000 96.2000 5.2000 ;
	    RECT 103.0000 4.8000 103.4000 5.2000 ;
	    RECT 111.8000 5.1000 112.1000 6.8000 ;
	    RECT 113.8000 6.7000 114.2000 6.8000 ;
	    RECT 112.6000 5.1000 113.0000 5.2000 ;
	    RECT 113.4000 5.1000 113.8000 5.2000 ;
	    RECT 115.2000 5.1000 115.5000 7.5000 ;
	    RECT 115.8000 7.2000 116.1000 8.8000 ;
	    RECT 116.6000 7.8000 117.0000 8.2000 ;
	    RECT 120.6000 7.8000 121.0000 8.2000 ;
	    RECT 121.4000 8.1000 121.8000 8.2000 ;
	    RECT 122.2000 8.1000 122.6000 8.2000 ;
	    RECT 121.4000 7.8000 122.6000 8.1000 ;
	    RECT 123.0000 7.8000 123.4000 8.2000 ;
	    RECT 115.8000 6.8000 116.2000 7.2000 ;
	    RECT 111.8000 4.7000 112.2000 5.1000 ;
	    RECT 112.6000 4.8000 113.8000 5.1000 ;
	    RECT 115.1000 4.7000 115.5000 5.1000 ;
	    RECT 116.6000 5.2000 116.9000 7.8000 ;
	    RECT 118.2000 6.8000 118.6000 7.2000 ;
	    RECT 118.2000 6.2000 118.5000 6.8000 ;
	    RECT 120.6000 6.2000 120.9000 7.8000 ;
	    RECT 117.4000 5.8000 117.8000 6.2000 ;
	    RECT 118.2000 5.8000 118.6000 6.2000 ;
	    RECT 120.6000 5.8000 121.0000 6.2000 ;
	    RECT 122.2000 5.8000 122.6000 6.2000 ;
	    RECT 116.6000 4.8000 117.0000 5.2000 ;
	    RECT 117.4000 5.1000 117.7000 5.8000 ;
	    RECT 122.2000 5.2000 122.5000 5.8000 ;
	    RECT 123.0000 5.2000 123.3000 7.8000 ;
	    RECT 124.6000 7.2000 124.9000 9.8000 ;
	    RECT 125.4000 9.2000 125.7000 11.8000 ;
	    RECT 132.6000 11.8000 133.0000 12.2000 ;
	    RECT 132.6000 9.2000 132.9000 11.8000 ;
	    RECT 134.2000 9.2000 134.5000 12.8000 ;
	    RECT 125.4000 8.8000 125.8000 9.2000 ;
	    RECT 130.2000 8.8000 130.6000 9.2000 ;
	    RECT 132.6000 8.8000 133.0000 9.2000 ;
	    RECT 134.2000 8.8000 134.6000 9.2000 ;
	    RECT 125.4000 7.8000 125.8000 8.2000 ;
	    RECT 125.4000 7.2000 125.7000 7.8000 ;
	    RECT 126.2000 7.5000 126.6000 7.9000 ;
	    RECT 129.3000 7.8000 129.7000 7.9000 ;
	    RECT 126.9000 7.5000 129.7000 7.8000 ;
	    RECT 124.6000 6.8000 125.0000 7.2000 ;
	    RECT 125.4000 6.8000 125.8000 7.2000 ;
	    RECT 126.2000 7.1000 126.5000 7.5000 ;
	    RECT 126.9000 7.4000 127.3000 7.5000 ;
	    RECT 128.6000 7.4000 129.0000 7.5000 ;
	    RECT 126.2000 6.8000 129.0000 7.1000 ;
	    RECT 118.2000 5.1000 118.6000 5.2000 ;
	    RECT 117.4000 4.8000 118.6000 5.1000 ;
	    RECT 122.2000 4.8000 122.6000 5.2000 ;
	    RECT 123.0000 4.8000 123.4000 5.2000 ;
	    RECT 126.2000 5.1000 126.5000 6.8000 ;
	    RECT 127.0000 5.8000 127.4000 6.2000 ;
	    RECT 128.7000 6.1000 129.0000 6.8000 ;
	    RECT 127.0000 5.2000 127.3000 5.8000 ;
	    RECT 128.7000 5.7000 129.1000 6.1000 ;
	    RECT 126.2000 4.7000 126.6000 5.1000 ;
	    RECT 127.0000 4.8000 127.4000 5.2000 ;
	    RECT 129.4000 5.1000 129.7000 7.5000 ;
	    RECT 130.2000 7.2000 130.5000 8.8000 ;
	    RECT 136.6000 8.2000 136.9000 12.8000 ;
	    RECT 140.6000 11.8000 141.0000 12.2000 ;
	    RECT 141.4000 11.8000 141.8000 12.2000 ;
	    RECT 139.8000 8.8000 140.2000 9.2000 ;
	    RECT 139.8000 8.2000 140.1000 8.8000 ;
	    RECT 131.8000 7.8000 132.2000 8.2000 ;
	    RECT 134.2000 8.1000 134.6000 8.2000 ;
	    RECT 135.0000 8.1000 135.4000 8.2000 ;
	    RECT 134.2000 7.8000 135.4000 8.1000 ;
	    RECT 136.6000 7.8000 137.0000 8.2000 ;
	    RECT 139.8000 7.8000 140.2000 8.2000 ;
	    RECT 131.8000 7.2000 132.1000 7.8000 ;
	    RECT 136.6000 7.2000 136.9000 7.8000 ;
	    RECT 130.2000 6.8000 130.6000 7.2000 ;
	    RECT 131.0000 6.8000 131.4000 7.2000 ;
	    RECT 131.8000 6.8000 132.2000 7.2000 ;
	    RECT 136.6000 6.8000 137.0000 7.2000 ;
	    RECT 137.4000 7.1000 137.8000 7.2000 ;
	    RECT 138.2000 7.1000 138.6000 7.2000 ;
	    RECT 137.4000 6.8000 138.6000 7.1000 ;
	    RECT 131.0000 6.2000 131.3000 6.8000 ;
	    RECT 131.0000 5.8000 131.4000 6.2000 ;
	    RECT 135.8000 5.8000 136.2000 6.2000 ;
	    RECT 138.2000 5.8000 138.6000 6.2000 ;
	    RECT 129.3000 4.7000 129.7000 5.1000 ;
	    RECT 135.8000 5.2000 136.1000 5.8000 ;
	    RECT 138.2000 5.2000 138.5000 5.8000 ;
	    RECT 140.6000 5.2000 140.9000 11.8000 ;
	    RECT 141.4000 9.2000 141.7000 11.8000 ;
	    RECT 143.8000 11.2000 144.1000 12.8000 ;
	    RECT 143.8000 10.8000 144.2000 11.2000 ;
	    RECT 141.4000 8.8000 141.8000 9.2000 ;
	    RECT 143.0000 9.1000 143.4000 9.2000 ;
	    RECT 143.8000 9.1000 144.1000 10.8000 ;
	    RECT 143.0000 8.8000 144.1000 9.1000 ;
	    RECT 142.2000 6.8000 142.6000 7.2000 ;
	    RECT 142.2000 5.2000 142.5000 6.8000 ;
	    RECT 135.8000 4.8000 136.2000 5.2000 ;
	    RECT 138.2000 4.8000 138.6000 5.2000 ;
	    RECT 140.6000 4.8000 141.0000 5.2000 ;
	    RECT 142.2000 4.8000 142.6000 5.2000 ;
	    RECT 145.4000 3.1000 145.8000 8.9000 ;
	    RECT 147.0000 6.2000 147.3000 12.8000 ;
	    RECT 153.4000 11.8000 153.8000 12.2000 ;
	    RECT 153.4000 10.2000 153.7000 11.8000 ;
	    RECT 151.0000 9.8000 151.4000 10.2000 ;
	    RECT 153.4000 9.8000 153.8000 10.2000 ;
	    RECT 147.0000 5.8000 147.4000 6.2000 ;
	    RECT 150.2000 3.1000 150.6000 8.9000 ;
	    RECT 151.0000 7.2000 151.3000 9.8000 ;
	    RECT 158.2000 9.2000 158.5000 12.8000 ;
	    RECT 159.0000 10.2000 159.3000 25.8000 ;
	    RECT 160.6000 23.1000 161.0000 28.9000 ;
	    RECT 161.4000 22.2000 161.7000 31.8000 ;
	    RECT 175.0000 30.2000 175.3000 32.8000 ;
	    RECT 163.0000 29.8000 163.4000 30.2000 ;
	    RECT 166.2000 29.8000 166.6000 30.2000 ;
	    RECT 175.0000 29.8000 175.4000 30.2000 ;
	    RECT 163.0000 29.2000 163.3000 29.8000 ;
	    RECT 163.0000 28.8000 163.4000 29.2000 ;
	    RECT 165.4000 27.8000 165.8000 28.2000 ;
	    RECT 165.4000 27.2000 165.7000 27.8000 ;
	    RECT 165.4000 26.8000 165.8000 27.2000 ;
	    RECT 166.2000 26.2000 166.5000 29.8000 ;
	    RECT 177.4000 29.2000 177.7000 32.8000 ;
	    RECT 180.6000 32.1000 181.0000 37.9000 ;
	    RECT 181.4000 35.8000 181.8000 36.2000 ;
	    RECT 181.4000 35.1000 181.7000 35.8000 ;
	    RECT 181.4000 34.7000 181.8000 35.1000 ;
	    RECT 185.4000 32.1000 185.8000 37.9000 ;
	    RECT 187.8000 36.8000 188.2000 37.2000 ;
	    RECT 187.8000 36.2000 188.1000 36.8000 ;
	    RECT 194.2000 36.2000 194.5000 47.8000 ;
	    RECT 195.8000 46.2000 196.1000 50.8000 ;
	    RECT 199.8000 49.2000 200.1000 50.8000 ;
	    RECT 195.8000 45.8000 196.2000 46.2000 ;
	    RECT 187.8000 35.8000 188.2000 36.2000 ;
	    RECT 189.4000 35.8000 189.8000 36.2000 ;
	    RECT 191.8000 35.8000 192.2000 36.2000 ;
	    RECT 194.2000 35.8000 194.6000 36.2000 ;
	    RECT 188.6000 34.8000 189.0000 35.2000 ;
	    RECT 188.6000 34.2000 188.9000 34.8000 ;
	    RECT 189.4000 34.2000 189.7000 35.8000 ;
	    RECT 191.8000 35.2000 192.1000 35.8000 ;
	    RECT 191.8000 34.8000 192.2000 35.2000 ;
	    RECT 188.6000 33.8000 189.0000 34.2000 ;
	    RECT 189.4000 33.8000 189.8000 34.2000 ;
	    RECT 191.0000 34.1000 191.4000 34.2000 ;
	    RECT 191.8000 34.1000 192.2000 34.2000 ;
	    RECT 191.0000 33.8000 192.2000 34.1000 ;
	    RECT 193.4000 33.8000 193.8000 34.2000 ;
	    RECT 193.4000 33.2000 193.7000 33.8000 ;
	    RECT 191.0000 33.1000 191.4000 33.2000 ;
	    RECT 191.8000 33.1000 192.2000 33.2000 ;
	    RECT 191.0000 32.8000 192.2000 33.1000 ;
	    RECT 193.4000 32.8000 193.8000 33.2000 ;
	    RECT 190.2000 31.8000 190.6000 32.2000 ;
	    RECT 186.2000 30.8000 186.6000 31.2000 ;
	    RECT 178.2000 29.8000 178.6000 30.2000 ;
	    RECT 167.8000 28.8000 168.2000 29.2000 ;
	    RECT 167.8000 28.2000 168.1000 28.8000 ;
	    RECT 167.8000 27.8000 168.2000 28.2000 ;
	    RECT 166.2000 25.8000 166.6000 26.2000 ;
	    RECT 167.0000 25.1000 167.4000 25.2000 ;
	    RECT 167.8000 25.1000 168.2000 25.2000 ;
	    RECT 168.6000 25.1000 169.0000 27.9000 ;
	    RECT 169.4000 26.8000 169.8000 27.2000 ;
	    RECT 167.0000 24.8000 168.2000 25.1000 ;
	    RECT 161.4000 21.8000 161.8000 22.2000 ;
	    RECT 169.4000 19.2000 169.7000 26.8000 ;
	    RECT 170.2000 23.1000 170.6000 28.9000 ;
	    RECT 171.8000 26.8000 172.2000 27.2000 ;
	    RECT 171.8000 26.2000 172.1000 26.8000 ;
	    RECT 171.8000 25.8000 172.2000 26.2000 ;
	    RECT 175.0000 23.1000 175.4000 28.9000 ;
	    RECT 177.4000 28.8000 177.8000 29.2000 ;
	    RECT 178.2000 28.2000 178.5000 29.8000 ;
	    RECT 178.2000 27.8000 178.6000 28.2000 ;
	    RECT 181.4000 28.1000 181.8000 28.2000 ;
	    RECT 182.2000 28.1000 182.6000 28.2000 ;
	    RECT 181.4000 27.8000 182.6000 28.1000 ;
	    RECT 181.4000 25.2000 181.7000 27.8000 ;
	    RECT 181.4000 24.8000 181.8000 25.2000 ;
	    RECT 179.0000 24.1000 179.4000 24.2000 ;
	    RECT 179.8000 24.1000 180.2000 24.2000 ;
	    RECT 179.0000 23.8000 180.2000 24.1000 ;
	    RECT 169.4000 18.8000 169.8000 19.2000 ;
	    RECT 169.4000 16.2000 169.7000 18.8000 ;
	    RECT 173.4000 16.8000 173.8000 17.2000 ;
	    RECT 169.4000 15.8000 169.8000 16.2000 ;
	    RECT 173.4000 15.2000 173.7000 16.8000 ;
	    RECT 163.0000 15.1000 163.4000 15.2000 ;
	    RECT 162.2000 14.8000 163.4000 15.1000 ;
	    RECT 172.6000 15.1000 173.0000 15.2000 ;
	    RECT 173.4000 15.1000 173.8000 15.2000 ;
	    RECT 172.6000 14.8000 173.8000 15.1000 ;
	    RECT 162.2000 13.2000 162.5000 14.8000 ;
	    RECT 162.2000 12.8000 162.6000 13.2000 ;
	    RECT 163.0000 12.8000 163.4000 13.2000 ;
	    RECT 169.4000 12.8000 169.8000 13.2000 ;
	    RECT 159.0000 9.8000 159.4000 10.2000 ;
	    RECT 154.2000 8.8000 154.6000 9.2000 ;
	    RECT 158.2000 8.8000 158.6000 9.2000 ;
	    RECT 151.0000 6.8000 151.4000 7.2000 ;
	    RECT 151.8000 5.1000 152.2000 7.9000 ;
	    RECT 152.6000 7.8000 153.0000 8.2000 ;
	    RECT 152.6000 7.2000 152.9000 7.8000 ;
	    RECT 153.4000 7.5000 153.8000 7.9000 ;
	    RECT 154.2000 7.8000 154.5000 8.8000 ;
	    RECT 154.1000 7.5000 156.2000 7.8000 ;
	    RECT 156.7000 7.5000 157.1000 7.9000 ;
	    RECT 152.6000 6.8000 153.0000 7.2000 ;
	    RECT 153.4000 7.1000 153.7000 7.5000 ;
	    RECT 154.1000 7.4000 154.5000 7.5000 ;
	    RECT 155.8000 7.4000 156.2000 7.5000 ;
	    RECT 153.4000 6.8000 155.8000 7.1000 ;
	    RECT 153.4000 5.1000 153.7000 6.8000 ;
	    RECT 155.4000 6.7000 155.8000 6.8000 ;
	    RECT 153.4000 4.7000 153.8000 5.1000 ;
	    RECT 154.2000 4.8000 154.6000 5.2000 ;
	    RECT 156.8000 5.1000 157.1000 7.5000 ;
	    RECT 154.2000 4.2000 154.5000 4.8000 ;
	    RECT 156.7000 4.7000 157.1000 5.1000 ;
	    RECT 154.2000 3.8000 154.6000 4.2000 ;
	    RECT 162.2000 3.1000 162.6000 8.9000 ;
	    RECT 163.0000 8.1000 163.3000 12.8000 ;
	    RECT 164.6000 9.8000 165.0000 10.2000 ;
	    RECT 163.0000 7.8000 164.1000 8.1000 ;
	    RECT 163.8000 6.2000 164.1000 7.8000 ;
	    RECT 164.6000 7.2000 164.9000 9.8000 ;
	    RECT 164.6000 6.8000 165.0000 7.2000 ;
	    RECT 163.8000 5.8000 164.2000 6.2000 ;
	    RECT 167.0000 3.1000 167.4000 8.9000 ;
	    RECT 169.4000 8.2000 169.7000 12.8000 ;
	    RECT 175.8000 12.1000 176.2000 17.9000 ;
	    RECT 176.6000 15.8000 177.0000 16.2000 ;
	    RECT 176.6000 15.2000 176.9000 15.8000 ;
	    RECT 176.6000 14.8000 177.0000 15.2000 ;
	    RECT 179.8000 14.7000 180.2000 15.1000 ;
	    RECT 179.8000 14.2000 180.1000 14.7000 ;
	    RECT 179.8000 13.8000 180.2000 14.2000 ;
	    RECT 180.6000 12.1000 181.0000 17.9000 ;
	    RECT 181.4000 13.8000 181.8000 14.2000 ;
	    RECT 181.4000 10.2000 181.7000 13.8000 ;
	    RECT 182.2000 13.1000 182.6000 15.9000 ;
	    RECT 186.2000 15.2000 186.5000 30.8000 ;
	    RECT 189.4000 25.1000 189.8000 27.9000 ;
	    RECT 190.2000 27.2000 190.5000 31.8000 ;
	    RECT 190.2000 26.8000 190.6000 27.2000 ;
	    RECT 191.0000 23.1000 191.4000 28.9000 ;
	    RECT 194.2000 28.2000 194.5000 35.8000 ;
	    RECT 195.0000 33.1000 195.4000 35.9000 ;
	    RECT 195.8000 34.2000 196.1000 45.8000 ;
	    RECT 196.6000 43.1000 197.0000 48.9000 ;
	    RECT 199.0000 48.8000 199.4000 49.2000 ;
	    RECT 199.8000 48.8000 200.2000 49.2000 ;
	    RECT 199.0000 47.2000 199.3000 48.8000 ;
	    RECT 204.6000 47.2000 204.9000 52.8000 ;
	    RECT 205.4000 52.2000 205.7000 52.8000 ;
	    RECT 205.4000 51.8000 205.8000 52.2000 ;
	    RECT 207.0000 51.2000 207.3000 54.8000 ;
	    RECT 209.4000 53.1000 209.8000 55.9000 ;
	    RECT 210.2000 54.8000 210.6000 55.2000 ;
	    RECT 210.2000 54.2000 210.5000 54.8000 ;
	    RECT 210.2000 53.8000 210.6000 54.2000 ;
	    RECT 211.0000 52.1000 211.4000 57.9000 ;
	    RECT 211.8000 54.7000 212.2000 55.1000 ;
	    RECT 211.8000 53.2000 212.1000 54.7000 ;
	    RECT 211.8000 52.8000 212.2000 53.2000 ;
	    RECT 215.8000 52.1000 216.2000 57.9000 ;
	    RECT 216.6000 54.2000 216.9000 61.8000 ;
	    RECT 218.2000 56.8000 218.6000 57.2000 ;
	    RECT 218.2000 55.2000 218.5000 56.8000 ;
	    RECT 218.2000 54.8000 218.6000 55.2000 ;
	    RECT 216.6000 53.8000 217.0000 54.2000 ;
	    RECT 219.0000 53.1000 219.4000 55.9000 ;
	    RECT 219.0000 51.8000 219.4000 52.2000 ;
	    RECT 220.6000 52.1000 221.0000 57.9000 ;
	    RECT 221.4000 55.1000 221.7000 65.8000 ;
	    RECT 223.8000 65.1000 224.1000 65.8000 ;
	    RECT 227.0000 65.2000 227.3000 66.8000 ;
	    RECT 228.6000 65.8000 229.0000 66.2000 ;
	    RECT 229.4000 65.8000 229.8000 66.2000 ;
	    RECT 231.0000 65.8000 231.4000 66.2000 ;
	    RECT 228.6000 65.2000 228.9000 65.8000 ;
	    RECT 229.4000 65.2000 229.7000 65.8000 ;
	    RECT 224.6000 65.1000 225.0000 65.2000 ;
	    RECT 223.8000 64.8000 225.0000 65.1000 ;
	    RECT 227.0000 64.8000 227.4000 65.2000 ;
	    RECT 228.6000 64.8000 229.0000 65.2000 ;
	    RECT 229.4000 64.8000 229.8000 65.2000 ;
	    RECT 227.0000 59.1000 227.3000 64.8000 ;
	    RECT 231.0000 62.2000 231.3000 65.8000 ;
	    RECT 229.4000 61.8000 229.8000 62.2000 ;
	    RECT 231.0000 61.8000 231.4000 62.2000 ;
	    RECT 229.4000 59.2000 229.7000 61.8000 ;
	    RECT 233.4000 59.2000 233.7000 66.8000 ;
	    RECT 235.8000 65.8000 236.2000 66.2000 ;
	    RECT 235.8000 64.2000 236.1000 65.8000 ;
	    RECT 236.6000 65.2000 236.9000 66.8000 ;
	    RECT 237.4000 66.1000 237.8000 66.2000 ;
	    RECT 238.2000 66.1000 238.6000 66.2000 ;
	    RECT 237.4000 65.8000 238.6000 66.1000 ;
	    RECT 236.6000 64.8000 237.0000 65.2000 ;
	    RECT 235.8000 63.8000 236.2000 64.2000 ;
	    RECT 235.8000 62.2000 236.1000 63.8000 ;
	    RECT 235.8000 61.8000 236.2000 62.2000 ;
	    RECT 227.8000 59.1000 228.2000 59.2000 ;
	    RECT 227.0000 58.8000 228.2000 59.1000 ;
	    RECT 229.4000 58.8000 229.8000 59.2000 ;
	    RECT 233.4000 58.8000 233.8000 59.2000 ;
	    RECT 234.2000 59.1000 234.6000 59.2000 ;
	    RECT 235.0000 59.1000 235.4000 59.2000 ;
	    RECT 234.2000 58.8000 235.4000 59.1000 ;
	    RECT 221.4000 54.7000 221.8000 55.1000 ;
	    RECT 222.2000 53.8000 222.6000 54.2000 ;
	    RECT 207.0000 50.8000 207.4000 51.2000 ;
	    RECT 219.0000 49.2000 219.3000 51.8000 ;
	    RECT 206.2000 47.8000 206.6000 48.2000 ;
	    RECT 199.0000 46.8000 199.4000 47.2000 ;
	    RECT 201.4000 46.8000 201.8000 47.2000 ;
	    RECT 204.6000 46.8000 205.0000 47.2000 ;
	    RECT 201.4000 46.2000 201.7000 46.8000 ;
	    RECT 206.2000 46.2000 206.5000 47.8000 ;
	    RECT 209.4000 46.8000 209.8000 47.2000 ;
	    RECT 209.4000 46.2000 209.7000 46.8000 ;
	    RECT 201.4000 45.8000 201.8000 46.2000 ;
	    RECT 202.2000 45.8000 202.6000 46.2000 ;
	    RECT 203.0000 46.1000 203.4000 46.2000 ;
	    RECT 203.8000 46.1000 204.2000 46.2000 ;
	    RECT 203.0000 45.8000 204.2000 46.1000 ;
	    RECT 206.2000 45.8000 206.6000 46.2000 ;
	    RECT 209.4000 45.8000 209.8000 46.2000 ;
	    RECT 202.2000 39.2000 202.5000 45.8000 ;
	    RECT 202.2000 38.8000 202.6000 39.2000 ;
	    RECT 195.8000 33.8000 196.2000 34.2000 ;
	    RECT 195.8000 32.1000 196.1000 33.8000 ;
	    RECT 196.6000 32.1000 197.0000 37.9000 ;
	    RECT 197.4000 36.8000 197.8000 37.2000 ;
	    RECT 197.4000 35.1000 197.7000 36.8000 ;
	    RECT 197.4000 34.7000 197.8000 35.1000 ;
	    RECT 200.6000 33.8000 201.0000 34.2000 ;
	    RECT 200.6000 33.2000 200.9000 33.8000 ;
	    RECT 200.6000 32.8000 201.0000 33.2000 ;
	    RECT 201.4000 32.1000 201.8000 37.9000 ;
	    RECT 203.8000 36.8000 204.2000 37.2000 ;
	    RECT 203.8000 35.2000 204.1000 36.8000 ;
	    RECT 206.2000 36.2000 206.5000 45.8000 ;
	    RECT 210.2000 45.1000 210.6000 47.9000 ;
	    RECT 211.8000 43.1000 212.2000 48.9000 ;
	    RECT 212.6000 46.8000 213.0000 47.2000 ;
	    RECT 212.6000 46.3000 212.9000 46.8000 ;
	    RECT 212.6000 45.9000 213.0000 46.3000 ;
	    RECT 215.0000 46.1000 215.4000 46.2000 ;
	    RECT 215.8000 46.1000 216.2000 46.2000 ;
	    RECT 215.0000 45.8000 216.2000 46.1000 ;
	    RECT 216.6000 43.1000 217.0000 48.9000 ;
	    RECT 219.0000 48.8000 219.4000 49.2000 ;
	    RECT 219.8000 45.1000 220.2000 47.9000 ;
	    RECT 221.4000 43.1000 221.8000 48.9000 ;
	    RECT 222.2000 48.2000 222.5000 53.8000 ;
	    RECT 225.4000 52.1000 225.8000 57.9000 ;
	    RECT 228.6000 54.8000 229.0000 55.2000 ;
	    RECT 231.0000 55.1000 231.4000 55.2000 ;
	    RECT 231.8000 55.1000 232.2000 55.2000 ;
	    RECT 231.0000 54.8000 232.2000 55.1000 ;
	    RECT 228.6000 54.2000 228.9000 54.8000 ;
	    RECT 228.6000 53.8000 229.0000 54.2000 ;
	    RECT 230.2000 52.8000 230.6000 53.2000 ;
	    RECT 230.2000 52.2000 230.5000 52.8000 ;
	    RECT 230.2000 51.8000 230.6000 52.2000 ;
	    RECT 236.6000 52.1000 237.0000 57.9000 ;
	    RECT 239.0000 53.2000 239.3000 71.8000 ;
	    RECT 239.8000 65.2000 240.1000 73.8000 ;
	    RECT 247.1000 73.5000 247.4000 75.9000 ;
	    RECT 247.7000 74.9000 248.1000 75.3000 ;
	    RECT 247.8000 74.2000 248.1000 74.9000 ;
	    RECT 250.3000 74.2000 250.6000 75.9000 ;
	    RECT 255.0000 75.8000 255.4000 76.2000 ;
	    RECT 253.4000 75.1000 253.8000 75.2000 ;
	    RECT 253.4000 74.8000 254.5000 75.1000 ;
	    RECT 247.8000 73.9000 250.6000 74.2000 ;
	    RECT 247.8000 73.5000 248.2000 73.6000 ;
	    RECT 249.5000 73.5000 249.9000 73.6000 ;
	    RECT 250.3000 73.5000 250.6000 73.9000 ;
	    RECT 247.1000 73.2000 249.9000 73.5000 ;
	    RECT 240.6000 72.8000 241.0000 73.2000 ;
	    RECT 243.0000 73.1000 243.4000 73.2000 ;
	    RECT 243.8000 73.1000 244.2000 73.2000 ;
	    RECT 247.1000 73.1000 247.5000 73.2000 ;
	    RECT 250.2000 73.1000 250.6000 73.5000 ;
	    RECT 243.0000 72.8000 244.2000 73.1000 ;
	    RECT 240.6000 72.2000 240.9000 72.8000 ;
	    RECT 240.6000 71.8000 241.0000 72.2000 ;
	    RECT 242.2000 72.1000 242.6000 72.2000 ;
	    RECT 243.0000 72.1000 243.4000 72.2000 ;
	    RECT 242.2000 71.8000 243.4000 72.1000 ;
	    RECT 247.8000 72.1000 248.2000 72.2000 ;
	    RECT 248.6000 72.1000 249.0000 72.2000 ;
	    RECT 247.8000 71.8000 249.0000 72.1000 ;
	    RECT 243.8000 69.8000 244.2000 70.2000 ;
	    RECT 243.8000 68.2000 244.1000 69.8000 ;
	    RECT 242.2000 68.1000 242.6000 68.2000 ;
	    RECT 243.0000 68.1000 243.4000 68.2000 ;
	    RECT 242.2000 67.8000 243.4000 68.1000 ;
	    RECT 243.8000 67.8000 244.2000 68.2000 ;
	    RECT 245.4000 67.8000 245.8000 68.2000 ;
	    RECT 247.8000 67.8000 248.2000 68.2000 ;
	    RECT 249.4000 67.8000 249.8000 68.2000 ;
	    RECT 251.8000 67.8000 252.2000 68.2000 ;
	    RECT 245.4000 67.2000 245.7000 67.8000 ;
	    RECT 247.8000 67.2000 248.1000 67.8000 ;
	    RECT 241.4000 66.8000 241.8000 67.2000 ;
	    RECT 245.4000 66.8000 245.8000 67.2000 ;
	    RECT 247.8000 66.8000 248.2000 67.2000 ;
	    RECT 241.4000 66.2000 241.7000 66.8000 ;
	    RECT 241.4000 65.8000 241.8000 66.2000 ;
	    RECT 247.8000 66.1000 248.2000 66.2000 ;
	    RECT 248.6000 66.1000 249.0000 66.2000 ;
	    RECT 247.8000 65.8000 249.0000 66.1000 ;
	    RECT 239.8000 64.8000 240.2000 65.2000 ;
	    RECT 239.8000 59.2000 240.1000 64.8000 ;
	    RECT 248.6000 63.8000 249.0000 64.2000 ;
	    RECT 248.6000 63.2000 248.9000 63.8000 ;
	    RECT 244.6000 62.8000 245.0000 63.2000 ;
	    RECT 248.6000 62.8000 249.0000 63.2000 ;
	    RECT 244.6000 62.2000 244.9000 62.8000 ;
	    RECT 243.0000 61.8000 243.4000 62.2000 ;
	    RECT 244.6000 61.8000 245.0000 62.2000 ;
	    RECT 239.8000 58.8000 240.2000 59.2000 ;
	    RECT 240.6000 56.8000 241.0000 57.2000 ;
	    RECT 240.6000 55.1000 240.9000 56.8000 ;
	    RECT 240.6000 54.7000 241.0000 55.1000 ;
	    RECT 239.0000 52.8000 239.4000 53.2000 ;
	    RECT 229.4000 50.8000 229.8000 51.2000 ;
	    RECT 229.4000 49.2000 229.7000 50.8000 ;
	    RECT 239.0000 49.2000 239.3000 52.8000 ;
	    RECT 241.4000 52.1000 241.8000 57.9000 ;
	    RECT 243.0000 57.2000 243.3000 61.8000 ;
	    RECT 243.0000 56.8000 243.4000 57.2000 ;
	    RECT 242.2000 53.8000 242.6000 54.2000 ;
	    RECT 227.8000 49.1000 228.2000 49.2000 ;
	    RECT 228.6000 49.1000 229.0000 49.2000 ;
	    RECT 222.2000 47.8000 222.6000 48.2000 ;
	    RECT 222.2000 45.9000 222.6000 46.3000 ;
	    RECT 222.2000 42.1000 222.5000 45.9000 ;
	    RECT 221.4000 41.8000 222.5000 42.1000 ;
	    RECT 225.4000 45.8000 225.8000 46.2000 ;
	    RECT 221.4000 39.2000 221.7000 41.8000 ;
	    RECT 217.4000 39.1000 217.8000 39.2000 ;
	    RECT 218.2000 39.1000 218.6000 39.2000 ;
	    RECT 217.4000 38.8000 218.6000 39.1000 ;
	    RECT 221.4000 38.8000 221.8000 39.2000 ;
	    RECT 204.6000 35.8000 205.0000 36.2000 ;
	    RECT 206.2000 35.8000 206.6000 36.2000 ;
	    RECT 203.8000 34.8000 204.2000 35.2000 ;
	    RECT 204.6000 34.2000 204.9000 35.8000 ;
	    RECT 205.4000 35.1000 205.8000 35.2000 ;
	    RECT 206.2000 35.1000 206.6000 35.2000 ;
	    RECT 205.4000 34.8000 206.6000 35.1000 ;
	    RECT 207.8000 35.1000 208.2000 35.2000 ;
	    RECT 208.6000 35.1000 209.0000 35.2000 ;
	    RECT 207.8000 34.8000 209.0000 35.1000 ;
	    RECT 204.6000 33.8000 205.0000 34.2000 ;
	    RECT 209.4000 33.1000 209.8000 35.9000 ;
	    RECT 210.2000 33.8000 210.6000 34.2000 ;
	    RECT 210.2000 33.2000 210.5000 33.8000 ;
	    RECT 210.2000 32.8000 210.6000 33.2000 ;
	    RECT 195.0000 31.8000 196.1000 32.1000 ;
	    RECT 205.4000 31.8000 205.8000 32.2000 ;
	    RECT 211.0000 32.1000 211.4000 37.9000 ;
	    RECT 211.8000 35.8000 212.2000 36.2000 ;
	    RECT 211.8000 35.1000 212.1000 35.8000 ;
	    RECT 211.8000 34.7000 212.2000 35.1000 ;
	    RECT 215.8000 32.1000 216.2000 37.9000 ;
	    RECT 219.8000 34.8000 220.2000 35.2000 ;
	    RECT 219.0000 33.8000 219.4000 34.2000 ;
	    RECT 219.0000 33.2000 219.3000 33.8000 ;
	    RECT 219.0000 32.8000 219.4000 33.2000 ;
	    RECT 194.2000 27.8000 194.6000 28.2000 ;
	    RECT 195.0000 27.2000 195.3000 31.8000 ;
	    RECT 205.4000 29.2000 205.7000 31.8000 ;
	    RECT 219.8000 31.2000 220.1000 34.8000 ;
	    RECT 222.2000 33.1000 222.6000 35.9000 ;
	    RECT 223.0000 32.8000 223.4000 33.2000 ;
	    RECT 215.8000 30.8000 216.2000 31.2000 ;
	    RECT 219.8000 30.8000 220.2000 31.2000 ;
	    RECT 215.8000 29.2000 216.1000 30.8000 ;
	    RECT 223.0000 29.2000 223.3000 32.8000 ;
	    RECT 223.8000 32.1000 224.2000 37.9000 ;
	    RECT 224.6000 34.7000 225.0000 35.1000 ;
	    RECT 224.6000 34.2000 224.9000 34.7000 ;
	    RECT 225.4000 34.2000 225.7000 45.8000 ;
	    RECT 226.2000 43.1000 226.6000 48.9000 ;
	    RECT 227.8000 48.8000 229.0000 49.1000 ;
	    RECT 229.4000 48.8000 229.8000 49.2000 ;
	    RECT 231.8000 43.1000 232.2000 48.9000 ;
	    RECT 233.4000 48.8000 233.8000 49.2000 ;
	    RECT 232.6000 45.8000 233.0000 46.2000 ;
	    RECT 232.6000 45.2000 232.9000 45.8000 ;
	    RECT 232.6000 44.8000 233.0000 45.2000 ;
	    RECT 229.4000 41.8000 229.8000 42.2000 ;
	    RECT 224.6000 33.8000 225.0000 34.2000 ;
	    RECT 225.4000 33.8000 225.8000 34.2000 ;
	    RECT 224.6000 32.8000 225.0000 33.2000 ;
	    RECT 191.8000 26.8000 192.2000 27.2000 ;
	    RECT 192.6000 26.8000 193.0000 27.2000 ;
	    RECT 195.0000 26.8000 195.4000 27.2000 ;
	    RECT 187.8000 21.8000 188.2000 22.2000 ;
	    RECT 187.8000 16.2000 188.1000 21.8000 ;
	    RECT 187.8000 15.8000 188.2000 16.2000 ;
	    RECT 183.0000 14.8000 183.4000 15.2000 ;
	    RECT 184.6000 14.8000 185.0000 15.2000 ;
	    RECT 186.2000 14.8000 186.6000 15.2000 ;
	    RECT 188.6000 14.8000 189.0000 15.2000 ;
	    RECT 183.0000 13.2000 183.3000 14.8000 ;
	    RECT 184.6000 14.2000 184.9000 14.8000 ;
	    RECT 184.6000 13.8000 185.0000 14.2000 ;
	    RECT 183.0000 12.8000 183.4000 13.2000 ;
	    RECT 175.8000 9.8000 176.2000 10.2000 ;
	    RECT 181.4000 9.8000 181.8000 10.2000 ;
	    RECT 170.2000 8.8000 170.6000 9.2000 ;
	    RECT 171.8000 9.1000 172.2000 9.2000 ;
	    RECT 172.6000 9.1000 173.0000 9.2000 ;
	    RECT 171.8000 8.8000 173.0000 9.1000 ;
	    RECT 168.6000 5.1000 169.0000 7.9000 ;
	    RECT 169.4000 7.8000 169.8000 8.2000 ;
	    RECT 170.2000 7.2000 170.5000 8.8000 ;
	    RECT 170.2000 6.8000 170.6000 7.2000 ;
	    RECT 170.2000 6.2000 170.5000 6.8000 ;
	    RECT 170.2000 5.8000 170.6000 6.2000 ;
	    RECT 171.8000 5.8000 172.2000 6.2000 ;
	    RECT 171.8000 5.2000 172.1000 5.8000 ;
	    RECT 171.8000 4.8000 172.2000 5.2000 ;
	    RECT 175.0000 3.1000 175.4000 8.9000 ;
	    RECT 175.8000 6.2000 176.1000 9.8000 ;
	    RECT 175.8000 5.8000 176.2000 6.2000 ;
	    RECT 177.4000 6.1000 177.8000 6.2000 ;
	    RECT 178.2000 6.1000 178.6000 6.2000 ;
	    RECT 177.4000 5.8000 178.6000 6.1000 ;
	    RECT 179.8000 3.1000 180.2000 8.9000 ;
	    RECT 184.6000 8.8000 185.0000 9.2000 ;
	    RECT 184.6000 8.2000 184.9000 8.8000 ;
	    RECT 181.4000 5.1000 181.8000 7.9000 ;
	    RECT 184.6000 7.8000 185.0000 8.2000 ;
	    RECT 186.2000 5.2000 186.5000 14.8000 ;
	    RECT 188.6000 14.2000 188.9000 14.8000 ;
	    RECT 188.6000 13.8000 189.0000 14.2000 ;
	    RECT 189.4000 13.8000 189.8000 14.2000 ;
	    RECT 188.6000 13.1000 189.0000 13.2000 ;
	    RECT 189.4000 13.1000 189.7000 13.8000 ;
	    RECT 188.6000 12.8000 189.7000 13.1000 ;
	    RECT 189.4000 9.2000 189.7000 12.8000 ;
	    RECT 191.0000 10.1000 191.4000 10.2000 ;
	    RECT 191.8000 10.1000 192.1000 26.8000 ;
	    RECT 192.6000 26.2000 192.9000 26.8000 ;
	    RECT 192.6000 25.8000 193.0000 26.2000 ;
	    RECT 195.8000 23.1000 196.2000 28.9000 ;
	    RECT 204.6000 28.8000 205.0000 29.2000 ;
	    RECT 205.4000 28.8000 205.8000 29.2000 ;
	    RECT 215.8000 28.8000 216.2000 29.2000 ;
	    RECT 223.0000 28.8000 223.4000 29.2000 ;
	    RECT 200.6000 27.1000 201.0000 27.2000 ;
	    RECT 201.4000 27.1000 201.8000 27.2000 ;
	    RECT 200.6000 26.8000 201.8000 27.1000 ;
	    RECT 204.6000 26.2000 204.9000 28.8000 ;
	    RECT 207.8000 27.8000 208.2000 28.2000 ;
	    RECT 210.2000 27.8000 210.6000 28.2000 ;
	    RECT 214.2000 27.8000 214.6000 28.2000 ;
	    RECT 217.4000 27.8000 217.8000 28.2000 ;
	    RECT 207.8000 27.2000 208.1000 27.8000 ;
	    RECT 210.2000 27.2000 210.5000 27.8000 ;
	    RECT 207.8000 26.8000 208.2000 27.2000 ;
	    RECT 208.6000 26.8000 209.0000 27.2000 ;
	    RECT 210.2000 26.8000 210.6000 27.2000 ;
	    RECT 200.6000 26.1000 201.0000 26.2000 ;
	    RECT 201.4000 26.1000 201.8000 26.2000 ;
	    RECT 200.6000 25.8000 201.8000 26.1000 ;
	    RECT 203.8000 25.8000 204.2000 26.2000 ;
	    RECT 204.6000 25.8000 205.0000 26.2000 ;
	    RECT 207.0000 25.8000 207.4000 26.2000 ;
	    RECT 192.6000 15.1000 193.0000 15.2000 ;
	    RECT 193.4000 15.1000 193.8000 15.2000 ;
	    RECT 192.6000 14.8000 193.8000 15.1000 ;
	    RECT 195.0000 12.8000 195.4000 13.2000 ;
	    RECT 195.8000 13.1000 196.2000 15.9000 ;
	    RECT 195.0000 12.2000 195.3000 12.8000 ;
	    RECT 195.0000 11.8000 195.4000 12.2000 ;
	    RECT 197.4000 12.1000 197.8000 17.9000 ;
	    RECT 198.2000 15.8000 198.6000 16.2000 ;
	    RECT 200.6000 15.8000 201.0000 16.2000 ;
	    RECT 198.2000 14.2000 198.5000 15.8000 ;
	    RECT 199.0000 15.1000 199.4000 15.2000 ;
	    RECT 199.8000 15.1000 200.2000 15.2000 ;
	    RECT 199.0000 14.8000 200.2000 15.1000 ;
	    RECT 198.2000 13.8000 198.6000 14.2000 ;
	    RECT 191.0000 9.8000 192.1000 10.1000 ;
	    RECT 186.2000 4.8000 186.6000 5.2000 ;
	    RECT 187.0000 3.1000 187.4000 8.9000 ;
	    RECT 189.4000 8.8000 189.8000 9.2000 ;
	    RECT 191.0000 8.2000 191.3000 9.8000 ;
	    RECT 191.0000 7.8000 191.4000 8.2000 ;
	    RECT 191.0000 6.8000 191.4000 7.2000 ;
	    RECT 191.0000 6.3000 191.3000 6.8000 ;
	    RECT 191.0000 5.9000 191.4000 6.3000 ;
	    RECT 191.8000 3.1000 192.2000 8.9000 ;
	    RECT 198.2000 8.2000 198.5000 13.8000 ;
	    RECT 193.4000 5.1000 193.8000 7.9000 ;
	    RECT 194.2000 7.8000 194.6000 8.2000 ;
	    RECT 198.2000 7.8000 198.6000 8.2000 ;
	    RECT 194.2000 7.2000 194.5000 7.8000 ;
	    RECT 194.2000 6.8000 194.6000 7.2000 ;
	    RECT 195.8000 6.8000 196.2000 7.2000 ;
	    RECT 198.2000 6.8000 198.6000 7.2000 ;
	    RECT 195.8000 6.2000 196.1000 6.8000 ;
	    RECT 198.2000 6.2000 198.5000 6.8000 ;
	    RECT 200.6000 6.2000 200.9000 15.8000 ;
	    RECT 202.2000 12.1000 202.6000 17.9000 ;
	    RECT 203.8000 14.2000 204.1000 25.8000 ;
	    RECT 207.0000 24.2000 207.3000 25.8000 ;
	    RECT 207.0000 23.8000 207.4000 24.2000 ;
	    RECT 207.0000 19.2000 207.3000 23.8000 ;
	    RECT 207.0000 18.8000 207.4000 19.2000 ;
	    RECT 204.6000 17.1000 205.0000 17.2000 ;
	    RECT 205.4000 17.1000 205.8000 17.2000 ;
	    RECT 204.6000 16.8000 205.8000 17.1000 ;
	    RECT 208.6000 15.2000 208.9000 26.8000 ;
	    RECT 209.4000 25.8000 209.8000 26.2000 ;
	    RECT 209.4000 25.2000 209.7000 25.8000 ;
	    RECT 209.4000 24.8000 209.8000 25.2000 ;
	    RECT 211.0000 24.8000 211.4000 25.2000 ;
	    RECT 211.8000 25.1000 212.2000 25.2000 ;
	    RECT 212.6000 25.1000 213.0000 25.2000 ;
	    RECT 211.8000 24.8000 213.0000 25.1000 ;
	    RECT 211.0000 23.2000 211.3000 24.8000 ;
	    RECT 214.2000 24.2000 214.5000 27.8000 ;
	    RECT 217.4000 27.2000 217.7000 27.8000 ;
	    RECT 216.6000 26.8000 217.0000 27.2000 ;
	    RECT 217.4000 26.8000 217.8000 27.2000 ;
	    RECT 219.0000 27.1000 219.4000 27.2000 ;
	    RECT 219.8000 27.1000 220.2000 27.2000 ;
	    RECT 219.0000 26.8000 220.2000 27.1000 ;
	    RECT 221.4000 26.8000 221.8000 27.2000 ;
	    RECT 215.0000 24.8000 215.4000 25.2000 ;
	    RECT 214.2000 23.8000 214.6000 24.2000 ;
	    RECT 211.0000 22.8000 211.4000 23.2000 ;
	    RECT 215.0000 19.2000 215.3000 24.8000 ;
	    RECT 216.6000 24.2000 216.9000 26.8000 ;
	    RECT 221.4000 26.2000 221.7000 26.8000 ;
	    RECT 219.0000 25.8000 219.4000 26.2000 ;
	    RECT 221.4000 25.8000 221.8000 26.2000 ;
	    RECT 216.6000 23.8000 217.0000 24.2000 ;
	    RECT 215.0000 18.8000 215.4000 19.2000 ;
	    RECT 209.4000 16.8000 209.8000 17.2000 ;
	    RECT 209.4000 15.2000 209.7000 16.8000 ;
	    RECT 213.4000 15.8000 213.8000 16.2000 ;
	    RECT 205.4000 14.8000 205.8000 15.2000 ;
	    RECT 206.2000 14.8000 206.6000 15.2000 ;
	    RECT 207.8000 15.1000 208.2000 15.2000 ;
	    RECT 208.6000 15.1000 209.0000 15.2000 ;
	    RECT 207.8000 14.8000 209.0000 15.1000 ;
	    RECT 209.4000 14.8000 209.8000 15.2000 ;
	    RECT 210.2000 15.1000 210.6000 15.2000 ;
	    RECT 211.0000 15.1000 211.4000 15.2000 ;
	    RECT 210.2000 14.8000 211.4000 15.1000 ;
	    RECT 205.4000 14.2000 205.7000 14.8000 ;
	    RECT 206.2000 14.2000 206.5000 14.8000 ;
	    RECT 203.8000 13.8000 204.2000 14.2000 ;
	    RECT 205.4000 13.8000 205.8000 14.2000 ;
	    RECT 206.2000 13.8000 206.6000 14.2000 ;
	    RECT 210.2000 13.8000 210.6000 14.2000 ;
	    RECT 210.2000 13.2000 210.5000 13.8000 ;
	    RECT 210.2000 12.8000 210.6000 13.2000 ;
	    RECT 213.4000 12.2000 213.7000 15.8000 ;
	    RECT 218.2000 14.8000 218.6000 15.2000 ;
	    RECT 218.2000 14.2000 218.5000 14.8000 ;
	    RECT 219.0000 14.2000 219.3000 25.8000 ;
	    RECT 224.6000 25.1000 224.9000 32.8000 ;
	    RECT 225.4000 31.8000 225.8000 32.2000 ;
	    RECT 228.6000 32.1000 229.0000 37.9000 ;
	    RECT 229.4000 36.2000 229.7000 41.8000 ;
	    RECT 231.0000 39.1000 231.4000 39.2000 ;
	    RECT 231.8000 39.1000 232.2000 39.2000 ;
	    RECT 231.0000 38.8000 232.2000 39.1000 ;
	    RECT 233.4000 37.2000 233.7000 48.8000 ;
	    RECT 235.8000 45.9000 236.2000 46.3000 ;
	    RECT 235.8000 45.2000 236.1000 45.9000 ;
	    RECT 235.8000 44.8000 236.2000 45.2000 ;
	    RECT 236.6000 43.1000 237.0000 48.9000 ;
	    RECT 239.0000 48.8000 239.4000 49.2000 ;
	    RECT 238.2000 45.1000 238.6000 47.9000 ;
	    RECT 239.0000 44.8000 239.4000 45.2000 ;
	    RECT 233.4000 36.8000 233.8000 37.2000 ;
	    RECT 229.4000 35.8000 229.8000 36.2000 ;
	    RECT 231.8000 35.8000 232.2000 36.2000 ;
	    RECT 231.8000 35.1000 232.1000 35.8000 ;
	    RECT 231.0000 34.8000 232.1000 35.1000 ;
	    RECT 233.4000 35.2000 233.7000 36.8000 ;
	    RECT 238.2000 35.8000 238.6000 36.2000 ;
	    RECT 233.4000 34.8000 233.8000 35.2000 ;
	    RECT 234.2000 34.8000 234.6000 35.2000 ;
	    RECT 231.0000 33.2000 231.3000 34.8000 ;
	    RECT 234.2000 34.2000 234.5000 34.8000 ;
	    RECT 231.8000 34.1000 232.2000 34.2000 ;
	    RECT 232.6000 34.1000 233.0000 34.2000 ;
	    RECT 231.8000 33.8000 233.0000 34.1000 ;
	    RECT 234.2000 33.8000 234.6000 34.2000 ;
	    RECT 235.8000 33.8000 236.2000 34.2000 ;
	    RECT 235.8000 33.2000 236.1000 33.8000 ;
	    RECT 231.0000 32.8000 231.4000 33.2000 ;
	    RECT 235.8000 32.8000 236.2000 33.2000 ;
	    RECT 236.6000 31.8000 237.0000 32.2000 ;
	    RECT 225.4000 26.2000 225.7000 31.8000 ;
	    RECT 236.6000 31.2000 236.9000 31.8000 ;
	    RECT 236.6000 30.8000 237.0000 31.2000 ;
	    RECT 238.2000 30.2000 238.5000 35.8000 ;
	    RECT 239.0000 34.1000 239.3000 44.8000 ;
	    RECT 241.4000 43.1000 241.8000 48.9000 ;
	    RECT 242.2000 46.2000 242.5000 53.8000 ;
	    RECT 243.0000 53.1000 243.4000 55.9000 ;
	    RECT 245.4000 55.8000 245.8000 56.2000 ;
	    RECT 245.4000 55.1000 245.7000 55.8000 ;
	    RECT 246.2000 55.1000 246.6000 55.2000 ;
	    RECT 245.4000 54.8000 246.6000 55.1000 ;
	    RECT 249.4000 54.2000 249.7000 67.8000 ;
	    RECT 251.0000 66.8000 251.4000 67.2000 ;
	    RECT 251.0000 66.2000 251.3000 66.8000 ;
	    RECT 251.8000 66.2000 252.1000 67.8000 ;
	    RECT 254.2000 67.2000 254.5000 74.8000 ;
	    RECT 255.0000 68.2000 255.3000 75.8000 ;
	    RECT 255.8000 73.2000 256.1000 85.8000 ;
	    RECT 256.6000 85.1000 257.0000 85.2000 ;
	    RECT 257.4000 85.1000 257.8000 85.2000 ;
	    RECT 256.6000 84.8000 257.8000 85.1000 ;
	    RECT 259.1000 85.1000 259.4000 87.5000 ;
	    RECT 259.8000 87.4000 260.2000 87.5000 ;
	    RECT 261.5000 87.4000 261.9000 87.5000 ;
	    RECT 262.3000 87.1000 262.6000 87.5000 ;
	    RECT 259.8000 86.8000 262.6000 87.1000 ;
	    RECT 259.8000 86.1000 260.1000 86.8000 ;
	    RECT 259.7000 85.7000 260.1000 86.1000 ;
	    RECT 262.3000 85.1000 262.6000 86.8000 ;
	    RECT 259.1000 84.7000 259.5000 85.1000 ;
	    RECT 262.2000 84.7000 262.6000 85.1000 ;
	    RECT 264.6000 87.5000 265.0000 87.9000 ;
	    RECT 267.0000 87.8000 267.3000 93.8000 ;
	    RECT 268.6000 91.8000 269.0000 92.2000 ;
	    RECT 268.6000 90.2000 268.9000 91.8000 ;
	    RECT 268.6000 89.8000 269.0000 90.2000 ;
	    RECT 265.3000 87.5000 267.4000 87.8000 ;
	    RECT 267.9000 87.5000 268.3000 87.9000 ;
	    RECT 264.6000 87.1000 264.9000 87.5000 ;
	    RECT 265.3000 87.4000 265.7000 87.5000 ;
	    RECT 267.0000 87.4000 267.4000 87.5000 ;
	    RECT 264.6000 86.8000 267.0000 87.1000 ;
	    RECT 264.6000 85.1000 264.9000 86.8000 ;
	    RECT 266.6000 86.7000 267.0000 86.8000 ;
	    RECT 268.0000 85.1000 268.3000 87.5000 ;
	    RECT 264.6000 84.7000 265.0000 85.1000 ;
	    RECT 267.9000 84.7000 268.3000 85.1000 ;
	    RECT 268.6000 86.8000 269.0000 87.2000 ;
	    RECT 268.6000 84.1000 268.9000 86.8000 ;
	    RECT 267.8000 83.8000 268.9000 84.1000 ;
	    RECT 262.2000 82.8000 262.6000 83.2000 ;
	    RECT 256.6000 79.8000 257.0000 80.2000 ;
	    RECT 256.6000 75.2000 256.9000 79.8000 ;
	    RECT 262.2000 79.2000 262.5000 82.8000 ;
	    RECT 262.2000 78.8000 262.6000 79.2000 ;
	    RECT 257.4000 77.8000 257.8000 78.2000 ;
	    RECT 259.8000 77.8000 260.2000 78.2000 ;
	    RECT 257.4000 76.2000 257.7000 77.8000 ;
	    RECT 257.4000 75.8000 257.8000 76.2000 ;
	    RECT 259.0000 75.8000 259.4000 76.2000 ;
	    RECT 259.0000 75.2000 259.3000 75.8000 ;
	    RECT 256.6000 74.8000 257.0000 75.2000 ;
	    RECT 259.0000 74.8000 259.4000 75.2000 ;
	    RECT 259.8000 74.2000 260.1000 77.8000 ;
	    RECT 260.6000 76.8000 261.0000 77.2000 ;
	    RECT 260.6000 76.2000 260.9000 76.8000 ;
	    RECT 267.8000 76.2000 268.1000 83.8000 ;
	    RECT 268.6000 78.8000 269.0000 79.2000 ;
	    RECT 268.6000 78.2000 268.9000 78.8000 ;
	    RECT 268.6000 77.8000 269.0000 78.2000 ;
	    RECT 260.6000 75.8000 261.0000 76.2000 ;
	    RECT 265.4000 75.8000 265.8000 76.2000 ;
	    RECT 267.0000 76.1000 267.4000 76.2000 ;
	    RECT 267.8000 76.1000 268.2000 76.2000 ;
	    RECT 267.0000 75.8000 268.2000 76.1000 ;
	    RECT 265.4000 75.2000 265.7000 75.8000 ;
	    RECT 265.4000 74.8000 265.8000 75.2000 ;
	    RECT 259.8000 73.8000 260.2000 74.2000 ;
	    RECT 263.0000 73.8000 263.4000 74.2000 ;
	    RECT 263.0000 73.2000 263.3000 73.8000 ;
	    RECT 255.8000 72.8000 256.2000 73.2000 ;
	    RECT 259.0000 72.8000 259.4000 73.2000 ;
	    RECT 263.0000 72.8000 263.4000 73.2000 ;
	    RECT 259.0000 69.2000 259.3000 72.8000 ;
	    RECT 265.4000 71.2000 265.7000 74.8000 ;
	    RECT 269.4000 73.1000 269.8000 73.2000 ;
	    RECT 268.6000 72.8000 269.8000 73.1000 ;
	    RECT 267.0000 72.1000 267.4000 72.2000 ;
	    RECT 267.8000 72.1000 268.2000 72.2000 ;
	    RECT 267.0000 71.8000 268.2000 72.1000 ;
	    RECT 265.4000 70.8000 265.8000 71.2000 ;
	    RECT 267.8000 70.8000 268.2000 71.2000 ;
	    RECT 259.0000 68.8000 259.4000 69.2000 ;
	    RECT 255.0000 67.8000 255.4000 68.2000 ;
	    RECT 257.4000 67.8000 257.8000 68.2000 ;
	    RECT 257.4000 67.2000 257.7000 67.8000 ;
	    RECT 258.1000 67.5000 258.5000 67.9000 ;
	    RECT 259.0000 67.5000 261.1000 67.8000 ;
	    RECT 261.4000 67.5000 261.8000 67.9000 ;
	    RECT 252.6000 66.8000 253.0000 67.2000 ;
	    RECT 254.2000 66.8000 254.6000 67.2000 ;
	    RECT 257.4000 66.8000 257.8000 67.2000 ;
	    RECT 250.2000 65.8000 250.6000 66.2000 ;
	    RECT 251.0000 65.8000 251.4000 66.2000 ;
	    RECT 251.8000 65.8000 252.2000 66.2000 ;
	    RECT 250.2000 65.2000 250.5000 65.8000 ;
	    RECT 250.2000 64.8000 250.6000 65.2000 ;
	    RECT 251.8000 64.2000 252.1000 65.8000 ;
	    RECT 252.6000 65.2000 252.9000 66.8000 ;
	    RECT 252.6000 64.8000 253.0000 65.2000 ;
	    RECT 258.1000 65.1000 258.4000 67.5000 ;
	    RECT 259.0000 67.4000 259.4000 67.5000 ;
	    RECT 260.7000 67.4000 261.1000 67.5000 ;
	    RECT 261.5000 67.1000 261.8000 67.5000 ;
	    RECT 259.4000 66.8000 261.8000 67.1000 ;
	    RECT 259.4000 66.7000 259.8000 66.8000 ;
	    RECT 261.5000 65.1000 261.8000 66.8000 ;
	    RECT 263.0000 66.8000 263.4000 67.2000 ;
	    RECT 263.0000 66.2000 263.3000 66.8000 ;
	    RECT 263.0000 65.8000 263.4000 66.2000 ;
	    RECT 258.1000 64.7000 258.5000 65.1000 ;
	    RECT 261.4000 64.7000 261.8000 65.1000 ;
	    RECT 251.8000 63.8000 252.2000 64.2000 ;
	    RECT 261.4000 56.8000 261.8000 57.2000 ;
	    RECT 261.4000 56.2000 261.7000 56.8000 ;
	    RECT 259.8000 55.8000 260.2000 56.2000 ;
	    RECT 261.4000 55.8000 261.8000 56.2000 ;
	    RECT 259.8000 55.2000 260.1000 55.8000 ;
	    RECT 255.0000 54.8000 255.4000 55.2000 ;
	    RECT 259.8000 54.8000 260.2000 55.2000 ;
	    RECT 260.6000 54.8000 261.0000 55.2000 ;
	    RECT 244.6000 54.1000 245.0000 54.2000 ;
	    RECT 245.4000 54.1000 245.8000 54.2000 ;
	    RECT 244.6000 53.8000 245.8000 54.1000 ;
	    RECT 249.4000 53.8000 249.8000 54.2000 ;
	    RECT 243.8000 52.8000 244.2000 53.2000 ;
	    RECT 250.2000 53.1000 250.6000 53.2000 ;
	    RECT 251.0000 53.1000 251.4000 53.2000 ;
	    RECT 250.2000 52.8000 251.4000 53.1000 ;
	    RECT 243.8000 52.2000 244.1000 52.8000 ;
	    RECT 255.0000 52.2000 255.3000 54.8000 ;
	    RECT 260.6000 54.2000 260.9000 54.8000 ;
	    RECT 257.4000 53.8000 257.8000 54.2000 ;
	    RECT 258.2000 53.8000 258.6000 54.2000 ;
	    RECT 259.0000 54.1000 259.4000 54.2000 ;
	    RECT 259.8000 54.1000 260.2000 54.2000 ;
	    RECT 259.0000 53.8000 260.2000 54.1000 ;
	    RECT 260.6000 53.8000 261.0000 54.2000 ;
	    RECT 257.4000 53.2000 257.7000 53.8000 ;
	    RECT 258.2000 53.2000 258.5000 53.8000 ;
	    RECT 260.6000 53.2000 260.9000 53.8000 ;
	    RECT 256.6000 52.8000 257.0000 53.2000 ;
	    RECT 257.4000 52.8000 257.8000 53.2000 ;
	    RECT 258.2000 52.8000 258.6000 53.2000 ;
	    RECT 260.6000 52.8000 261.0000 53.2000 ;
	    RECT 243.8000 51.8000 244.2000 52.2000 ;
	    RECT 250.2000 51.8000 250.6000 52.2000 ;
	    RECT 251.8000 51.8000 252.2000 52.2000 ;
	    RECT 255.0000 51.8000 255.4000 52.2000 ;
	    RECT 255.8000 51.8000 256.2000 52.2000 ;
	    RECT 245.4000 47.8000 245.8000 48.2000 ;
	    RECT 243.0000 46.8000 243.4000 47.2000 ;
	    RECT 242.2000 45.8000 242.6000 46.2000 ;
	    RECT 242.2000 45.2000 242.5000 45.8000 ;
	    RECT 242.2000 44.8000 242.6000 45.2000 ;
	    RECT 239.8000 36.8000 240.2000 37.2000 ;
	    RECT 239.8000 35.2000 240.1000 36.8000 ;
	    RECT 243.0000 35.2000 243.3000 46.8000 ;
	    RECT 245.4000 46.3000 245.7000 47.8000 ;
	    RECT 245.4000 45.9000 245.8000 46.3000 ;
	    RECT 246.2000 43.1000 246.6000 48.9000 ;
	    RECT 250.2000 48.2000 250.5000 51.8000 ;
	    RECT 251.8000 49.2000 252.1000 51.8000 ;
	    RECT 255.8000 49.2000 256.1000 51.8000 ;
	    RECT 256.6000 49.2000 256.9000 52.8000 ;
	    RECT 259.8000 50.8000 260.2000 51.2000 ;
	    RECT 251.0000 48.8000 251.4000 49.2000 ;
	    RECT 251.8000 48.8000 252.2000 49.2000 ;
	    RECT 255.0000 48.8000 255.4000 49.2000 ;
	    RECT 255.8000 48.8000 256.2000 49.2000 ;
	    RECT 256.6000 48.8000 257.0000 49.2000 ;
	    RECT 251.0000 48.2000 251.3000 48.8000 ;
	    RECT 247.8000 45.1000 248.2000 47.9000 ;
	    RECT 250.2000 47.8000 250.6000 48.2000 ;
	    RECT 251.0000 47.8000 251.4000 48.2000 ;
	    RECT 248.6000 46.8000 249.0000 47.2000 ;
	    RECT 253.4000 47.1000 253.8000 47.2000 ;
	    RECT 254.2000 47.1000 254.6000 47.2000 ;
	    RECT 253.4000 46.8000 254.6000 47.1000 ;
	    RECT 248.6000 46.2000 248.9000 46.8000 ;
	    RECT 248.6000 45.8000 249.0000 46.2000 ;
	    RECT 253.4000 45.8000 253.8000 46.2000 ;
	    RECT 253.4000 45.2000 253.7000 45.8000 ;
	    RECT 250.2000 44.8000 250.6000 45.2000 ;
	    RECT 251.8000 45.1000 252.2000 45.2000 ;
	    RECT 252.6000 45.1000 253.0000 45.2000 ;
	    RECT 251.8000 44.8000 253.0000 45.1000 ;
	    RECT 253.4000 44.8000 253.8000 45.2000 ;
	    RECT 250.2000 43.2000 250.5000 44.8000 ;
	    RECT 250.2000 42.8000 250.6000 43.2000 ;
	    RECT 246.2000 35.8000 246.6000 36.2000 ;
	    RECT 246.2000 35.2000 246.5000 35.8000 ;
	    RECT 239.8000 34.8000 240.2000 35.2000 ;
	    RECT 243.0000 34.8000 243.4000 35.2000 ;
	    RECT 246.2000 34.8000 246.6000 35.2000 ;
	    RECT 247.0000 34.8000 247.4000 35.2000 ;
	    RECT 239.0000 33.8000 240.1000 34.1000 ;
	    RECT 238.2000 29.8000 238.6000 30.2000 ;
	    RECT 239.8000 29.2000 240.1000 33.8000 ;
	    RECT 240.6000 33.8000 241.0000 34.2000 ;
	    RECT 242.2000 33.8000 242.6000 34.2000 ;
	    RECT 240.6000 30.2000 240.9000 33.8000 ;
	    RECT 242.2000 33.2000 242.5000 33.8000 ;
	    RECT 242.2000 32.8000 242.6000 33.2000 ;
	    RECT 242.2000 32.1000 242.6000 32.2000 ;
	    RECT 243.0000 32.1000 243.3000 34.8000 ;
	    RECT 247.0000 34.2000 247.3000 34.8000 ;
	    RECT 245.4000 34.1000 245.8000 34.2000 ;
	    RECT 246.2000 34.1000 246.6000 34.2000 ;
	    RECT 245.4000 33.8000 246.6000 34.1000 ;
	    RECT 247.0000 33.8000 247.4000 34.2000 ;
	    RECT 243.8000 33.1000 244.2000 33.2000 ;
	    RECT 244.6000 33.1000 245.0000 33.2000 ;
	    RECT 243.8000 32.8000 245.0000 33.1000 ;
	    RECT 242.2000 31.8000 243.3000 32.1000 ;
	    RECT 244.6000 31.8000 245.0000 32.2000 ;
	    RECT 240.6000 29.8000 241.0000 30.2000 ;
	    RECT 242.2000 29.2000 242.5000 31.8000 ;
	    RECT 243.0000 29.8000 243.4000 30.2000 ;
	    RECT 232.6000 29.1000 233.0000 29.2000 ;
	    RECT 233.4000 29.1000 233.8000 29.2000 ;
	    RECT 232.6000 28.8000 233.8000 29.1000 ;
	    RECT 239.0000 28.8000 239.4000 29.2000 ;
	    RECT 239.8000 28.8000 240.2000 29.2000 ;
	    RECT 242.2000 28.8000 242.6000 29.2000 ;
	    RECT 228.6000 28.1000 229.0000 28.2000 ;
	    RECT 229.4000 28.1000 229.8000 28.2000 ;
	    RECT 228.6000 27.8000 229.8000 28.1000 ;
	    RECT 231.0000 28.1000 231.4000 28.2000 ;
	    RECT 231.8000 28.1000 232.2000 28.2000 ;
	    RECT 231.0000 27.8000 232.2000 28.1000 ;
	    RECT 232.6000 27.8000 233.0000 28.2000 ;
	    RECT 237.4000 27.8000 237.8000 28.2000 ;
	    RECT 232.6000 27.2000 232.9000 27.8000 ;
	    RECT 237.4000 27.2000 237.7000 27.8000 ;
	    RECT 239.0000 27.2000 239.3000 28.8000 ;
	    RECT 240.6000 27.8000 241.0000 28.2000 ;
	    RECT 226.2000 26.8000 226.6000 27.2000 ;
	    RECT 227.0000 26.8000 227.4000 27.2000 ;
	    RECT 229.4000 27.1000 229.8000 27.2000 ;
	    RECT 230.2000 27.1000 230.6000 27.2000 ;
	    RECT 229.4000 26.8000 230.6000 27.1000 ;
	    RECT 232.6000 26.8000 233.0000 27.2000 ;
	    RECT 234.2000 26.8000 234.6000 27.2000 ;
	    RECT 237.4000 26.8000 237.8000 27.2000 ;
	    RECT 239.0000 26.8000 239.4000 27.2000 ;
	    RECT 226.2000 26.2000 226.5000 26.8000 ;
	    RECT 227.0000 26.2000 227.3000 26.8000 ;
	    RECT 225.4000 25.8000 225.8000 26.2000 ;
	    RECT 226.2000 25.8000 226.6000 26.2000 ;
	    RECT 227.0000 25.8000 227.4000 26.2000 ;
	    RECT 227.8000 26.1000 228.2000 26.2000 ;
	    RECT 228.6000 26.1000 229.0000 26.2000 ;
	    RECT 227.8000 25.8000 229.0000 26.1000 ;
	    RECT 224.6000 24.8000 225.7000 25.1000 ;
	    RECT 224.6000 18.8000 225.0000 19.2000 ;
	    RECT 222.2000 17.1000 222.6000 17.2000 ;
	    RECT 223.0000 17.1000 223.4000 17.2000 ;
	    RECT 222.2000 16.8000 223.4000 17.1000 ;
	    RECT 224.6000 16.2000 224.9000 18.8000 ;
	    RECT 224.6000 15.8000 225.0000 16.2000 ;
	    RECT 219.8000 14.8000 220.2000 15.2000 ;
	    RECT 222.2000 15.1000 222.6000 15.2000 ;
	    RECT 223.0000 15.1000 223.4000 15.2000 ;
	    RECT 222.2000 14.8000 223.4000 15.1000 ;
	    RECT 223.8000 15.1000 224.2000 15.2000 ;
	    RECT 224.6000 15.1000 225.0000 15.2000 ;
	    RECT 223.8000 14.8000 225.0000 15.1000 ;
	    RECT 219.8000 14.2000 220.1000 14.8000 ;
	    RECT 214.2000 13.8000 214.6000 14.2000 ;
	    RECT 215.8000 13.8000 216.2000 14.2000 ;
	    RECT 216.6000 13.8000 217.0000 14.2000 ;
	    RECT 218.2000 13.8000 218.6000 14.2000 ;
	    RECT 219.0000 13.8000 219.4000 14.2000 ;
	    RECT 219.8000 13.8000 220.2000 14.2000 ;
	    RECT 213.4000 11.8000 213.8000 12.2000 ;
	    RECT 205.4000 9.8000 205.8000 10.2000 ;
	    RECT 203.8000 7.8000 204.2000 8.2000 ;
	    RECT 203.8000 7.2000 204.1000 7.8000 ;
	    RECT 202.2000 6.8000 202.6000 7.2000 ;
	    RECT 203.8000 6.8000 204.2000 7.2000 ;
	    RECT 202.2000 6.2000 202.5000 6.8000 ;
	    RECT 195.8000 5.8000 196.2000 6.2000 ;
	    RECT 197.4000 5.8000 197.8000 6.2000 ;
	    RECT 198.2000 5.8000 198.6000 6.2000 ;
	    RECT 200.6000 5.8000 201.0000 6.2000 ;
	    RECT 202.2000 5.8000 202.6000 6.2000 ;
	    RECT 197.4000 5.2000 197.7000 5.8000 ;
	    RECT 200.6000 5.2000 200.9000 5.8000 ;
	    RECT 197.4000 4.8000 197.8000 5.2000 ;
	    RECT 200.6000 4.8000 201.0000 5.2000 ;
	    RECT 204.6000 5.1000 205.0000 7.9000 ;
	    RECT 205.4000 7.2000 205.7000 9.8000 ;
	    RECT 214.2000 9.2000 214.5000 13.8000 ;
	    RECT 215.8000 11.2000 216.1000 13.8000 ;
	    RECT 216.6000 13.2000 216.9000 13.8000 ;
	    RECT 216.6000 12.8000 217.0000 13.2000 ;
	    RECT 223.8000 13.1000 224.2000 13.2000 ;
	    RECT 224.6000 13.1000 225.0000 13.2000 ;
	    RECT 223.8000 12.8000 225.0000 13.1000 ;
	    RECT 221.4000 11.8000 221.8000 12.2000 ;
	    RECT 215.8000 10.8000 216.2000 11.2000 ;
	    RECT 221.4000 10.2000 221.7000 11.8000 ;
	    RECT 221.4000 9.8000 221.8000 10.2000 ;
	    RECT 205.4000 6.8000 205.8000 7.2000 ;
	    RECT 206.2000 3.1000 206.6000 8.9000 ;
	    RECT 207.0000 5.9000 207.4000 6.3000 ;
	    RECT 207.0000 5.2000 207.3000 5.9000 ;
	    RECT 207.0000 4.8000 207.4000 5.2000 ;
	    RECT 211.0000 3.1000 211.4000 8.9000 ;
	    RECT 213.4000 8.8000 213.8000 9.2000 ;
	    RECT 214.2000 8.8000 214.6000 9.2000 ;
	    RECT 217.4000 9.1000 217.8000 9.2000 ;
	    RECT 218.2000 9.1000 218.6000 9.2000 ;
	    RECT 217.4000 8.8000 218.6000 9.1000 ;
	    RECT 213.4000 7.2000 213.7000 8.8000 ;
	    RECT 213.4000 6.8000 213.8000 7.2000 ;
	    RECT 215.8000 6.1000 216.2000 6.2000 ;
	    RECT 216.6000 6.1000 217.0000 6.2000 ;
	    RECT 215.8000 5.8000 217.0000 6.1000 ;
	    RECT 219.8000 3.1000 220.2000 8.9000 ;
	    RECT 222.2000 7.8000 222.6000 8.2000 ;
	    RECT 223.8000 7.8000 224.2000 8.2000 ;
	    RECT 222.2000 7.2000 222.5000 7.8000 ;
	    RECT 222.2000 6.8000 222.6000 7.2000 ;
	    RECT 223.8000 6.3000 224.1000 7.8000 ;
	    RECT 223.8000 5.9000 224.2000 6.3000 ;
	    RECT 224.6000 3.1000 225.0000 8.9000 ;
	    RECT 225.4000 7.2000 225.7000 24.8000 ;
	    RECT 228.6000 24.8000 229.0000 25.2000 ;
	    RECT 232.6000 24.8000 233.0000 25.2000 ;
	    RECT 234.2000 25.1000 234.5000 26.8000 ;
	    RECT 236.6000 26.1000 237.0000 26.2000 ;
	    RECT 237.4000 26.1000 237.8000 26.2000 ;
	    RECT 236.6000 25.8000 237.8000 26.1000 ;
	    RECT 238.2000 25.8000 238.6000 26.2000 ;
	    RECT 238.2000 25.2000 238.5000 25.8000 ;
	    RECT 235.0000 25.1000 235.4000 25.2000 ;
	    RECT 234.2000 24.8000 235.4000 25.1000 ;
	    RECT 236.6000 25.1000 237.0000 25.2000 ;
	    RECT 237.4000 25.1000 237.8000 25.2000 ;
	    RECT 236.6000 24.8000 237.8000 25.1000 ;
	    RECT 238.2000 24.8000 238.6000 25.2000 ;
	    RECT 228.6000 24.1000 228.9000 24.8000 ;
	    RECT 228.6000 23.8000 229.7000 24.1000 ;
	    RECT 227.8000 17.1000 228.2000 17.2000 ;
	    RECT 228.6000 17.1000 229.0000 17.2000 ;
	    RECT 227.8000 16.8000 229.0000 17.1000 ;
	    RECT 228.6000 14.8000 229.0000 15.2000 ;
	    RECT 228.6000 14.2000 228.9000 14.8000 ;
	    RECT 229.4000 14.2000 229.7000 23.8000 ;
	    RECT 231.0000 16.8000 231.4000 17.2000 ;
	    RECT 231.0000 16.2000 231.3000 16.8000 ;
	    RECT 231.0000 15.8000 231.4000 16.2000 ;
	    RECT 226.2000 14.1000 226.6000 14.2000 ;
	    RECT 227.0000 14.1000 227.4000 14.2000 ;
	    RECT 226.2000 13.8000 227.4000 14.1000 ;
	    RECT 228.6000 13.8000 229.0000 14.2000 ;
	    RECT 229.4000 13.8000 229.8000 14.2000 ;
	    RECT 229.4000 13.2000 229.7000 13.8000 ;
	    RECT 229.4000 12.8000 229.8000 13.2000 ;
	    RECT 232.6000 10.1000 232.9000 24.8000 ;
	    RECT 234.2000 22.8000 234.6000 23.2000 ;
	    RECT 234.2000 19.2000 234.5000 22.8000 ;
	    RECT 234.2000 18.8000 234.6000 19.2000 ;
	    RECT 235.0000 17.2000 235.3000 24.8000 ;
	    RECT 240.6000 17.2000 240.9000 27.8000 ;
	    RECT 243.0000 27.2000 243.3000 29.8000 ;
	    RECT 244.6000 29.2000 244.9000 31.8000 ;
	    RECT 244.6000 28.8000 245.0000 29.2000 ;
	    RECT 244.5000 27.5000 244.9000 27.9000 ;
	    RECT 245.4000 27.5000 247.5000 27.8000 ;
	    RECT 247.8000 27.5000 248.2000 27.9000 ;
	    RECT 243.0000 27.1000 243.4000 27.2000 ;
	    RECT 242.2000 26.8000 243.4000 27.1000 ;
	    RECT 243.8000 26.8000 244.2000 27.2000 ;
	    RECT 235.0000 16.8000 235.4000 17.2000 ;
	    RECT 240.6000 16.8000 241.0000 17.2000 ;
	    RECT 237.4000 15.8000 237.8000 16.2000 ;
	    RECT 235.8000 15.1000 236.2000 15.2000 ;
	    RECT 236.6000 15.1000 237.0000 15.2000 ;
	    RECT 235.8000 14.8000 237.0000 15.1000 ;
	    RECT 234.2000 13.8000 234.6000 14.2000 ;
	    RECT 234.2000 11.2000 234.5000 13.8000 ;
	    RECT 237.4000 13.2000 237.7000 15.8000 ;
	    RECT 240.6000 15.2000 240.9000 16.8000 ;
	    RECT 239.0000 15.1000 239.4000 15.2000 ;
	    RECT 239.8000 15.1000 240.2000 15.2000 ;
	    RECT 239.0000 14.8000 240.2000 15.1000 ;
	    RECT 240.6000 14.8000 241.0000 15.2000 ;
	    RECT 237.4000 12.8000 237.8000 13.2000 ;
	    RECT 234.2000 10.8000 234.6000 11.2000 ;
	    RECT 233.4000 10.1000 233.8000 10.2000 ;
	    RECT 232.6000 9.8000 233.8000 10.1000 ;
	    RECT 227.0000 8.8000 227.4000 9.2000 ;
	    RECT 227.0000 8.2000 227.3000 8.8000 ;
	    RECT 233.4000 8.2000 233.7000 9.8000 ;
	    RECT 225.4000 6.8000 225.8000 7.2000 ;
	    RECT 226.2000 5.1000 226.6000 7.9000 ;
	    RECT 227.0000 7.8000 227.4000 8.2000 ;
	    RECT 229.4000 7.8000 229.8000 8.2000 ;
	    RECT 233.4000 7.8000 233.8000 8.2000 ;
	    RECT 229.4000 7.2000 229.7000 7.8000 ;
	    RECT 227.8000 7.1000 228.2000 7.2000 ;
	    RECT 228.6000 7.1000 229.0000 7.2000 ;
	    RECT 227.8000 6.8000 229.0000 7.1000 ;
	    RECT 229.4000 6.8000 229.8000 7.2000 ;
	    RECT 231.8000 6.8000 232.2000 7.2000 ;
	    RECT 231.8000 6.2000 232.1000 6.8000 ;
	    RECT 239.0000 6.2000 239.3000 14.8000 ;
	    RECT 242.2000 14.2000 242.5000 26.8000 ;
	    RECT 243.8000 26.2000 244.1000 26.8000 ;
	    RECT 243.8000 25.8000 244.2000 26.2000 ;
	    RECT 244.5000 25.1000 244.8000 27.5000 ;
	    RECT 245.4000 27.4000 245.8000 27.5000 ;
	    RECT 247.1000 27.4000 247.5000 27.5000 ;
	    RECT 247.9000 27.1000 248.2000 27.5000 ;
	    RECT 245.8000 26.8000 248.2000 27.1000 ;
	    RECT 248.6000 27.8000 249.0000 28.2000 ;
	    RECT 248.6000 27.2000 248.9000 27.8000 ;
	    RECT 248.6000 26.8000 249.0000 27.2000 ;
	    RECT 245.8000 26.7000 246.2000 26.8000 ;
	    RECT 246.2000 25.8000 246.6000 26.2000 ;
	    RECT 244.5000 24.7000 244.9000 25.1000 ;
	    RECT 243.0000 23.8000 243.4000 24.2000 ;
	    RECT 244.6000 23.8000 245.0000 24.2000 ;
	    RECT 243.0000 16.2000 243.3000 23.8000 ;
	    RECT 243.0000 15.8000 243.4000 16.2000 ;
	    RECT 240.6000 14.1000 241.0000 14.2000 ;
	    RECT 241.4000 14.1000 241.8000 14.2000 ;
	    RECT 240.6000 13.8000 241.8000 14.1000 ;
	    RECT 242.2000 13.8000 242.6000 14.2000 ;
	    RECT 242.2000 13.2000 242.5000 13.8000 ;
	    RECT 242.2000 12.8000 242.6000 13.2000 ;
	    RECT 241.4000 11.8000 241.8000 12.2000 ;
	    RECT 243.8000 11.8000 244.2000 12.2000 ;
	    RECT 241.4000 10.2000 241.7000 11.8000 ;
	    RECT 241.4000 9.8000 241.8000 10.2000 ;
	    RECT 241.4000 8.8000 241.8000 9.2000 ;
	    RECT 241.4000 8.2000 241.7000 8.8000 ;
	    RECT 241.4000 7.8000 241.8000 8.2000 ;
	    RECT 243.8000 6.2000 244.1000 11.8000 ;
	    RECT 244.6000 7.2000 244.9000 23.8000 ;
	    RECT 246.2000 19.2000 246.5000 25.8000 ;
	    RECT 247.9000 25.1000 248.2000 26.8000 ;
	    RECT 247.8000 24.7000 248.2000 25.1000 ;
	    RECT 248.6000 25.8000 249.0000 26.2000 ;
	    RECT 248.6000 25.2000 248.9000 25.8000 ;
	    RECT 248.6000 24.8000 249.0000 25.2000 ;
	    RECT 249.4000 25.1000 249.8000 27.9000 ;
	    RECT 250.2000 27.2000 250.5000 42.8000 ;
	    RECT 254.2000 38.2000 254.5000 46.8000 ;
	    RECT 255.0000 46.2000 255.3000 48.8000 ;
	    RECT 256.6000 48.1000 257.0000 48.2000 ;
	    RECT 257.4000 48.1000 257.8000 48.2000 ;
	    RECT 256.6000 47.8000 257.8000 48.1000 ;
	    RECT 255.8000 46.8000 256.2000 47.2000 ;
	    RECT 255.0000 45.8000 255.4000 46.2000 ;
	    RECT 254.2000 37.8000 254.6000 38.2000 ;
	    RECT 255.0000 36.1000 255.3000 45.8000 ;
	    RECT 255.8000 45.2000 256.1000 46.8000 ;
	    RECT 255.8000 44.8000 256.2000 45.2000 ;
	    RECT 255.8000 40.2000 256.1000 44.8000 ;
	    RECT 258.2000 42.1000 258.6000 42.2000 ;
	    RECT 259.0000 42.1000 259.4000 42.2000 ;
	    RECT 258.2000 41.8000 259.4000 42.1000 ;
	    RECT 255.8000 39.8000 256.2000 40.2000 ;
	    RECT 259.0000 37.8000 259.4000 38.2000 ;
	    RECT 255.8000 36.1000 256.2000 36.2000 ;
	    RECT 255.0000 35.8000 256.2000 36.1000 ;
	    RECT 258.2000 35.8000 258.6000 36.2000 ;
	    RECT 258.2000 35.2000 258.5000 35.8000 ;
	    RECT 254.2000 34.8000 254.6000 35.2000 ;
	    RECT 258.2000 34.8000 258.6000 35.2000 ;
	    RECT 254.2000 29.2000 254.5000 34.8000 ;
	    RECT 259.0000 34.2000 259.3000 37.8000 ;
	    RECT 255.0000 34.1000 255.4000 34.2000 ;
	    RECT 255.8000 34.1000 256.2000 34.2000 ;
	    RECT 255.0000 33.8000 256.2000 34.1000 ;
	    RECT 259.0000 33.8000 259.4000 34.2000 ;
	    RECT 256.6000 31.8000 257.0000 32.2000 ;
	    RECT 256.6000 31.2000 256.9000 31.8000 ;
	    RECT 256.6000 30.8000 257.0000 31.2000 ;
	    RECT 259.0000 29.8000 259.4000 30.2000 ;
	    RECT 250.2000 26.8000 250.6000 27.2000 ;
	    RECT 251.0000 23.1000 251.4000 28.9000 ;
	    RECT 254.2000 28.8000 254.6000 29.2000 ;
	    RECT 257.4000 29.1000 257.8000 29.2000 ;
	    RECT 258.2000 29.1000 258.6000 29.2000 ;
	    RECT 254.2000 28.2000 254.5000 28.8000 ;
	    RECT 254.2000 27.8000 254.6000 28.2000 ;
	    RECT 255.0000 27.8000 255.4000 28.2000 ;
	    RECT 255.0000 27.2000 255.3000 27.8000 ;
	    RECT 255.0000 26.8000 255.4000 27.2000 ;
	    RECT 251.8000 25.9000 252.2000 26.3000 ;
	    RECT 251.8000 25.2000 252.1000 25.9000 ;
	    RECT 251.8000 24.8000 252.2000 25.2000 ;
	    RECT 255.8000 23.1000 256.2000 28.9000 ;
	    RECT 257.4000 28.8000 258.6000 29.1000 ;
	    RECT 259.0000 28.2000 259.3000 29.8000 ;
	    RECT 259.8000 29.2000 260.1000 50.8000 ;
	    RECT 265.4000 50.2000 265.7000 70.8000 ;
	    RECT 267.8000 69.2000 268.1000 70.8000 ;
	    RECT 267.8000 68.8000 268.2000 69.2000 ;
	    RECT 266.2000 66.8000 266.6000 67.2000 ;
	    RECT 266.2000 66.2000 266.5000 66.8000 ;
	    RECT 266.2000 65.8000 266.6000 66.2000 ;
	    RECT 266.2000 54.1000 266.6000 54.2000 ;
	    RECT 267.0000 54.1000 267.4000 54.2000 ;
	    RECT 266.2000 53.8000 267.4000 54.1000 ;
	    RECT 267.0000 53.1000 267.4000 53.2000 ;
	    RECT 267.8000 53.1000 268.2000 53.2000 ;
	    RECT 267.0000 52.8000 268.2000 53.1000 ;
	    RECT 265.4000 49.8000 265.8000 50.2000 ;
	    RECT 267.8000 49.8000 268.2000 50.2000 ;
	    RECT 260.6000 43.1000 261.0000 48.9000 ;
	    RECT 261.4000 45.8000 261.8000 46.2000 ;
	    RECT 264.6000 45.9000 265.0000 46.3000 ;
	    RECT 261.4000 43.2000 261.7000 45.8000 ;
	    RECT 261.4000 42.8000 261.8000 43.2000 ;
	    RECT 261.4000 39.8000 261.8000 40.2000 ;
	    RECT 261.4000 36.2000 261.7000 39.8000 ;
	    RECT 264.6000 39.2000 264.9000 45.9000 ;
	    RECT 265.4000 43.1000 265.8000 48.9000 ;
	    RECT 267.0000 45.1000 267.4000 47.9000 ;
	    RECT 267.8000 45.2000 268.1000 49.8000 ;
	    RECT 268.6000 49.2000 268.9000 72.8000 ;
	    RECT 268.6000 48.8000 269.0000 49.2000 ;
	    RECT 269.4000 47.8000 269.8000 48.2000 ;
	    RECT 267.8000 44.8000 268.2000 45.2000 ;
	    RECT 264.6000 38.8000 265.0000 39.2000 ;
	    RECT 261.4000 35.8000 261.8000 36.2000 ;
	    RECT 262.2000 35.8000 262.6000 36.2000 ;
	    RECT 267.8000 35.8000 268.2000 36.2000 ;
	    RECT 261.4000 35.2000 261.7000 35.8000 ;
	    RECT 262.2000 35.2000 262.5000 35.8000 ;
	    RECT 260.6000 34.8000 261.0000 35.2000 ;
	    RECT 261.4000 34.8000 261.8000 35.2000 ;
	    RECT 262.2000 34.8000 262.6000 35.2000 ;
	    RECT 260.6000 34.2000 260.9000 34.8000 ;
	    RECT 260.6000 33.8000 261.0000 34.2000 ;
	    RECT 262.2000 30.1000 262.5000 34.8000 ;
	    RECT 263.0000 34.1000 263.4000 34.2000 ;
	    RECT 263.8000 34.1000 264.2000 34.2000 ;
	    RECT 263.0000 33.8000 264.2000 34.1000 ;
	    RECT 266.2000 33.8000 266.6000 34.2000 ;
	    RECT 263.8000 32.8000 264.2000 33.2000 ;
	    RECT 264.6000 32.8000 265.0000 33.2000 ;
	    RECT 263.8000 32.2000 264.1000 32.8000 ;
	    RECT 263.8000 31.8000 264.2000 32.2000 ;
	    RECT 262.2000 29.8000 263.3000 30.1000 ;
	    RECT 259.8000 28.8000 260.2000 29.2000 ;
	    RECT 257.4000 27.8000 257.8000 28.2000 ;
	    RECT 259.0000 27.8000 259.4000 28.2000 ;
	    RECT 255.8000 21.8000 256.2000 22.2000 ;
	    RECT 255.8000 19.2000 256.1000 21.8000 ;
	    RECT 257.4000 19.2000 257.7000 27.8000 ;
	    RECT 260.6000 25.1000 261.0000 27.9000 ;
	    RECT 261.4000 26.8000 261.8000 27.2000 ;
	    RECT 261.4000 26.2000 261.7000 26.8000 ;
	    RECT 261.4000 25.8000 261.8000 26.2000 ;
	    RECT 246.2000 18.8000 246.6000 19.2000 ;
	    RECT 247.8000 18.8000 248.2000 19.2000 ;
	    RECT 250.2000 18.8000 250.6000 19.2000 ;
	    RECT 255.8000 18.8000 256.2000 19.2000 ;
	    RECT 257.4000 18.8000 257.8000 19.2000 ;
	    RECT 247.8000 16.2000 248.1000 18.8000 ;
	    RECT 247.8000 15.8000 248.2000 16.2000 ;
	    RECT 246.2000 15.1000 246.6000 15.2000 ;
	    RECT 247.0000 15.1000 247.4000 15.2000 ;
	    RECT 246.2000 14.8000 247.4000 15.1000 ;
	    RECT 248.6000 14.8000 249.0000 15.2000 ;
	    RECT 248.6000 14.2000 248.9000 14.8000 ;
	    RECT 250.2000 14.2000 250.5000 18.8000 ;
	    RECT 251.0000 17.8000 251.4000 18.2000 ;
	    RECT 251.0000 17.2000 251.3000 17.8000 ;
	    RECT 251.0000 16.8000 251.4000 17.2000 ;
	    RECT 251.8000 15.8000 252.2000 16.2000 ;
	    RECT 252.6000 15.8000 253.0000 16.2000 ;
	    RECT 251.8000 15.2000 252.1000 15.8000 ;
	    RECT 252.6000 15.2000 252.9000 15.8000 ;
	    RECT 251.8000 14.8000 252.2000 15.2000 ;
	    RECT 252.6000 14.8000 253.0000 15.2000 ;
	    RECT 259.0000 14.8000 259.4000 15.2000 ;
	    RECT 259.0000 14.2000 259.3000 14.8000 ;
	    RECT 245.4000 14.1000 245.8000 14.2000 ;
	    RECT 246.2000 14.1000 246.6000 14.2000 ;
	    RECT 245.4000 13.8000 246.6000 14.1000 ;
	    RECT 248.6000 13.8000 249.0000 14.2000 ;
	    RECT 250.2000 13.8000 250.6000 14.2000 ;
	    RECT 256.6000 13.8000 257.0000 14.2000 ;
	    RECT 259.0000 13.8000 259.4000 14.2000 ;
	    RECT 248.6000 12.8000 249.0000 13.2000 ;
	    RECT 248.6000 7.2000 248.9000 12.8000 ;
	    RECT 249.4000 7.8000 249.8000 8.2000 ;
	    RECT 244.6000 6.8000 245.0000 7.2000 ;
	    RECT 245.4000 6.8000 245.8000 7.2000 ;
	    RECT 248.6000 6.8000 249.0000 7.2000 ;
	    RECT 245.4000 6.2000 245.7000 6.8000 ;
	    RECT 249.4000 6.2000 249.7000 7.8000 ;
	    RECT 250.2000 7.2000 250.5000 13.8000 ;
	    RECT 256.6000 13.2000 256.9000 13.8000 ;
	    RECT 252.6000 12.8000 253.0000 13.2000 ;
	    RECT 255.0000 12.8000 255.4000 13.2000 ;
	    RECT 256.6000 12.8000 257.0000 13.2000 ;
	    RECT 257.4000 12.8000 257.8000 13.2000 ;
	    RECT 260.6000 13.1000 261.0000 15.9000 ;
	    RECT 261.4000 14.2000 261.7000 25.8000 ;
	    RECT 262.2000 23.1000 262.6000 28.9000 ;
	    RECT 261.4000 13.8000 261.8000 14.2000 ;
	    RECT 251.0000 11.8000 251.4000 12.2000 ;
	    RECT 251.0000 8.2000 251.3000 11.8000 ;
	    RECT 252.6000 9.2000 252.9000 12.8000 ;
	    RECT 255.0000 12.2000 255.3000 12.8000 ;
	    RECT 255.0000 11.8000 255.4000 12.2000 ;
	    RECT 255.0000 10.8000 255.4000 11.2000 ;
	    RECT 253.4000 9.8000 253.8000 10.2000 ;
	    RECT 252.6000 8.8000 253.0000 9.2000 ;
	    RECT 253.4000 8.2000 253.7000 9.8000 ;
	    RECT 255.0000 9.2000 255.3000 10.8000 ;
	    RECT 257.4000 10.2000 257.7000 12.8000 ;
	    RECT 262.2000 12.1000 262.6000 17.9000 ;
	    RECT 257.4000 9.8000 257.8000 10.2000 ;
	    RECT 255.0000 8.8000 255.4000 9.2000 ;
	    RECT 257.4000 8.8000 257.8000 9.2000 ;
	    RECT 261.4000 9.1000 261.8000 9.2000 ;
	    RECT 262.2000 9.1000 262.6000 9.2000 ;
	    RECT 261.4000 8.8000 262.6000 9.1000 ;
	    RECT 257.4000 8.2000 257.7000 8.8000 ;
	    RECT 251.0000 7.8000 251.4000 8.2000 ;
	    RECT 252.6000 8.1000 253.0000 8.2000 ;
	    RECT 253.4000 8.1000 253.8000 8.2000 ;
	    RECT 252.6000 7.8000 253.8000 8.1000 ;
	    RECT 255.8000 8.1000 256.2000 8.2000 ;
	    RECT 256.6000 8.1000 257.0000 8.2000 ;
	    RECT 255.8000 7.8000 257.0000 8.1000 ;
	    RECT 257.4000 7.8000 257.8000 8.2000 ;
	    RECT 259.0000 8.1000 259.4000 8.2000 ;
	    RECT 259.8000 8.1000 260.2000 8.2000 ;
	    RECT 259.0000 7.8000 260.2000 8.1000 ;
	    RECT 250.2000 6.8000 250.6000 7.2000 ;
	    RECT 251.8000 6.8000 252.2000 7.2000 ;
	    RECT 255.8000 6.8000 256.2000 7.2000 ;
	    RECT 251.8000 6.2000 252.1000 6.8000 ;
	    RECT 255.8000 6.2000 256.1000 6.8000 ;
	    RECT 263.0000 6.2000 263.3000 29.8000 ;
	    RECT 263.8000 26.8000 264.2000 27.2000 ;
	    RECT 263.8000 26.2000 264.1000 26.8000 ;
	    RECT 263.8000 25.8000 264.2000 26.2000 ;
	    RECT 263.8000 15.8000 264.2000 16.2000 ;
	    RECT 263.8000 15.2000 264.1000 15.8000 ;
	    RECT 263.8000 14.8000 264.2000 15.2000 ;
	    RECT 264.6000 9.2000 264.9000 32.8000 ;
	    RECT 265.4000 31.8000 265.8000 32.2000 ;
	    RECT 264.6000 8.8000 265.0000 9.2000 ;
	    RECT 265.4000 8.2000 265.7000 31.8000 ;
	    RECT 266.2000 28.2000 266.5000 33.8000 ;
	    RECT 267.8000 33.2000 268.1000 35.8000 ;
	    RECT 267.8000 32.8000 268.2000 33.2000 ;
	    RECT 269.4000 29.2000 269.7000 47.8000 ;
	    RECT 266.2000 27.8000 266.6000 28.2000 ;
	    RECT 267.0000 23.1000 267.4000 28.9000 ;
	    RECT 269.4000 28.8000 269.8000 29.2000 ;
	    RECT 267.0000 12.1000 267.4000 17.9000 ;
	    RECT 267.8000 11.8000 268.2000 12.2000 ;
	    RECT 268.6000 12.1000 269.0000 12.2000 ;
	    RECT 269.4000 12.1000 269.8000 12.2000 ;
	    RECT 268.6000 11.8000 269.8000 12.1000 ;
	    RECT 263.8000 7.8000 264.2000 8.2000 ;
	    RECT 265.4000 7.8000 265.8000 8.2000 ;
	    RECT 263.8000 7.2000 264.1000 7.8000 ;
	    RECT 263.8000 6.8000 264.2000 7.2000 ;
	    RECT 228.6000 6.1000 229.0000 6.2000 ;
	    RECT 229.4000 6.1000 229.8000 6.2000 ;
	    RECT 228.6000 5.8000 229.8000 6.1000 ;
	    RECT 231.8000 5.8000 232.2000 6.2000 ;
	    RECT 232.6000 6.1000 233.0000 6.2000 ;
	    RECT 233.4000 6.1000 233.8000 6.2000 ;
	    RECT 232.6000 5.8000 233.8000 6.1000 ;
	    RECT 235.8000 6.1000 236.2000 6.2000 ;
	    RECT 236.6000 6.1000 237.0000 6.2000 ;
	    RECT 235.8000 5.8000 237.0000 6.1000 ;
	    RECT 239.0000 5.8000 239.4000 6.2000 ;
	    RECT 239.8000 5.8000 240.2000 6.2000 ;
	    RECT 242.2000 6.1000 242.6000 6.2000 ;
	    RECT 243.0000 6.1000 243.4000 6.2000 ;
	    RECT 242.2000 5.8000 243.4000 6.1000 ;
	    RECT 243.8000 5.8000 244.2000 6.2000 ;
	    RECT 245.4000 5.8000 245.8000 6.2000 ;
	    RECT 249.4000 5.8000 249.8000 6.2000 ;
	    RECT 251.8000 5.8000 252.2000 6.2000 ;
	    RECT 254.2000 6.1000 254.6000 6.2000 ;
	    RECT 255.0000 6.1000 255.4000 6.2000 ;
	    RECT 254.2000 5.8000 255.4000 6.1000 ;
	    RECT 255.8000 5.8000 256.2000 6.2000 ;
	    RECT 260.6000 5.8000 261.0000 6.2000 ;
	    RECT 263.0000 5.8000 263.4000 6.2000 ;
	    RECT 239.8000 5.2000 240.1000 5.8000 ;
	    RECT 260.6000 5.2000 260.9000 5.8000 ;
	    RECT 265.4000 5.2000 265.7000 7.8000 ;
	    RECT 267.8000 6.2000 268.1000 11.8000 ;
	    RECT 269.4000 10.8000 269.8000 11.2000 ;
	    RECT 269.4000 9.2000 269.7000 10.8000 ;
	    RECT 268.6000 8.8000 269.0000 9.2000 ;
	    RECT 269.4000 8.8000 269.8000 9.2000 ;
	    RECT 268.6000 8.2000 268.9000 8.8000 ;
	    RECT 268.6000 7.8000 269.0000 8.2000 ;
	    RECT 267.8000 5.8000 268.2000 6.2000 ;
	    RECT 239.8000 4.8000 240.2000 5.2000 ;
	    RECT 246.2000 5.1000 246.6000 5.2000 ;
	    RECT 247.0000 5.1000 247.4000 5.2000 ;
	    RECT 246.2000 4.8000 247.4000 5.1000 ;
	    RECT 260.6000 4.8000 261.0000 5.2000 ;
	    RECT 261.4000 5.1000 261.8000 5.2000 ;
	    RECT 262.2000 5.1000 262.6000 5.2000 ;
	    RECT 261.4000 4.8000 262.6000 5.1000 ;
	    RECT 265.4000 4.8000 265.8000 5.2000 ;
         LAYER metal3 ;
	    RECT 202.2000 178.1000 202.6000 178.2000 ;
	    RECT 215.8000 178.1000 216.2000 178.2000 ;
	    RECT 250.2000 178.1000 250.6000 178.2000 ;
	    RECT 202.2000 177.8000 250.6000 178.1000 ;
	    RECT 183.8000 177.1000 184.2000 177.2000 ;
	    RECT 187.0000 177.1000 187.4000 177.2000 ;
	    RECT 183.8000 176.8000 187.4000 177.1000 ;
	    RECT 205.4000 176.8000 205.8000 177.2000 ;
	    RECT 222.2000 176.8000 222.6000 177.2000 ;
	    RECT 1.4000 176.1000 1.8000 176.2000 ;
	    RECT 5.4000 176.1000 5.8000 176.2000 ;
	    RECT 1.4000 175.8000 5.8000 176.1000 ;
	    RECT 9.4000 176.1000 9.8000 176.2000 ;
	    RECT 10.2000 176.1000 10.6000 176.2000 ;
	    RECT 9.4000 175.8000 10.6000 176.1000 ;
	    RECT 89.4000 176.1000 89.8000 176.2000 ;
	    RECT 93.4000 176.1000 93.8000 176.2000 ;
	    RECT 89.4000 175.8000 93.8000 176.1000 ;
	    RECT 205.4000 176.1000 205.7000 176.8000 ;
	    RECT 208.6000 176.1000 209.0000 176.2000 ;
	    RECT 205.4000 175.8000 209.0000 176.1000 ;
	    RECT 222.2000 176.1000 222.5000 176.8000 ;
	    RECT 238.2000 176.1000 238.6000 176.2000 ;
	    RECT 222.2000 175.8000 238.6000 176.1000 ;
	    RECT 254.2000 176.1000 254.6000 176.2000 ;
	    RECT 266.2000 176.1000 266.6000 176.2000 ;
	    RECT 254.2000 175.8000 266.6000 176.1000 ;
	    RECT 65.4000 175.1000 65.8000 175.2000 ;
	    RECT 58.2000 174.8000 65.8000 175.1000 ;
	    RECT 83.8000 175.1000 84.2000 175.2000 ;
	    RECT 91.0000 175.1000 91.4000 175.2000 ;
	    RECT 83.8000 174.8000 91.4000 175.1000 ;
	    RECT 91.8000 175.1000 92.2000 175.2000 ;
	    RECT 92.6000 175.1000 93.0000 175.2000 ;
	    RECT 91.8000 174.8000 93.0000 175.1000 ;
	    RECT 106.2000 175.1000 106.6000 175.2000 ;
	    RECT 107.0000 175.1000 107.4000 175.2000 ;
	    RECT 106.2000 174.8000 107.4000 175.1000 ;
	    RECT 114.2000 175.1000 114.6000 175.2000 ;
	    RECT 129.4000 175.1000 129.8000 175.2000 ;
	    RECT 114.2000 174.8000 129.8000 175.1000 ;
	    RECT 154.2000 175.1000 154.6000 175.2000 ;
	    RECT 165.4000 175.1000 165.8000 175.2000 ;
	    RECT 166.2000 175.1000 166.6000 175.2000 ;
	    RECT 154.2000 174.8000 166.6000 175.1000 ;
	    RECT 183.8000 175.1000 184.2000 175.2000 ;
	    RECT 219.0000 175.1000 219.4000 175.2000 ;
	    RECT 183.8000 174.8000 219.4000 175.1000 ;
	    RECT 219.8000 175.1000 220.2000 175.2000 ;
	    RECT 223.0000 175.1000 223.4000 175.2000 ;
	    RECT 219.8000 174.8000 223.4000 175.1000 ;
	    RECT 223.8000 175.1000 224.2000 175.2000 ;
	    RECT 224.6000 175.1000 225.0000 175.2000 ;
	    RECT 223.8000 174.8000 225.0000 175.1000 ;
	    RECT 227.8000 175.1000 228.2000 175.2000 ;
	    RECT 239.8000 175.1000 240.2000 175.2000 ;
	    RECT 243.0000 175.1000 243.4000 175.2000 ;
	    RECT 227.8000 174.8000 232.2000 175.1000 ;
	    RECT 239.8000 174.8000 243.4000 175.1000 ;
	    RECT 255.0000 175.1000 255.4000 175.2000 ;
	    RECT 255.0000 174.8000 259.3000 175.1000 ;
	    RECT 58.2000 174.2000 58.5000 174.8000 ;
	    RECT 231.8000 174.7000 232.2000 174.8000 ;
	    RECT 259.0000 174.2000 259.3000 174.8000 ;
	    RECT 6.2000 174.1000 6.6000 174.2000 ;
	    RECT 8.6000 174.1000 9.0000 174.2000 ;
	    RECT 6.2000 173.8000 9.0000 174.1000 ;
	    RECT 26.2000 174.1000 26.6000 174.2000 ;
	    RECT 30.2000 174.1000 30.6000 174.2000 ;
	    RECT 26.2000 173.8000 30.6000 174.1000 ;
	    RECT 58.2000 173.8000 58.6000 174.2000 ;
	    RECT 91.8000 174.1000 92.2000 174.2000 ;
	    RECT 101.4000 174.1000 101.8000 174.2000 ;
	    RECT 119.8000 174.1000 120.2000 174.2000 ;
	    RECT 91.8000 173.8000 99.3000 174.1000 ;
	    RECT 101.4000 173.8000 120.2000 174.1000 ;
	    RECT 120.6000 174.1000 121.0000 174.2000 ;
	    RECT 127.0000 174.1000 127.4000 174.2000 ;
	    RECT 120.6000 173.8000 127.4000 174.1000 ;
	    RECT 160.6000 174.1000 161.0000 174.2000 ;
	    RECT 167.0000 174.1000 167.4000 174.2000 ;
	    RECT 160.6000 173.8000 167.4000 174.1000 ;
	    RECT 171.8000 174.1000 172.2000 174.2000 ;
	    RECT 185.4000 174.1000 185.8000 174.2000 ;
	    RECT 171.8000 173.8000 185.8000 174.1000 ;
	    RECT 199.0000 174.1000 199.4000 174.2000 ;
	    RECT 199.8000 174.1000 200.2000 174.2000 ;
	    RECT 199.0000 173.8000 200.2000 174.1000 ;
	    RECT 200.6000 173.8000 201.0000 174.2000 ;
	    RECT 217.4000 174.1000 217.8000 174.2000 ;
	    RECT 219.0000 174.1000 219.4000 174.2000 ;
	    RECT 217.4000 173.8000 219.4000 174.1000 ;
	    RECT 222.2000 174.1000 222.6000 174.2000 ;
	    RECT 223.0000 174.1000 223.4000 174.2000 ;
	    RECT 222.2000 173.8000 223.4000 174.1000 ;
	    RECT 223.8000 174.1000 224.2000 174.2000 ;
	    RECT 225.4000 174.1000 225.8000 174.2000 ;
	    RECT 223.8000 173.8000 225.8000 174.1000 ;
	    RECT 239.0000 174.1000 239.4000 174.2000 ;
	    RECT 240.6000 174.1000 241.0000 174.2000 ;
	    RECT 239.0000 173.8000 241.0000 174.1000 ;
	    RECT 243.0000 174.1000 243.4000 174.2000 ;
	    RECT 247.0000 174.1000 247.4000 174.2000 ;
	    RECT 248.6000 174.1000 249.0000 174.2000 ;
	    RECT 243.0000 173.8000 249.0000 174.1000 ;
	    RECT 259.0000 173.8000 259.4000 174.2000 ;
	    RECT 99.0000 173.2000 99.3000 173.8000 ;
	    RECT 200.6000 173.2000 200.9000 173.8000 ;
	    RECT 99.0000 172.8000 99.4000 173.2000 ;
	    RECT 164.6000 173.1000 165.0000 173.2000 ;
	    RECT 175.0000 173.1000 175.4000 173.2000 ;
	    RECT 164.6000 172.8000 175.4000 173.1000 ;
	    RECT 177.4000 173.1000 177.8000 173.2000 ;
	    RECT 183.8000 173.1000 184.2000 173.2000 ;
	    RECT 177.4000 172.8000 184.2000 173.1000 ;
	    RECT 200.6000 172.8000 201.0000 173.2000 ;
	    RECT 205.4000 173.1000 205.8000 173.2000 ;
	    RECT 227.0000 173.1000 227.4000 173.2000 ;
	    RECT 205.4000 172.8000 227.4000 173.1000 ;
	    RECT 242.2000 173.1000 242.6000 173.2000 ;
	    RECT 245.4000 173.1000 245.8000 173.2000 ;
	    RECT 242.2000 172.8000 245.8000 173.1000 ;
	    RECT 249.4000 173.1000 249.8000 173.2000 ;
	    RECT 250.2000 173.1000 250.6000 173.2000 ;
	    RECT 249.4000 172.8000 250.6000 173.1000 ;
	    RECT 265.4000 173.1000 265.8000 173.2000 ;
	    RECT 267.0000 173.1000 267.4000 173.2000 ;
	    RECT 265.4000 172.8000 267.4000 173.1000 ;
	    RECT 13.4000 172.1000 13.8000 172.2000 ;
	    RECT 14.2000 172.1000 14.6000 172.2000 ;
	    RECT 20.6000 172.1000 21.0000 172.2000 ;
	    RECT 27.0000 172.1000 27.4000 172.2000 ;
	    RECT 30.2000 172.1000 30.6000 172.2000 ;
	    RECT 13.4000 171.8000 14.6000 172.1000 ;
	    RECT 19.8000 171.8000 30.6000 172.1000 ;
	    RECT 49.4000 172.1000 49.8000 172.2000 ;
	    RECT 52.6000 172.1000 53.0000 172.2000 ;
	    RECT 62.2000 172.1000 62.6000 172.2000 ;
	    RECT 49.4000 171.8000 62.6000 172.1000 ;
	    RECT 107.8000 172.1000 108.2000 172.2000 ;
	    RECT 111.8000 172.1000 112.2000 172.2000 ;
	    RECT 107.8000 171.8000 112.2000 172.1000 ;
	    RECT 120.6000 172.1000 121.0000 172.2000 ;
	    RECT 129.4000 172.1000 129.8000 172.2000 ;
	    RECT 133.4000 172.1000 133.8000 172.2000 ;
	    RECT 120.6000 171.8000 133.8000 172.1000 ;
	    RECT 139.8000 172.1000 140.2000 172.2000 ;
	    RECT 140.6000 172.1000 141.0000 172.2000 ;
	    RECT 147.0000 172.1000 147.4000 172.2000 ;
	    RECT 139.8000 171.8000 147.4000 172.1000 ;
	    RECT 175.0000 172.1000 175.3000 172.8000 ;
	    RECT 191.0000 172.1000 191.4000 172.2000 ;
	    RECT 175.0000 171.8000 191.4000 172.1000 ;
	    RECT 203.8000 172.1000 204.2000 172.2000 ;
	    RECT 215.8000 172.1000 216.2000 172.2000 ;
	    RECT 203.8000 171.8000 216.2000 172.1000 ;
	    RECT 219.0000 172.1000 219.4000 172.2000 ;
	    RECT 220.6000 172.1000 221.0000 172.2000 ;
	    RECT 219.0000 171.8000 221.0000 172.1000 ;
	    RECT 222.2000 172.1000 222.6000 172.2000 ;
	    RECT 224.6000 172.1000 225.0000 172.2000 ;
	    RECT 222.2000 171.8000 225.0000 172.1000 ;
	    RECT 239.0000 172.1000 239.4000 172.2000 ;
	    RECT 243.0000 172.1000 243.4000 172.2000 ;
	    RECT 246.2000 172.1000 246.6000 172.2000 ;
	    RECT 260.6000 172.1000 261.0000 172.2000 ;
	    RECT 239.0000 171.8000 243.4000 172.1000 ;
	    RECT 245.4000 171.8000 261.0000 172.1000 ;
	    RECT 111.8000 171.1000 112.2000 171.2000 ;
	    RECT 116.6000 171.1000 117.0000 171.2000 ;
	    RECT 111.8000 170.8000 117.0000 171.1000 ;
	    RECT 203.0000 171.1000 203.4000 171.2000 ;
	    RECT 207.0000 171.1000 207.4000 171.2000 ;
	    RECT 203.0000 170.8000 207.4000 171.1000 ;
	    RECT 219.0000 171.1000 219.4000 171.2000 ;
	    RECT 252.6000 171.1000 253.0000 171.2000 ;
	    RECT 219.0000 170.8000 253.0000 171.1000 ;
	    RECT 121.4000 169.8000 121.8000 170.2000 ;
	    RECT 193.4000 170.1000 193.8000 170.2000 ;
	    RECT 206.2000 170.1000 206.6000 170.2000 ;
	    RECT 193.4000 169.8000 206.6000 170.1000 ;
	    RECT 214.2000 170.1000 214.6000 170.2000 ;
	    RECT 215.0000 170.1000 215.4000 170.2000 ;
	    RECT 214.2000 169.8000 215.4000 170.1000 ;
	    RECT 215.8000 170.1000 216.2000 170.2000 ;
	    RECT 220.6000 170.1000 221.0000 170.2000 ;
	    RECT 215.8000 169.8000 221.0000 170.1000 ;
	    RECT 222.2000 170.1000 222.6000 170.2000 ;
	    RECT 263.8000 170.1000 264.2000 170.2000 ;
	    RECT 222.2000 169.8000 264.2000 170.1000 ;
	    RECT 106.2000 169.1000 106.6000 169.2000 ;
	    RECT 115.0000 169.1000 115.4000 169.2000 ;
	    RECT 106.2000 168.8000 115.4000 169.1000 ;
	    RECT 121.4000 169.1000 121.7000 169.8000 ;
	    RECT 125.4000 169.1000 125.8000 169.2000 ;
	    RECT 131.0000 169.1000 131.4000 169.2000 ;
	    RECT 121.4000 168.8000 131.4000 169.1000 ;
	    RECT 153.4000 169.1000 153.8000 169.2000 ;
	    RECT 154.2000 169.1000 154.6000 169.2000 ;
	    RECT 153.4000 168.8000 154.6000 169.1000 ;
	    RECT 171.8000 169.1000 172.2000 169.2000 ;
	    RECT 180.6000 169.1000 181.0000 169.2000 ;
	    RECT 171.8000 168.8000 181.0000 169.1000 ;
	    RECT 200.6000 169.1000 201.0000 169.2000 ;
	    RECT 208.6000 169.1000 209.0000 169.2000 ;
	    RECT 218.2000 169.1000 218.6000 169.2000 ;
	    RECT 200.6000 168.8000 218.6000 169.1000 ;
	    RECT 223.0000 169.1000 223.4000 169.2000 ;
	    RECT 227.0000 169.1000 227.4000 169.2000 ;
	    RECT 235.8000 169.1000 236.2000 169.2000 ;
	    RECT 239.0000 169.1000 239.4000 169.2000 ;
	    RECT 240.6000 169.1000 241.0000 169.2000 ;
	    RECT 244.6000 169.1000 245.0000 169.2000 ;
	    RECT 223.0000 168.8000 227.4000 169.1000 ;
	    RECT 235.0000 168.8000 239.4000 169.1000 ;
	    RECT 239.8000 168.8000 245.0000 169.1000 ;
	    RECT 245.4000 169.1000 245.8000 169.2000 ;
	    RECT 247.0000 169.1000 247.4000 169.2000 ;
	    RECT 245.4000 168.8000 247.4000 169.1000 ;
	    RECT 247.8000 169.1000 248.2000 169.2000 ;
	    RECT 253.4000 169.1000 253.8000 169.2000 ;
	    RECT 247.8000 168.8000 253.8000 169.1000 ;
	    RECT 255.8000 169.1000 256.2000 169.2000 ;
	    RECT 257.4000 169.1000 257.8000 169.2000 ;
	    RECT 255.8000 168.8000 257.8000 169.1000 ;
	    RECT 31.8000 168.1000 32.2000 168.2000 ;
	    RECT 35.0000 168.1000 35.4000 168.2000 ;
	    RECT 31.8000 167.8000 35.4000 168.1000 ;
	    RECT 43.0000 168.1000 43.4000 168.2000 ;
	    RECT 47.0000 168.1000 47.4000 168.2000 ;
	    RECT 51.0000 168.1000 51.4000 168.2000 ;
	    RECT 43.0000 167.8000 51.4000 168.1000 ;
	    RECT 67.8000 168.1000 68.2000 168.2000 ;
	    RECT 72.6000 168.1000 73.0000 168.2000 ;
	    RECT 88.6000 168.1000 89.0000 168.2000 ;
	    RECT 67.8000 167.8000 89.0000 168.1000 ;
	    RECT 107.8000 167.8000 108.2000 168.2000 ;
	    RECT 120.6000 168.1000 121.0000 168.2000 ;
	    RECT 133.4000 168.1000 133.8000 168.2000 ;
	    RECT 134.2000 168.1000 134.6000 168.2000 ;
	    RECT 120.6000 167.8000 134.6000 168.1000 ;
	    RECT 173.4000 167.8000 173.8000 168.2000 ;
	    RECT 207.0000 168.1000 207.4000 168.2000 ;
	    RECT 229.4000 168.1000 229.8000 168.2000 ;
	    RECT 257.4000 168.1000 257.8000 168.2000 ;
	    RECT 207.0000 167.8000 257.8000 168.1000 ;
	    RECT 6.2000 167.1000 6.6000 167.2000 ;
	    RECT 11.0000 167.1000 11.4000 167.2000 ;
	    RECT 6.2000 166.8000 11.4000 167.1000 ;
	    RECT 35.8000 167.1000 36.2000 167.2000 ;
	    RECT 42.2000 167.1000 42.6000 167.2000 ;
	    RECT 35.8000 166.8000 42.6000 167.1000 ;
	    RECT 52.6000 167.1000 53.0000 167.2000 ;
	    RECT 55.0000 167.1000 55.4000 167.2000 ;
	    RECT 52.6000 166.8000 55.4000 167.1000 ;
	    RECT 56.6000 167.1000 57.0000 167.2000 ;
	    RECT 61.4000 167.1000 61.8000 167.2000 ;
	    RECT 56.6000 166.8000 61.8000 167.1000 ;
	    RECT 89.4000 167.1000 89.8000 167.2000 ;
	    RECT 97.4000 167.1000 97.8000 167.2000 ;
	    RECT 89.4000 166.8000 97.8000 167.1000 ;
	    RECT 101.4000 166.8000 101.8000 167.2000 ;
	    RECT 103.8000 167.1000 104.2000 167.2000 ;
	    RECT 107.8000 167.1000 108.1000 167.8000 ;
	    RECT 103.8000 166.8000 108.1000 167.1000 ;
	    RECT 127.8000 166.8000 128.2000 167.2000 ;
	    RECT 153.4000 167.1000 153.8000 167.2000 ;
	    RECT 158.2000 167.1000 158.6000 167.2000 ;
	    RECT 173.4000 167.1000 173.7000 167.8000 ;
	    RECT 153.4000 166.8000 173.7000 167.1000 ;
	    RECT 175.0000 166.8000 175.4000 167.2000 ;
	    RECT 210.2000 167.1000 210.6000 167.2000 ;
	    RECT 216.6000 167.1000 217.0000 167.2000 ;
	    RECT 210.2000 166.8000 217.0000 167.1000 ;
	    RECT 227.0000 167.1000 227.4000 167.2000 ;
	    RECT 228.6000 167.1000 229.0000 167.2000 ;
	    RECT 227.0000 166.8000 229.0000 167.1000 ;
	    RECT 231.8000 167.1000 232.2000 167.2000 ;
	    RECT 232.6000 167.1000 233.0000 167.2000 ;
	    RECT 231.8000 166.8000 233.0000 167.1000 ;
	    RECT 236.6000 167.1000 237.0000 167.2000 ;
	    RECT 240.6000 167.1000 241.0000 167.2000 ;
	    RECT 244.6000 167.1000 245.0000 167.2000 ;
	    RECT 249.4000 167.1000 249.8000 167.2000 ;
	    RECT 236.6000 166.8000 249.8000 167.1000 ;
	    RECT 23.8000 166.1000 24.2000 166.2000 ;
	    RECT 25.4000 166.1000 25.8000 166.2000 ;
	    RECT 23.8000 165.8000 25.8000 166.1000 ;
	    RECT 29.4000 166.1000 29.8000 166.2000 ;
	    RECT 32.6000 166.1000 33.0000 166.2000 ;
	    RECT 29.4000 165.8000 33.0000 166.1000 ;
	    RECT 50.2000 166.1000 50.6000 166.2000 ;
	    RECT 53.4000 166.1000 53.8000 166.2000 ;
	    RECT 58.2000 166.1000 58.6000 166.2000 ;
	    RECT 50.2000 165.8000 58.6000 166.1000 ;
	    RECT 71.8000 166.1000 72.2000 166.2000 ;
	    RECT 80.6000 166.1000 81.0000 166.2000 ;
	    RECT 71.8000 165.8000 81.0000 166.1000 ;
	    RECT 82.2000 166.1000 82.6000 166.2000 ;
	    RECT 92.6000 166.1000 93.0000 166.2000 ;
	    RECT 98.2000 166.1000 98.6000 166.2000 ;
	    RECT 82.2000 165.8000 98.6000 166.1000 ;
	    RECT 101.4000 166.1000 101.7000 166.8000 ;
	    RECT 110.2000 166.1000 110.6000 166.3000 ;
	    RECT 101.4000 165.9000 110.6000 166.1000 ;
	    RECT 127.8000 166.1000 128.1000 166.8000 ;
	    RECT 132.6000 166.1000 133.0000 166.2000 ;
	    RECT 101.4000 165.8000 110.5000 165.9000 ;
	    RECT 127.8000 165.8000 133.0000 166.1000 ;
	    RECT 141.4000 166.1000 141.8000 166.2000 ;
	    RECT 147.8000 166.1000 148.2000 166.2000 ;
	    RECT 141.4000 165.8000 148.2000 166.1000 ;
	    RECT 151.8000 166.1000 152.2000 166.2000 ;
	    RECT 159.8000 166.1000 160.2000 166.2000 ;
	    RECT 151.8000 165.8000 160.2000 166.1000 ;
	    RECT 170.2000 166.1000 170.6000 166.2000 ;
	    RECT 175.0000 166.1000 175.3000 166.8000 ;
	    RECT 170.2000 165.8000 175.3000 166.1000 ;
	    RECT 183.8000 166.1000 184.2000 166.2000 ;
	    RECT 191.0000 166.1000 191.4000 166.2000 ;
	    RECT 183.8000 165.8000 191.4000 166.1000 ;
	    RECT 208.6000 166.1000 209.0000 166.2000 ;
	    RECT 214.2000 166.1000 214.6000 166.2000 ;
	    RECT 235.8000 166.1000 236.2000 166.2000 ;
	    RECT 245.4000 166.1000 245.8000 166.2000 ;
	    RECT 208.6000 165.8000 214.6000 166.1000 ;
	    RECT 227.8000 165.8000 230.5000 166.1000 ;
	    RECT 235.8000 165.8000 245.8000 166.1000 ;
	    RECT 246.2000 166.1000 246.6000 166.2000 ;
	    RECT 247.0000 166.1000 247.4000 166.2000 ;
	    RECT 246.2000 165.8000 247.4000 166.1000 ;
	    RECT 247.8000 166.1000 248.2000 166.2000 ;
	    RECT 257.4000 166.1000 257.8000 166.2000 ;
	    RECT 247.8000 165.8000 257.8000 166.1000 ;
	    RECT 227.8000 165.2000 228.1000 165.8000 ;
	    RECT 230.2000 165.2000 230.5000 165.8000 ;
	    RECT 13.4000 164.8000 13.8000 165.2000 ;
	    RECT 38.2000 165.1000 38.6000 165.2000 ;
	    RECT 55.0000 165.1000 55.4000 165.2000 ;
	    RECT 38.2000 164.8000 55.4000 165.1000 ;
	    RECT 62.2000 165.1000 62.6000 165.2000 ;
	    RECT 72.6000 165.1000 73.0000 165.2000 ;
	    RECT 62.2000 164.8000 73.0000 165.1000 ;
	    RECT 91.0000 165.1000 91.4000 165.2000 ;
	    RECT 99.8000 165.1000 100.2000 165.2000 ;
	    RECT 91.0000 164.8000 100.2000 165.1000 ;
	    RECT 158.2000 165.1000 158.6000 165.2000 ;
	    RECT 167.8000 165.1000 168.2000 165.2000 ;
	    RECT 182.2000 165.1000 182.6000 165.2000 ;
	    RECT 158.2000 164.8000 182.6000 165.1000 ;
	    RECT 184.6000 165.1000 185.0000 165.2000 ;
	    RECT 198.2000 165.1000 198.6000 165.2000 ;
	    RECT 184.6000 164.8000 198.6000 165.1000 ;
	    RECT 199.0000 165.1000 199.4000 165.2000 ;
	    RECT 215.8000 165.1000 216.2000 165.2000 ;
	    RECT 223.0000 165.1000 223.4000 165.2000 ;
	    RECT 199.0000 164.8000 223.4000 165.1000 ;
	    RECT 227.8000 164.8000 228.2000 165.2000 ;
	    RECT 230.2000 164.8000 230.6000 165.2000 ;
	    RECT 231.0000 165.1000 231.4000 165.2000 ;
	    RECT 234.2000 165.1000 234.6000 165.2000 ;
	    RECT 237.4000 165.1000 237.8000 165.2000 ;
	    RECT 231.0000 164.8000 234.6000 165.1000 ;
	    RECT 236.6000 164.8000 237.8000 165.1000 ;
	    RECT 238.2000 165.1000 238.6000 165.2000 ;
	    RECT 239.8000 165.1000 240.2000 165.2000 ;
	    RECT 238.2000 164.8000 240.2000 165.1000 ;
	    RECT 240.6000 165.1000 241.0000 165.2000 ;
	    RECT 241.4000 165.1000 241.8000 165.2000 ;
	    RECT 240.6000 164.8000 241.8000 165.1000 ;
	    RECT 10.2000 164.1000 10.6000 164.2000 ;
	    RECT 13.4000 164.1000 13.7000 164.8000 ;
	    RECT 238.2000 164.2000 238.5000 164.8000 ;
	    RECT 10.2000 163.8000 13.7000 164.1000 ;
	    RECT 43.0000 164.1000 43.4000 164.2000 ;
	    RECT 47.8000 164.1000 48.2000 164.2000 ;
	    RECT 43.0000 163.8000 48.2000 164.1000 ;
	    RECT 61.4000 164.1000 61.8000 164.2000 ;
	    RECT 64.6000 164.1000 65.0000 164.2000 ;
	    RECT 68.6000 164.1000 69.0000 164.2000 ;
	    RECT 73.4000 164.1000 73.8000 164.2000 ;
	    RECT 84.6000 164.1000 85.0000 164.2000 ;
	    RECT 102.2000 164.1000 102.6000 164.2000 ;
	    RECT 119.0000 164.1000 119.4000 164.2000 ;
	    RECT 136.6000 164.1000 137.0000 164.2000 ;
	    RECT 138.2000 164.1000 138.6000 164.2000 ;
	    RECT 61.4000 163.8000 138.6000 164.1000 ;
	    RECT 187.8000 164.1000 188.2000 164.2000 ;
	    RECT 203.8000 164.1000 204.2000 164.2000 ;
	    RECT 235.8000 164.1000 236.2000 164.2000 ;
	    RECT 187.8000 163.8000 236.2000 164.1000 ;
	    RECT 238.2000 163.8000 238.6000 164.2000 ;
	    RECT 241.4000 164.1000 241.8000 164.2000 ;
	    RECT 255.0000 164.1000 255.4000 164.2000 ;
	    RECT 259.0000 164.1000 259.4000 164.2000 ;
	    RECT 241.4000 163.8000 259.4000 164.1000 ;
	    RECT 99.0000 163.1000 99.4000 163.2000 ;
	    RECT 126.2000 163.1000 126.6000 163.2000 ;
	    RECT 134.2000 163.1000 134.6000 163.2000 ;
	    RECT 139.8000 163.1000 140.2000 163.2000 ;
	    RECT 99.0000 162.8000 140.2000 163.1000 ;
	    RECT 199.8000 163.1000 200.2000 163.2000 ;
	    RECT 219.8000 163.1000 220.2000 163.2000 ;
	    RECT 199.8000 162.8000 220.2000 163.1000 ;
	    RECT 71.0000 162.1000 71.4000 162.2000 ;
	    RECT 75.0000 162.1000 75.4000 162.2000 ;
	    RECT 71.0000 161.8000 75.4000 162.1000 ;
	    RECT 88.6000 162.1000 89.0000 162.2000 ;
	    RECT 120.6000 162.1000 121.0000 162.2000 ;
	    RECT 88.6000 161.8000 121.0000 162.1000 ;
	    RECT 132.6000 162.1000 133.0000 162.2000 ;
	    RECT 142.2000 162.1000 142.6000 162.2000 ;
	    RECT 132.6000 161.8000 142.6000 162.1000 ;
	    RECT 190.2000 162.1000 190.6000 162.2000 ;
	    RECT 219.0000 162.1000 219.4000 162.2000 ;
	    RECT 190.2000 161.8000 219.4000 162.1000 ;
	    RECT 219.8000 162.1000 220.2000 162.2000 ;
	    RECT 224.6000 162.1000 225.0000 162.2000 ;
	    RECT 229.4000 162.1000 229.8000 162.2000 ;
	    RECT 231.0000 162.1000 231.4000 162.2000 ;
	    RECT 219.8000 161.8000 231.4000 162.1000 ;
	    RECT 243.8000 162.1000 244.2000 162.2000 ;
	    RECT 246.2000 162.1000 246.6000 162.2000 ;
	    RECT 243.8000 161.8000 246.6000 162.1000 ;
	    RECT 193.4000 161.1000 193.8000 161.2000 ;
	    RECT 210.2000 161.1000 210.6000 161.2000 ;
	    RECT 193.4000 160.8000 210.6000 161.1000 ;
	    RECT 229.4000 161.1000 229.8000 161.2000 ;
	    RECT 251.8000 161.1000 252.2000 161.2000 ;
	    RECT 266.2000 161.1000 266.6000 161.2000 ;
	    RECT 267.8000 161.1000 268.2000 161.2000 ;
	    RECT 229.4000 160.8000 268.2000 161.1000 ;
	    RECT 223.0000 160.1000 223.4000 160.2000 ;
	    RECT 255.8000 160.1000 256.2000 160.2000 ;
	    RECT 223.0000 159.8000 256.2000 160.1000 ;
	    RECT 13.4000 159.1000 13.8000 159.2000 ;
	    RECT 16.6000 159.1000 17.0000 159.2000 ;
	    RECT 13.4000 158.8000 17.0000 159.1000 ;
	    RECT 222.2000 159.1000 222.6000 159.2000 ;
	    RECT 233.4000 159.1000 233.8000 159.2000 ;
	    RECT 259.0000 159.1000 259.4000 159.2000 ;
	    RECT 222.2000 158.8000 259.4000 159.1000 ;
	    RECT 26.2000 158.1000 26.6000 158.2000 ;
	    RECT 35.0000 158.1000 35.4000 158.2000 ;
	    RECT 26.2000 157.8000 35.4000 158.1000 ;
	    RECT 47.0000 158.1000 47.4000 158.2000 ;
	    RECT 50.2000 158.1000 50.6000 158.2000 ;
	    RECT 47.0000 157.8000 50.6000 158.1000 ;
	    RECT 195.8000 158.1000 196.2000 158.2000 ;
	    RECT 211.8000 158.1000 212.2000 158.2000 ;
	    RECT 235.0000 158.1000 235.4000 158.2000 ;
	    RECT 195.8000 157.8000 235.4000 158.1000 ;
	    RECT 247.8000 158.1000 248.2000 158.2000 ;
	    RECT 261.4000 158.1000 261.8000 158.2000 ;
	    RECT 247.8000 157.8000 261.8000 158.1000 ;
	    RECT 14.2000 156.8000 14.6000 157.2000 ;
	    RECT 16.6000 157.1000 17.0000 157.2000 ;
	    RECT 20.6000 157.1000 21.0000 157.2000 ;
	    RECT 16.6000 156.8000 21.0000 157.1000 ;
	    RECT 29.4000 157.1000 29.8000 157.2000 ;
	    RECT 35.8000 157.1000 36.2000 157.2000 ;
	    RECT 29.4000 156.8000 36.2000 157.1000 ;
	    RECT 49.4000 156.8000 49.8000 157.2000 ;
	    RECT 101.4000 156.8000 101.8000 157.2000 ;
	    RECT 151.0000 157.1000 151.4000 157.2000 ;
	    RECT 135.8000 156.8000 151.4000 157.1000 ;
	    RECT 159.8000 157.1000 160.2000 157.2000 ;
	    RECT 171.8000 157.1000 172.2000 157.2000 ;
	    RECT 159.8000 156.8000 172.2000 157.1000 ;
	    RECT 191.0000 157.1000 191.4000 157.2000 ;
	    RECT 199.8000 157.1000 200.2000 157.2000 ;
	    RECT 191.0000 156.8000 200.2000 157.1000 ;
	    RECT 217.4000 157.1000 217.8000 157.2000 ;
	    RECT 222.2000 157.1000 222.6000 157.2000 ;
	    RECT 217.4000 156.8000 222.6000 157.1000 ;
	    RECT 249.4000 156.8000 249.8000 157.2000 ;
	    RECT 14.2000 156.2000 14.5000 156.8000 ;
	    RECT 3.8000 156.1000 4.2000 156.2000 ;
	    RECT 4.6000 156.1000 5.0000 156.2000 ;
	    RECT 3.8000 155.8000 5.0000 156.1000 ;
	    RECT 14.2000 155.8000 14.6000 156.2000 ;
	    RECT 29.4000 156.1000 29.8000 156.2000 ;
	    RECT 33.4000 156.1000 33.8000 156.2000 ;
	    RECT 29.4000 155.8000 33.8000 156.1000 ;
	    RECT 35.0000 156.1000 35.4000 156.2000 ;
	    RECT 39.0000 156.1000 39.4000 156.2000 ;
	    RECT 35.0000 155.8000 39.4000 156.1000 ;
	    RECT 49.4000 156.1000 49.7000 156.8000 ;
	    RECT 56.6000 156.1000 57.0000 156.2000 ;
	    RECT 49.4000 155.8000 57.0000 156.1000 ;
	    RECT 64.6000 155.8000 65.0000 156.2000 ;
	    RECT 99.8000 156.1000 100.2000 156.2000 ;
	    RECT 101.4000 156.1000 101.7000 156.8000 ;
	    RECT 135.8000 156.2000 136.1000 156.8000 ;
	    RECT 103.8000 156.1000 104.2000 156.2000 ;
	    RECT 117.4000 156.1000 117.8000 156.2000 ;
	    RECT 99.8000 155.8000 101.7000 156.1000 ;
	    RECT 103.0000 155.8000 117.8000 156.1000 ;
	    RECT 135.8000 155.8000 136.2000 156.2000 ;
	    RECT 140.6000 156.1000 141.0000 156.2000 ;
	    RECT 150.2000 156.1000 150.6000 156.2000 ;
	    RECT 155.0000 156.1000 155.4000 156.2000 ;
	    RECT 140.6000 155.8000 155.4000 156.1000 ;
	    RECT 165.4000 155.8000 165.8000 156.2000 ;
	    RECT 172.6000 156.1000 173.0000 156.2000 ;
	    RECT 179.8000 156.1000 180.2000 156.2000 ;
	    RECT 172.6000 155.8000 180.2000 156.1000 ;
	    RECT 182.2000 156.1000 182.6000 156.2000 ;
	    RECT 183.8000 156.1000 184.2000 156.2000 ;
	    RECT 215.8000 156.1000 216.2000 156.2000 ;
	    RECT 219.8000 156.1000 220.2000 156.2000 ;
	    RECT 182.2000 155.8000 220.2000 156.1000 ;
	    RECT 221.4000 155.8000 228.1000 156.1000 ;
	    RECT 13.4000 155.1000 13.8000 155.2000 ;
	    RECT 14.2000 155.1000 14.6000 155.2000 ;
	    RECT 13.4000 154.8000 14.6000 155.1000 ;
	    RECT 21.4000 155.1000 21.8000 155.2000 ;
	    RECT 24.6000 155.1000 25.0000 155.2000 ;
	    RECT 21.4000 154.8000 25.0000 155.1000 ;
	    RECT 32.6000 155.1000 33.0000 155.2000 ;
	    RECT 36.6000 155.1000 37.0000 155.2000 ;
	    RECT 40.6000 155.1000 41.0000 155.2000 ;
	    RECT 32.6000 154.8000 41.0000 155.1000 ;
	    RECT 50.2000 155.1000 50.6000 155.2000 ;
	    RECT 51.0000 155.1000 51.4000 155.2000 ;
	    RECT 50.2000 154.8000 51.4000 155.1000 ;
	    RECT 63.0000 155.1000 63.4000 155.2000 ;
	    RECT 64.6000 155.1000 64.9000 155.8000 ;
	    RECT 63.0000 154.8000 64.9000 155.1000 ;
	    RECT 133.4000 155.1000 133.8000 155.2000 ;
	    RECT 135.8000 155.1000 136.2000 155.2000 ;
	    RECT 136.6000 155.1000 137.0000 155.2000 ;
	    RECT 165.4000 155.1000 165.7000 155.8000 ;
	    RECT 221.4000 155.2000 221.7000 155.8000 ;
	    RECT 227.8000 155.2000 228.1000 155.8000 ;
	    RECT 236.6000 155.8000 237.0000 156.2000 ;
	    RECT 249.4000 156.1000 249.7000 156.8000 ;
	    RECT 253.4000 156.1000 253.8000 156.2000 ;
	    RECT 249.4000 155.8000 253.8000 156.1000 ;
	    RECT 254.2000 156.1000 254.6000 156.2000 ;
	    RECT 255.8000 156.1000 256.2000 156.2000 ;
	    RECT 254.2000 155.8000 256.2000 156.1000 ;
	    RECT 257.4000 156.1000 257.8000 156.2000 ;
	    RECT 264.6000 156.1000 265.0000 156.2000 ;
	    RECT 269.4000 156.1000 269.8000 156.2000 ;
	    RECT 257.4000 155.8000 269.8000 156.1000 ;
	    RECT 168.6000 155.1000 169.0000 155.2000 ;
	    RECT 133.4000 154.8000 137.0000 155.1000 ;
	    RECT 137.4000 154.8000 145.0000 155.1000 ;
	    RECT 165.4000 154.8000 169.0000 155.1000 ;
	    RECT 173.4000 155.1000 173.8000 155.2000 ;
	    RECT 191.8000 155.1000 192.2000 155.2000 ;
	    RECT 173.4000 154.8000 192.2000 155.1000 ;
	    RECT 193.4000 154.8000 193.8000 155.2000 ;
	    RECT 199.0000 155.1000 199.4000 155.2000 ;
	    RECT 214.2000 155.1000 214.6000 155.2000 ;
	    RECT 219.0000 155.1000 219.4000 155.2000 ;
	    RECT 199.0000 154.8000 204.9000 155.1000 ;
	    RECT 214.2000 154.8000 219.4000 155.1000 ;
	    RECT 221.4000 154.8000 221.8000 155.2000 ;
	    RECT 227.8000 154.8000 228.2000 155.2000 ;
	    RECT 236.6000 155.1000 236.9000 155.8000 ;
	    RECT 246.2000 155.1000 246.6000 155.2000 ;
	    RECT 236.6000 154.8000 246.6000 155.1000 ;
	    RECT 250.2000 155.1000 250.6000 155.2000 ;
	    RECT 254.2000 155.1000 254.6000 155.2000 ;
	    RECT 250.2000 154.8000 254.6000 155.1000 ;
	    RECT 137.4000 154.2000 137.7000 154.8000 ;
	    RECT 144.6000 154.7000 145.0000 154.8000 ;
	    RECT 19.0000 154.1000 19.4000 154.2000 ;
	    RECT 23.8000 154.1000 24.2000 154.2000 ;
	    RECT 27.8000 154.1000 28.2000 154.2000 ;
	    RECT 19.0000 153.8000 28.2000 154.1000 ;
	    RECT 30.2000 154.1000 30.6000 154.2000 ;
	    RECT 38.2000 154.1000 38.6000 154.2000 ;
	    RECT 30.2000 153.8000 38.6000 154.1000 ;
	    RECT 78.2000 154.1000 78.6000 154.2000 ;
	    RECT 86.2000 154.1000 86.6000 154.2000 ;
	    RECT 78.2000 153.8000 86.6000 154.1000 ;
	    RECT 91.0000 154.1000 91.4000 154.2000 ;
	    RECT 135.0000 154.1000 135.4000 154.2000 ;
	    RECT 91.0000 153.8000 135.4000 154.1000 ;
	    RECT 137.4000 153.8000 137.8000 154.2000 ;
	    RECT 142.2000 154.1000 142.6000 154.2000 ;
	    RECT 152.6000 154.1000 153.0000 154.2000 ;
	    RECT 158.2000 154.1000 158.6000 154.2000 ;
	    RECT 142.2000 153.8000 158.6000 154.1000 ;
	    RECT 171.0000 154.1000 171.4000 154.2000 ;
	    RECT 176.6000 154.1000 177.0000 154.2000 ;
	    RECT 171.0000 153.8000 177.0000 154.1000 ;
	    RECT 178.2000 154.1000 178.6000 154.2000 ;
	    RECT 179.8000 154.1000 180.2000 154.2000 ;
	    RECT 178.2000 153.8000 180.2000 154.1000 ;
	    RECT 190.2000 154.1000 190.6000 154.2000 ;
	    RECT 193.4000 154.1000 193.7000 154.8000 ;
	    RECT 204.6000 154.2000 204.9000 154.8000 ;
	    RECT 190.2000 153.8000 193.7000 154.1000 ;
	    RECT 198.2000 154.1000 198.6000 154.2000 ;
	    RECT 199.0000 154.1000 199.4000 154.2000 ;
	    RECT 198.2000 153.8000 199.4000 154.1000 ;
	    RECT 204.6000 153.8000 205.0000 154.2000 ;
	    RECT 218.2000 154.1000 218.6000 154.2000 ;
	    RECT 221.4000 154.1000 221.8000 154.2000 ;
	    RECT 218.2000 153.8000 221.8000 154.1000 ;
	    RECT 259.0000 154.1000 259.4000 154.2000 ;
	    RECT 264.6000 154.1000 265.0000 154.2000 ;
	    RECT 259.0000 153.8000 265.0000 154.1000 ;
	    RECT 25.4000 153.1000 25.8000 153.2000 ;
	    RECT 39.0000 153.1000 39.4000 153.2000 ;
	    RECT 25.4000 152.8000 39.4000 153.1000 ;
	    RECT 41.4000 153.1000 41.8000 153.2000 ;
	    RECT 43.0000 153.1000 43.4000 153.2000 ;
	    RECT 41.4000 152.8000 43.4000 153.1000 ;
	    RECT 75.0000 153.1000 75.4000 153.2000 ;
	    RECT 77.4000 153.1000 77.8000 153.2000 ;
	    RECT 75.0000 152.8000 77.8000 153.1000 ;
	    RECT 95.0000 153.1000 95.4000 153.2000 ;
	    RECT 99.8000 153.1000 100.2000 153.2000 ;
	    RECT 95.0000 152.8000 100.2000 153.1000 ;
	    RECT 100.6000 153.1000 101.0000 153.2000 ;
	    RECT 103.0000 153.1000 103.4000 153.2000 ;
	    RECT 104.6000 153.1000 105.0000 153.2000 ;
	    RECT 100.6000 152.8000 105.0000 153.1000 ;
	    RECT 107.8000 153.1000 108.2000 153.2000 ;
	    RECT 111.8000 153.1000 112.2000 153.2000 ;
	    RECT 107.8000 152.8000 112.2000 153.1000 ;
	    RECT 119.8000 153.1000 120.2000 153.2000 ;
	    RECT 129.4000 153.1000 129.8000 153.2000 ;
	    RECT 147.0000 153.1000 147.4000 153.2000 ;
	    RECT 151.8000 153.1000 152.2000 153.2000 ;
	    RECT 119.8000 152.8000 152.2000 153.1000 ;
	    RECT 169.4000 153.1000 169.8000 153.2000 ;
	    RECT 184.6000 153.1000 185.0000 153.2000 ;
	    RECT 198.2000 153.1000 198.6000 153.2000 ;
	    RECT 205.4000 153.1000 205.8000 153.2000 ;
	    RECT 207.0000 153.1000 207.4000 153.2000 ;
	    RECT 169.4000 152.8000 207.4000 153.1000 ;
	    RECT 213.4000 153.1000 213.8000 153.2000 ;
	    RECT 215.8000 153.1000 216.2000 153.2000 ;
	    RECT 213.4000 152.8000 216.2000 153.1000 ;
	    RECT 229.4000 153.1000 229.8000 153.2000 ;
	    RECT 232.6000 153.1000 233.0000 153.2000 ;
	    RECT 229.4000 152.8000 233.0000 153.1000 ;
	    RECT 241.4000 153.1000 241.8000 153.2000 ;
	    RECT 243.0000 153.1000 243.4000 153.2000 ;
	    RECT 241.4000 152.8000 243.4000 153.1000 ;
	    RECT 251.0000 152.8000 251.4000 153.2000 ;
	    RECT 252.6000 153.1000 253.0000 153.2000 ;
	    RECT 260.6000 153.1000 261.0000 153.2000 ;
	    RECT 252.6000 152.8000 261.0000 153.1000 ;
	    RECT 251.0000 152.2000 251.3000 152.8000 ;
	    RECT 3.0000 152.1000 3.4000 152.2000 ;
	    RECT 15.8000 152.1000 16.2000 152.2000 ;
	    RECT 3.0000 151.8000 16.2000 152.1000 ;
	    RECT 60.6000 152.1000 61.0000 152.2000 ;
	    RECT 70.2000 152.1000 70.6000 152.2000 ;
	    RECT 60.6000 151.8000 70.6000 152.1000 ;
	    RECT 98.2000 152.1000 98.6000 152.2000 ;
	    RECT 106.2000 152.1000 106.6000 152.2000 ;
	    RECT 108.6000 152.1000 109.0000 152.2000 ;
	    RECT 98.2000 151.8000 109.0000 152.1000 ;
	    RECT 133.4000 152.1000 133.8000 152.2000 ;
	    RECT 136.6000 152.1000 137.0000 152.2000 ;
	    RECT 133.4000 151.8000 137.0000 152.1000 ;
	    RECT 173.4000 152.1000 173.8000 152.2000 ;
	    RECT 176.6000 152.1000 177.0000 152.2000 ;
	    RECT 173.4000 151.8000 177.0000 152.1000 ;
	    RECT 179.8000 152.1000 180.2000 152.2000 ;
	    RECT 182.2000 152.1000 182.6000 152.2000 ;
	    RECT 179.8000 151.8000 182.6000 152.1000 ;
	    RECT 189.4000 152.1000 189.8000 152.2000 ;
	    RECT 191.8000 152.1000 192.2000 152.2000 ;
	    RECT 189.4000 151.8000 192.2000 152.1000 ;
	    RECT 227.0000 152.1000 227.4000 152.2000 ;
	    RECT 250.2000 152.1000 250.6000 152.2000 ;
	    RECT 227.0000 151.8000 250.6000 152.1000 ;
	    RECT 251.0000 151.8000 251.4000 152.2000 ;
	    RECT 254.2000 152.1000 254.6000 152.2000 ;
	    RECT 262.2000 152.1000 262.6000 152.2000 ;
	    RECT 254.2000 151.8000 262.6000 152.1000 ;
	    RECT 127.0000 151.1000 127.4000 151.2000 ;
	    RECT 139.8000 151.1000 140.2000 151.2000 ;
	    RECT 127.0000 150.8000 140.2000 151.1000 ;
	    RECT 175.0000 151.1000 175.4000 151.2000 ;
	    RECT 178.2000 151.1000 178.6000 151.2000 ;
	    RECT 193.4000 151.1000 193.8000 151.2000 ;
	    RECT 199.8000 151.1000 200.2000 151.2000 ;
	    RECT 175.0000 150.8000 200.2000 151.1000 ;
	    RECT 238.2000 151.1000 238.6000 151.2000 ;
	    RECT 239.0000 151.1000 239.4000 151.2000 ;
	    RECT 238.2000 150.8000 239.4000 151.1000 ;
	    RECT 250.2000 151.1000 250.6000 151.2000 ;
	    RECT 251.8000 151.1000 252.2000 151.2000 ;
	    RECT 250.2000 150.8000 252.2000 151.1000 ;
	    RECT 5.4000 150.1000 5.8000 150.2000 ;
	    RECT 24.6000 150.1000 25.0000 150.2000 ;
	    RECT 5.4000 149.8000 25.0000 150.1000 ;
	    RECT 43.8000 150.1000 44.2000 150.2000 ;
	    RECT 53.4000 150.1000 53.8000 150.2000 ;
	    RECT 43.8000 149.8000 53.8000 150.1000 ;
	    RECT 111.8000 150.1000 112.2000 150.2000 ;
	    RECT 115.0000 150.1000 115.4000 150.2000 ;
	    RECT 111.8000 149.8000 115.4000 150.1000 ;
	    RECT 181.4000 150.1000 181.8000 150.2000 ;
	    RECT 187.8000 150.1000 188.2000 150.2000 ;
	    RECT 181.4000 149.8000 188.2000 150.1000 ;
	    RECT 218.2000 150.1000 218.6000 150.2000 ;
	    RECT 224.6000 150.1000 225.0000 150.2000 ;
	    RECT 218.2000 149.8000 225.0000 150.1000 ;
	    RECT 235.8000 150.1000 236.2000 150.2000 ;
	    RECT 239.0000 150.1000 239.4000 150.2000 ;
	    RECT 242.2000 150.1000 242.6000 150.2000 ;
	    RECT 244.6000 150.1000 245.0000 150.2000 ;
	    RECT 249.4000 150.1000 249.8000 150.2000 ;
	    RECT 254.2000 150.1000 254.6000 150.2000 ;
	    RECT 235.8000 149.8000 254.6000 150.1000 ;
	    RECT 261.4000 150.1000 261.8000 150.2000 ;
	    RECT 263.8000 150.1000 264.2000 150.2000 ;
	    RECT 261.4000 149.8000 264.2000 150.1000 ;
	    RECT 0.6000 149.1000 1.0000 149.2000 ;
	    RECT 8.6000 149.1000 9.0000 149.2000 ;
	    RECT 0.6000 148.8000 9.0000 149.1000 ;
	    RECT 10.2000 149.1000 10.6000 149.2000 ;
	    RECT 16.6000 149.1000 17.0000 149.2000 ;
	    RECT 10.2000 148.8000 17.0000 149.1000 ;
	    RECT 29.4000 148.8000 29.8000 149.2000 ;
	    RECT 43.8000 148.8000 44.2000 149.2000 ;
	    RECT 51.8000 149.1000 52.2000 149.2000 ;
	    RECT 67.8000 149.1000 68.2000 149.2000 ;
	    RECT 51.0000 148.8000 68.2000 149.1000 ;
	    RECT 72.6000 149.1000 73.0000 149.2000 ;
	    RECT 85.4000 149.1000 85.8000 149.2000 ;
	    RECT 72.6000 148.8000 85.8000 149.1000 ;
	    RECT 93.4000 149.1000 93.8000 149.2000 ;
	    RECT 94.2000 149.1000 94.6000 149.2000 ;
	    RECT 93.4000 148.8000 94.6000 149.1000 ;
	    RECT 99.8000 149.1000 100.2000 149.2000 ;
	    RECT 111.8000 149.1000 112.2000 149.2000 ;
	    RECT 99.8000 148.8000 112.2000 149.1000 ;
	    RECT 180.6000 149.1000 181.0000 149.2000 ;
	    RECT 182.2000 149.1000 182.6000 149.2000 ;
	    RECT 180.6000 148.8000 182.6000 149.1000 ;
	    RECT 183.8000 149.1000 184.2000 149.2000 ;
	    RECT 185.4000 149.1000 185.8000 149.2000 ;
	    RECT 183.8000 148.8000 185.8000 149.1000 ;
	    RECT 186.2000 148.8000 186.6000 149.2000 ;
	    RECT 198.2000 149.1000 198.6000 149.2000 ;
	    RECT 214.2000 149.1000 214.6000 149.2000 ;
	    RECT 198.2000 148.8000 214.6000 149.1000 ;
	    RECT 223.0000 149.1000 223.4000 149.2000 ;
	    RECT 226.2000 149.1000 226.6000 149.2000 ;
	    RECT 228.6000 149.1000 229.0000 149.2000 ;
	    RECT 223.0000 148.8000 229.0000 149.1000 ;
	    RECT 230.2000 149.1000 230.6000 149.2000 ;
	    RECT 248.6000 149.1000 249.0000 149.2000 ;
	    RECT 230.2000 148.8000 249.0000 149.1000 ;
	    RECT 251.0000 149.1000 251.4000 149.2000 ;
	    RECT 253.4000 149.1000 253.8000 149.2000 ;
	    RECT 251.0000 148.8000 253.8000 149.1000 ;
	    RECT 263.8000 149.1000 264.2000 149.2000 ;
	    RECT 268.6000 149.1000 269.0000 149.2000 ;
	    RECT 263.8000 148.8000 269.7000 149.1000 ;
	    RECT 270.2000 148.8000 270.6000 149.2000 ;
	    RECT 29.4000 148.2000 29.7000 148.8000 ;
	    RECT 18.2000 148.1000 18.6000 148.2000 ;
	    RECT 23.8000 148.1000 24.2000 148.2000 ;
	    RECT 18.2000 147.8000 24.2000 148.1000 ;
	    RECT 27.8000 147.8000 28.2000 148.2000 ;
	    RECT 29.4000 147.8000 29.8000 148.2000 ;
	    RECT 43.8000 148.1000 44.1000 148.8000 ;
	    RECT 50.2000 148.1000 50.6000 148.2000 ;
	    RECT 43.8000 147.8000 50.6000 148.1000 ;
	    RECT 63.0000 148.1000 63.4000 148.2000 ;
	    RECT 67.0000 148.1000 67.4000 148.2000 ;
	    RECT 63.0000 147.8000 67.4000 148.1000 ;
	    RECT 82.2000 147.8000 82.6000 148.2000 ;
	    RECT 87.0000 147.8000 87.4000 148.2000 ;
	    RECT 104.6000 148.1000 105.0000 148.2000 ;
	    RECT 109.4000 148.1000 109.8000 148.2000 ;
	    RECT 104.6000 147.8000 109.8000 148.1000 ;
	    RECT 112.6000 148.1000 113.0000 148.2000 ;
	    RECT 120.6000 148.1000 121.0000 148.2000 ;
	    RECT 122.2000 148.1000 122.6000 148.2000 ;
	    RECT 112.6000 147.8000 122.6000 148.1000 ;
	    RECT 171.0000 148.1000 171.4000 148.2000 ;
	    RECT 172.6000 148.1000 173.0000 148.2000 ;
	    RECT 180.6000 148.1000 181.0000 148.2000 ;
	    RECT 186.2000 148.1000 186.5000 148.8000 ;
	    RECT 171.0000 147.8000 186.5000 148.1000 ;
	    RECT 203.8000 148.1000 204.2000 148.2000 ;
	    RECT 208.6000 148.1000 209.0000 148.2000 ;
	    RECT 203.8000 147.8000 209.0000 148.1000 ;
	    RECT 211.8000 148.1000 212.2000 148.2000 ;
	    RECT 215.8000 148.1000 216.2000 148.2000 ;
	    RECT 257.4000 148.1000 257.8000 148.2000 ;
	    RECT 258.2000 148.1000 258.6000 148.2000 ;
	    RECT 211.8000 147.8000 258.6000 148.1000 ;
	    RECT 268.6000 148.1000 269.0000 148.2000 ;
	    RECT 270.2000 148.1000 270.5000 148.8000 ;
	    RECT 268.6000 147.8000 270.5000 148.1000 ;
	    RECT 21.4000 146.8000 21.8000 147.2000 ;
	    RECT 23.0000 147.1000 23.4000 147.2000 ;
	    RECT 27.8000 147.1000 28.1000 147.8000 ;
	    RECT 23.0000 146.8000 28.1000 147.1000 ;
	    RECT 43.8000 147.1000 44.2000 147.2000 ;
	    RECT 57.4000 147.1000 57.8000 147.2000 ;
	    RECT 63.0000 147.1000 63.4000 147.2000 ;
	    RECT 43.8000 146.8000 63.4000 147.1000 ;
	    RECT 77.4000 146.8000 77.8000 147.2000 ;
	    RECT 82.2000 147.1000 82.5000 147.8000 ;
	    RECT 87.0000 147.1000 87.3000 147.8000 ;
	    RECT 82.2000 146.8000 87.3000 147.1000 ;
	    RECT 95.0000 147.1000 95.4000 147.2000 ;
	    RECT 99.8000 147.1000 100.2000 147.2000 ;
	    RECT 95.0000 146.8000 100.2000 147.1000 ;
	    RECT 110.2000 147.1000 110.6000 147.2000 ;
	    RECT 119.0000 147.1000 119.4000 147.2000 ;
	    RECT 119.8000 147.1000 120.2000 147.2000 ;
	    RECT 110.2000 146.8000 120.2000 147.1000 ;
	    RECT 135.0000 147.1000 135.4000 147.2000 ;
	    RECT 138.2000 147.1000 138.6000 147.2000 ;
	    RECT 143.8000 147.1000 144.2000 147.2000 ;
	    RECT 153.4000 147.1000 153.8000 147.2000 ;
	    RECT 135.0000 146.8000 153.8000 147.1000 ;
	    RECT 179.0000 147.1000 179.4000 147.2000 ;
	    RECT 186.2000 147.1000 186.6000 147.2000 ;
	    RECT 188.6000 147.1000 189.0000 147.2000 ;
	    RECT 179.0000 146.8000 185.7000 147.1000 ;
	    RECT 186.2000 146.8000 189.0000 147.1000 ;
	    RECT 191.0000 147.1000 191.4000 147.2000 ;
	    RECT 212.6000 147.1000 213.0000 147.2000 ;
	    RECT 213.4000 147.1000 213.8000 147.2000 ;
	    RECT 191.0000 146.8000 212.1000 147.1000 ;
	    RECT 212.6000 146.8000 213.8000 147.1000 ;
	    RECT 214.2000 147.1000 214.6000 147.2000 ;
	    RECT 225.4000 147.1000 225.8000 147.2000 ;
	    RECT 214.2000 146.8000 225.8000 147.1000 ;
	    RECT 229.4000 147.1000 229.8000 147.2000 ;
	    RECT 239.8000 147.1000 240.2000 147.2000 ;
	    RECT 229.4000 146.8000 240.2000 147.1000 ;
	    RECT 242.2000 147.1000 242.6000 147.2000 ;
	    RECT 243.0000 147.1000 243.4000 147.2000 ;
	    RECT 242.2000 146.8000 243.4000 147.1000 ;
	    RECT 244.6000 147.1000 245.0000 147.2000 ;
	    RECT 253.4000 147.1000 253.8000 147.2000 ;
	    RECT 244.6000 146.8000 253.8000 147.1000 ;
	    RECT 254.2000 147.1000 254.6000 147.2000 ;
	    RECT 259.0000 147.1000 259.4000 147.2000 ;
	    RECT 254.2000 146.8000 259.4000 147.1000 ;
	    RECT 263.0000 147.1000 263.4000 147.2000 ;
	    RECT 264.6000 147.1000 265.0000 147.2000 ;
	    RECT 263.0000 146.8000 265.0000 147.1000 ;
	    RECT 3.8000 146.1000 4.2000 146.2000 ;
	    RECT 4.6000 146.1000 5.0000 146.2000 ;
	    RECT 3.8000 145.8000 5.0000 146.1000 ;
	    RECT 7.8000 146.1000 8.2000 146.2000 ;
	    RECT 21.4000 146.1000 21.7000 146.8000 ;
	    RECT 7.8000 145.8000 21.7000 146.1000 ;
	    RECT 51.0000 146.1000 51.4000 146.2000 ;
	    RECT 55.8000 146.1000 56.2000 146.2000 ;
	    RECT 51.0000 145.8000 56.2000 146.1000 ;
	    RECT 69.4000 146.1000 69.8000 146.2000 ;
	    RECT 77.4000 146.1000 77.7000 146.8000 ;
	    RECT 69.4000 145.8000 77.7000 146.1000 ;
	    RECT 83.8000 146.1000 84.2000 146.2000 ;
	    RECT 87.0000 146.1000 87.4000 146.2000 ;
	    RECT 83.8000 145.8000 87.4000 146.1000 ;
	    RECT 88.6000 146.1000 89.0000 146.2000 ;
	    RECT 95.8000 146.1000 96.2000 146.2000 ;
	    RECT 88.6000 145.8000 96.2000 146.1000 ;
	    RECT 104.6000 146.1000 105.0000 146.2000 ;
	    RECT 107.0000 146.1000 107.4000 146.2000 ;
	    RECT 104.6000 145.8000 107.4000 146.1000 ;
	    RECT 115.0000 146.1000 115.4000 146.2000 ;
	    RECT 117.4000 146.1000 117.8000 146.2000 ;
	    RECT 115.0000 145.8000 117.8000 146.1000 ;
	    RECT 140.6000 146.1000 141.0000 146.2000 ;
	    RECT 141.4000 146.1000 141.8000 146.2000 ;
	    RECT 140.6000 145.8000 141.8000 146.1000 ;
	    RECT 142.2000 146.1000 142.6000 146.2000 ;
	    RECT 143.0000 146.1000 143.4000 146.2000 ;
	    RECT 144.6000 146.1000 145.0000 146.2000 ;
	    RECT 152.6000 146.1000 153.0000 146.2000 ;
	    RECT 142.2000 145.8000 143.4000 146.1000 ;
	    RECT 143.8000 145.8000 153.0000 146.1000 ;
	    RECT 166.2000 146.1000 166.6000 146.2000 ;
	    RECT 173.4000 146.1000 173.8000 146.2000 ;
	    RECT 166.2000 145.8000 173.8000 146.1000 ;
	    RECT 181.4000 146.1000 181.8000 146.2000 ;
	    RECT 183.0000 146.1000 183.4000 146.2000 ;
	    RECT 181.4000 145.8000 183.4000 146.1000 ;
	    RECT 185.4000 146.1000 185.7000 146.8000 ;
	    RECT 188.6000 146.1000 189.0000 146.2000 ;
	    RECT 185.4000 145.8000 189.0000 146.1000 ;
	    RECT 191.8000 146.1000 192.2000 146.2000 ;
	    RECT 195.8000 146.1000 196.2000 146.2000 ;
	    RECT 208.6000 146.1000 209.0000 146.2000 ;
	    RECT 191.8000 145.8000 194.5000 146.1000 ;
	    RECT 195.8000 145.8000 209.0000 146.1000 ;
	    RECT 211.8000 146.1000 212.1000 146.8000 ;
	    RECT 220.6000 146.1000 221.0000 146.2000 ;
	    RECT 211.8000 145.8000 221.0000 146.1000 ;
	    RECT 221.4000 146.1000 221.8000 146.2000 ;
	    RECT 223.8000 146.1000 224.2000 146.2000 ;
	    RECT 231.8000 146.1000 232.2000 146.2000 ;
	    RECT 233.4000 146.1000 233.8000 146.2000 ;
	    RECT 221.4000 145.8000 228.9000 146.1000 ;
	    RECT 231.8000 145.8000 233.8000 146.1000 ;
	    RECT 239.0000 146.1000 239.4000 146.2000 ;
	    RECT 240.6000 146.1000 241.0000 146.2000 ;
	    RECT 239.0000 145.8000 241.0000 146.1000 ;
	    RECT 242.2000 146.1000 242.6000 146.2000 ;
	    RECT 251.0000 146.1000 251.4000 146.2000 ;
	    RECT 252.6000 146.1000 253.0000 146.2000 ;
	    RECT 242.2000 145.8000 253.0000 146.1000 ;
	    RECT 258.2000 146.1000 258.6000 146.2000 ;
	    RECT 261.4000 146.1000 261.8000 146.2000 ;
	    RECT 265.4000 146.1000 265.8000 146.2000 ;
	    RECT 268.6000 146.1000 269.0000 146.2000 ;
	    RECT 258.2000 145.8000 269.0000 146.1000 ;
	    RECT 194.2000 145.2000 194.5000 145.8000 ;
	    RECT 228.6000 145.2000 228.9000 145.8000 ;
	    RECT 6.2000 145.1000 6.6000 145.2000 ;
	    RECT 7.8000 145.1000 8.2000 145.2000 ;
	    RECT 6.2000 144.8000 8.2000 145.1000 ;
	    RECT 9.4000 145.1000 9.8000 145.2000 ;
	    RECT 11.0000 145.1000 11.4000 145.2000 ;
	    RECT 9.4000 144.8000 11.4000 145.1000 ;
	    RECT 14.2000 145.1000 14.6000 145.2000 ;
	    RECT 17.4000 145.1000 17.8000 145.2000 ;
	    RECT 14.2000 144.8000 17.8000 145.1000 ;
	    RECT 54.2000 145.1000 54.6000 145.2000 ;
	    RECT 72.6000 145.1000 73.0000 145.2000 ;
	    RECT 54.2000 144.8000 73.0000 145.1000 ;
	    RECT 83.8000 144.8000 84.2000 145.2000 ;
	    RECT 85.4000 145.1000 85.8000 145.2000 ;
	    RECT 97.4000 145.1000 97.8000 145.2000 ;
	    RECT 103.8000 145.1000 104.2000 145.2000 ;
	    RECT 85.4000 144.8000 104.2000 145.1000 ;
	    RECT 112.6000 145.1000 113.0000 145.2000 ;
	    RECT 127.8000 145.1000 128.2000 145.2000 ;
	    RECT 112.6000 144.8000 128.2000 145.1000 ;
	    RECT 159.8000 145.1000 160.2000 145.2000 ;
	    RECT 179.0000 145.1000 179.4000 145.2000 ;
	    RECT 159.8000 144.8000 179.4000 145.1000 ;
	    RECT 187.8000 145.1000 188.2000 145.2000 ;
	    RECT 189.4000 145.1000 189.8000 145.2000 ;
	    RECT 187.8000 144.8000 189.8000 145.1000 ;
	    RECT 194.2000 144.8000 194.6000 145.2000 ;
	    RECT 216.6000 145.1000 217.0000 145.2000 ;
	    RECT 223.8000 145.1000 224.2000 145.2000 ;
	    RECT 195.0000 144.8000 224.2000 145.1000 ;
	    RECT 224.6000 145.1000 225.0000 145.2000 ;
	    RECT 227.8000 145.1000 228.2000 145.2000 ;
	    RECT 224.6000 144.8000 228.2000 145.1000 ;
	    RECT 228.6000 144.8000 229.0000 145.2000 ;
	    RECT 230.2000 145.1000 230.6000 145.2000 ;
	    RECT 234.2000 145.1000 234.6000 145.2000 ;
	    RECT 230.2000 144.8000 234.6000 145.1000 ;
	    RECT 240.6000 145.1000 241.0000 145.2000 ;
	    RECT 243.0000 145.1000 243.4000 145.2000 ;
	    RECT 240.6000 144.8000 243.4000 145.1000 ;
	    RECT 251.0000 144.8000 251.4000 145.2000 ;
	    RECT 251.8000 145.1000 252.2000 145.2000 ;
	    RECT 255.0000 145.1000 255.4000 145.2000 ;
	    RECT 251.8000 144.8000 255.4000 145.1000 ;
	    RECT 35.8000 144.1000 36.2000 144.2000 ;
	    RECT 40.6000 144.1000 41.0000 144.2000 ;
	    RECT 35.8000 143.8000 41.0000 144.1000 ;
	    RECT 46.2000 144.1000 46.6000 144.2000 ;
	    RECT 55.0000 144.1000 55.4000 144.2000 ;
	    RECT 62.2000 144.1000 62.6000 144.2000 ;
	    RECT 46.2000 143.8000 62.6000 144.1000 ;
	    RECT 74.2000 144.1000 74.6000 144.2000 ;
	    RECT 83.8000 144.1000 84.1000 144.8000 ;
	    RECT 74.2000 143.8000 84.1000 144.1000 ;
	    RECT 88.6000 144.1000 89.0000 144.2000 ;
	    RECT 90.2000 144.1000 90.6000 144.2000 ;
	    RECT 116.6000 144.1000 117.0000 144.2000 ;
	    RECT 88.6000 143.8000 117.0000 144.1000 ;
	    RECT 177.4000 144.1000 177.8000 144.2000 ;
	    RECT 180.6000 144.1000 181.0000 144.2000 ;
	    RECT 190.2000 144.1000 190.6000 144.2000 ;
	    RECT 177.4000 143.8000 190.6000 144.1000 ;
	    RECT 191.0000 144.1000 191.4000 144.2000 ;
	    RECT 195.0000 144.1000 195.3000 144.8000 ;
	    RECT 191.0000 143.8000 195.3000 144.1000 ;
	    RECT 216.6000 144.1000 217.0000 144.2000 ;
	    RECT 227.0000 144.1000 227.4000 144.2000 ;
	    RECT 216.6000 143.8000 227.4000 144.1000 ;
	    RECT 227.8000 144.1000 228.2000 144.2000 ;
	    RECT 237.4000 144.1000 237.8000 144.2000 ;
	    RECT 227.8000 143.8000 237.8000 144.1000 ;
	    RECT 246.2000 144.1000 246.6000 144.2000 ;
	    RECT 251.0000 144.1000 251.3000 144.8000 ;
	    RECT 246.2000 143.8000 251.3000 144.1000 ;
	    RECT 118.2000 143.1000 118.6000 143.2000 ;
	    RECT 128.6000 143.1000 129.0000 143.2000 ;
	    RECT 118.2000 142.8000 129.0000 143.1000 ;
	    RECT 192.6000 143.1000 193.0000 143.2000 ;
	    RECT 210.2000 143.1000 210.6000 143.2000 ;
	    RECT 192.6000 142.8000 210.6000 143.1000 ;
	    RECT 244.6000 142.8000 245.0000 143.2000 ;
	    RECT 87.0000 142.1000 87.4000 142.2000 ;
	    RECT 159.8000 142.1000 160.2000 142.2000 ;
	    RECT 87.0000 141.8000 160.2000 142.1000 ;
	    RECT 163.8000 142.1000 164.2000 142.2000 ;
	    RECT 175.8000 142.1000 176.2000 142.2000 ;
	    RECT 163.8000 141.8000 176.2000 142.1000 ;
	    RECT 186.2000 142.1000 186.6000 142.2000 ;
	    RECT 200.6000 142.1000 201.0000 142.2000 ;
	    RECT 186.2000 141.8000 201.0000 142.1000 ;
	    RECT 214.2000 142.1000 214.6000 142.2000 ;
	    RECT 244.6000 142.1000 244.9000 142.8000 ;
	    RECT 214.2000 141.8000 244.9000 142.1000 ;
	    RECT 258.2000 142.1000 258.6000 142.2000 ;
	    RECT 261.4000 142.1000 261.8000 142.2000 ;
	    RECT 258.2000 141.8000 261.8000 142.1000 ;
	    RECT 39.0000 140.8000 39.4000 141.2000 ;
	    RECT 201.4000 141.1000 201.8000 141.2000 ;
	    RECT 242.2000 141.1000 242.6000 141.2000 ;
	    RECT 201.4000 140.8000 242.6000 141.1000 ;
	    RECT 39.0000 140.2000 39.3000 140.8000 ;
	    RECT 39.0000 139.8000 39.4000 140.2000 ;
	    RECT 135.8000 140.1000 136.2000 140.2000 ;
	    RECT 143.8000 140.1000 144.2000 140.2000 ;
	    RECT 135.8000 139.8000 144.2000 140.1000 ;
	    RECT 175.8000 140.1000 176.2000 140.2000 ;
	    RECT 176.6000 140.1000 177.0000 140.2000 ;
	    RECT 175.8000 139.8000 177.0000 140.1000 ;
	    RECT 187.0000 140.1000 187.4000 140.2000 ;
	    RECT 202.2000 140.1000 202.6000 140.2000 ;
	    RECT 187.0000 139.8000 202.6000 140.1000 ;
	    RECT 256.6000 140.1000 257.0000 140.2000 ;
	    RECT 262.2000 140.1000 262.6000 140.2000 ;
	    RECT 256.6000 139.8000 262.6000 140.1000 ;
	    RECT 26.2000 139.1000 26.6000 139.2000 ;
	    RECT 34.2000 139.1000 34.6000 139.2000 ;
	    RECT 26.2000 138.8000 34.6000 139.1000 ;
	    RECT 38.2000 139.1000 38.6000 139.2000 ;
	    RECT 50.2000 139.1000 50.6000 139.2000 ;
	    RECT 86.2000 139.1000 86.6000 139.2000 ;
	    RECT 38.2000 138.8000 86.6000 139.1000 ;
	    RECT 123.0000 139.1000 123.4000 139.2000 ;
	    RECT 131.8000 139.1000 132.2000 139.2000 ;
	    RECT 137.4000 139.1000 137.8000 139.2000 ;
	    RECT 123.0000 138.8000 137.8000 139.1000 ;
	    RECT 175.8000 139.1000 176.2000 139.2000 ;
	    RECT 200.6000 139.1000 201.0000 139.2000 ;
	    RECT 207.8000 139.1000 208.2000 139.2000 ;
	    RECT 224.6000 139.1000 225.0000 139.2000 ;
	    RECT 241.4000 139.1000 241.8000 139.2000 ;
	    RECT 175.8000 138.8000 208.2000 139.1000 ;
	    RECT 219.0000 138.8000 241.8000 139.1000 ;
	    RECT 242.2000 139.1000 242.6000 139.2000 ;
	    RECT 266.2000 139.1000 266.6000 139.2000 ;
	    RECT 242.2000 138.8000 266.6000 139.1000 ;
	    RECT 219.0000 138.2000 219.3000 138.8000 ;
	    RECT 1.4000 138.1000 1.8000 138.2000 ;
	    RECT 28.6000 138.1000 29.0000 138.2000 ;
	    RECT 31.0000 138.1000 31.4000 138.2000 ;
	    RECT 1.4000 137.8000 31.4000 138.1000 ;
	    RECT 83.8000 138.1000 84.2000 138.2000 ;
	    RECT 87.8000 138.1000 88.2000 138.2000 ;
	    RECT 83.8000 137.8000 88.2000 138.1000 ;
	    RECT 107.8000 138.1000 108.2000 138.2000 ;
	    RECT 118.2000 138.1000 118.6000 138.2000 ;
	    RECT 107.8000 137.8000 118.6000 138.1000 ;
	    RECT 195.0000 138.1000 195.4000 138.2000 ;
	    RECT 201.4000 138.1000 201.8000 138.2000 ;
	    RECT 195.0000 137.8000 201.8000 138.1000 ;
	    RECT 219.0000 137.8000 219.4000 138.2000 ;
	    RECT 237.4000 138.1000 237.8000 138.2000 ;
	    RECT 255.0000 138.1000 255.4000 138.2000 ;
	    RECT 258.2000 138.1000 258.6000 138.2000 ;
	    RECT 237.4000 137.8000 258.6000 138.1000 ;
	    RECT 259.0000 137.8000 259.4000 138.2000 ;
	    RECT 16.6000 137.1000 17.0000 137.2000 ;
	    RECT 25.4000 137.1000 25.8000 137.2000 ;
	    RECT 16.6000 136.8000 25.8000 137.1000 ;
	    RECT 27.0000 136.8000 27.4000 137.2000 ;
	    RECT 50.2000 136.8000 50.6000 137.2000 ;
	    RECT 177.4000 137.1000 177.8000 137.2000 ;
	    RECT 178.2000 137.1000 178.6000 137.2000 ;
	    RECT 194.2000 137.1000 194.6000 137.2000 ;
	    RECT 177.4000 136.8000 194.6000 137.1000 ;
	    RECT 199.0000 137.1000 199.4000 137.2000 ;
	    RECT 199.8000 137.1000 200.2000 137.2000 ;
	    RECT 199.0000 136.8000 200.2000 137.1000 ;
	    RECT 206.2000 136.8000 206.6000 137.2000 ;
	    RECT 210.2000 137.1000 210.6000 137.2000 ;
	    RECT 219.8000 137.1000 220.2000 137.2000 ;
	    RECT 210.2000 136.8000 220.2000 137.1000 ;
	    RECT 228.6000 137.1000 229.0000 137.2000 ;
	    RECT 233.4000 137.1000 233.8000 137.2000 ;
	    RECT 228.6000 136.8000 233.8000 137.1000 ;
	    RECT 235.0000 137.1000 235.4000 137.2000 ;
	    RECT 241.4000 137.1000 241.8000 137.2000 ;
	    RECT 247.0000 137.1000 247.4000 137.2000 ;
	    RECT 247.8000 137.1000 248.2000 137.2000 ;
	    RECT 235.0000 136.8000 248.2000 137.1000 ;
	    RECT 249.4000 137.1000 249.8000 137.2000 ;
	    RECT 259.0000 137.1000 259.3000 137.8000 ;
	    RECT 249.4000 136.8000 259.3000 137.1000 ;
	    RECT 27.0000 136.2000 27.3000 136.8000 ;
	    RECT 15.0000 136.1000 15.4000 136.2000 ;
	    RECT 15.8000 136.1000 16.2000 136.2000 ;
	    RECT 17.4000 136.1000 17.8000 136.2000 ;
	    RECT 19.0000 136.1000 19.4000 136.2000 ;
	    RECT 15.0000 135.8000 19.4000 136.1000 ;
	    RECT 27.0000 135.8000 27.4000 136.2000 ;
	    RECT 29.4000 136.1000 29.8000 136.2000 ;
	    RECT 33.4000 136.1000 33.8000 136.2000 ;
	    RECT 29.4000 135.8000 33.8000 136.1000 ;
	    RECT 42.2000 135.8000 42.6000 136.2000 ;
	    RECT 50.2000 136.1000 50.5000 136.8000 ;
	    RECT 55.8000 136.1000 56.2000 136.2000 ;
	    RECT 50.2000 135.8000 56.2000 136.1000 ;
	    RECT 100.6000 136.1000 101.0000 136.2000 ;
	    RECT 103.0000 136.1000 103.4000 136.2000 ;
	    RECT 112.6000 136.1000 113.0000 136.2000 ;
	    RECT 100.6000 135.8000 113.0000 136.1000 ;
	    RECT 169.4000 136.1000 169.8000 136.2000 ;
	    RECT 176.6000 136.1000 177.0000 136.2000 ;
	    RECT 195.8000 136.1000 196.2000 136.2000 ;
	    RECT 203.8000 136.1000 204.2000 136.2000 ;
	    RECT 169.4000 135.8000 204.2000 136.1000 ;
	    RECT 206.2000 136.1000 206.5000 136.8000 ;
	    RECT 228.6000 136.1000 228.9000 136.8000 ;
	    RECT 206.2000 135.8000 228.9000 136.1000 ;
	    RECT 232.6000 136.1000 233.0000 136.2000 ;
	    RECT 240.6000 136.1000 241.0000 136.2000 ;
	    RECT 241.4000 136.1000 241.8000 136.2000 ;
	    RECT 246.2000 136.1000 246.6000 136.2000 ;
	    RECT 251.0000 136.1000 251.4000 136.2000 ;
	    RECT 232.6000 135.8000 241.8000 136.1000 ;
	    RECT 245.4000 135.8000 251.4000 136.1000 ;
	    RECT 258.2000 136.1000 258.6000 136.2000 ;
	    RECT 260.6000 136.1000 261.0000 136.2000 ;
	    RECT 258.2000 135.8000 261.0000 136.1000 ;
	    RECT 266.2000 135.8000 266.6000 136.2000 ;
	    RECT 7.0000 135.1000 7.4000 135.2000 ;
	    RECT 10.2000 135.1000 10.6000 135.2000 ;
	    RECT 11.8000 135.1000 12.2000 135.2000 ;
	    RECT 7.0000 134.8000 12.2000 135.1000 ;
	    RECT 16.6000 135.1000 17.0000 135.2000 ;
	    RECT 20.6000 135.1000 21.0000 135.2000 ;
	    RECT 16.6000 134.8000 21.0000 135.1000 ;
	    RECT 23.8000 135.1000 24.2000 135.2000 ;
	    RECT 27.0000 135.1000 27.4000 135.2000 ;
	    RECT 29.4000 135.1000 29.8000 135.2000 ;
	    RECT 36.6000 135.1000 37.0000 135.2000 ;
	    RECT 42.2000 135.1000 42.5000 135.8000 ;
	    RECT 266.2000 135.2000 266.5000 135.8000 ;
	    RECT 23.8000 134.8000 29.8000 135.1000 ;
	    RECT 35.8000 134.8000 42.5000 135.1000 ;
	    RECT 51.8000 134.8000 52.2000 135.2000 ;
	    RECT 57.4000 135.1000 57.8000 135.2000 ;
	    RECT 66.2000 135.1000 66.6000 135.2000 ;
	    RECT 57.4000 134.8000 66.6000 135.1000 ;
	    RECT 67.8000 135.1000 68.2000 135.2000 ;
	    RECT 92.6000 135.1000 93.0000 135.2000 ;
	    RECT 111.8000 135.1000 112.2000 135.2000 ;
	    RECT 67.8000 134.8000 79.3000 135.1000 ;
	    RECT 92.6000 134.8000 112.2000 135.1000 ;
	    RECT 117.4000 135.1000 117.8000 135.2000 ;
	    RECT 123.8000 135.1000 124.2000 135.2000 ;
	    RECT 117.4000 134.8000 124.2000 135.1000 ;
	    RECT 135.0000 135.1000 135.4000 135.2000 ;
	    RECT 142.2000 135.1000 142.6000 135.2000 ;
	    RECT 135.0000 134.8000 142.6000 135.1000 ;
	    RECT 158.2000 135.1000 158.6000 135.2000 ;
	    RECT 175.0000 135.1000 175.4000 135.2000 ;
	    RECT 158.2000 134.8000 175.4000 135.1000 ;
	    RECT 183.0000 135.1000 183.4000 135.2000 ;
	    RECT 185.4000 135.1000 185.8000 135.2000 ;
	    RECT 187.8000 135.1000 188.2000 135.2000 ;
	    RECT 183.0000 134.8000 188.2000 135.1000 ;
	    RECT 190.2000 135.1000 190.6000 135.2000 ;
	    RECT 196.6000 135.1000 197.0000 135.2000 ;
	    RECT 198.2000 135.1000 198.6000 135.2000 ;
	    RECT 190.2000 134.8000 198.6000 135.1000 ;
	    RECT 206.2000 135.1000 206.6000 135.2000 ;
	    RECT 217.4000 135.1000 217.8000 135.2000 ;
	    RECT 219.8000 135.1000 220.2000 135.2000 ;
	    RECT 224.6000 135.1000 225.0000 135.2000 ;
	    RECT 206.2000 134.8000 225.0000 135.1000 ;
	    RECT 225.4000 135.1000 225.8000 135.2000 ;
	    RECT 235.8000 135.1000 236.2000 135.2000 ;
	    RECT 242.2000 135.1000 242.6000 135.2000 ;
	    RECT 225.4000 134.8000 242.6000 135.1000 ;
	    RECT 246.2000 135.1000 246.6000 135.2000 ;
	    RECT 248.6000 135.1000 249.0000 135.2000 ;
	    RECT 246.2000 134.8000 249.0000 135.1000 ;
	    RECT 250.2000 135.1000 250.6000 135.2000 ;
	    RECT 251.8000 135.1000 252.2000 135.2000 ;
	    RECT 250.2000 134.8000 252.2000 135.1000 ;
	    RECT 253.4000 134.8000 253.8000 135.2000 ;
	    RECT 259.8000 134.8000 260.2000 135.2000 ;
	    RECT 266.2000 134.8000 266.6000 135.2000 ;
	    RECT 51.8000 134.1000 52.1000 134.8000 ;
	    RECT 48.6000 133.8000 52.1000 134.1000 ;
	    RECT 79.0000 134.2000 79.3000 134.8000 ;
	    RECT 79.0000 133.8000 79.4000 134.2000 ;
	    RECT 175.8000 134.1000 176.2000 134.2000 ;
	    RECT 176.6000 134.1000 177.0000 134.2000 ;
	    RECT 175.8000 133.8000 177.0000 134.1000 ;
	    RECT 180.6000 134.1000 181.0000 134.2000 ;
	    RECT 183.0000 134.1000 183.4000 134.2000 ;
	    RECT 192.6000 134.1000 193.0000 134.2000 ;
	    RECT 180.6000 133.8000 193.0000 134.1000 ;
	    RECT 194.2000 134.1000 194.6000 134.2000 ;
	    RECT 197.4000 134.1000 197.8000 134.2000 ;
	    RECT 194.2000 133.8000 197.8000 134.1000 ;
	    RECT 215.8000 134.1000 216.2000 134.2000 ;
	    RECT 226.2000 134.1000 226.6000 134.2000 ;
	    RECT 215.8000 133.8000 226.6000 134.1000 ;
	    RECT 230.2000 134.1000 230.6000 134.2000 ;
	    RECT 232.6000 134.1000 233.0000 134.2000 ;
	    RECT 230.2000 133.8000 233.0000 134.1000 ;
	    RECT 253.4000 134.1000 253.7000 134.8000 ;
	    RECT 256.6000 134.1000 257.0000 134.2000 ;
	    RECT 253.4000 133.8000 257.0000 134.1000 ;
	    RECT 259.8000 134.1000 260.1000 134.8000 ;
	    RECT 262.2000 134.1000 262.6000 134.2000 ;
	    RECT 259.8000 133.8000 262.6000 134.1000 ;
	    RECT 266.2000 134.1000 266.6000 134.2000 ;
	    RECT 267.8000 134.1000 268.2000 134.2000 ;
	    RECT 266.2000 133.8000 268.2000 134.1000 ;
	    RECT 48.6000 133.2000 48.9000 133.8000 ;
	    RECT 2.2000 133.1000 2.6000 133.2000 ;
	    RECT 7.0000 133.1000 7.4000 133.2000 ;
	    RECT 2.2000 132.8000 7.4000 133.1000 ;
	    RECT 10.2000 133.1000 10.6000 133.2000 ;
	    RECT 31.8000 133.1000 32.2000 133.2000 ;
	    RECT 10.2000 132.8000 32.2000 133.1000 ;
	    RECT 39.0000 133.1000 39.4000 133.2000 ;
	    RECT 48.6000 133.1000 49.0000 133.2000 ;
	    RECT 39.0000 132.8000 49.0000 133.1000 ;
	    RECT 51.0000 133.1000 51.4000 133.2000 ;
	    RECT 52.6000 133.1000 53.0000 133.2000 ;
	    RECT 51.0000 132.8000 53.0000 133.1000 ;
	    RECT 95.0000 133.1000 95.4000 133.2000 ;
	    RECT 98.2000 133.1000 98.6000 133.2000 ;
	    RECT 95.0000 132.8000 98.6000 133.1000 ;
	    RECT 103.8000 133.1000 104.2000 133.2000 ;
	    RECT 107.0000 133.1000 107.4000 133.2000 ;
	    RECT 103.8000 132.8000 107.4000 133.1000 ;
	    RECT 111.8000 133.1000 112.2000 133.2000 ;
	    RECT 117.4000 133.1000 117.8000 133.2000 ;
	    RECT 111.8000 132.8000 117.8000 133.1000 ;
	    RECT 118.2000 133.1000 118.6000 133.2000 ;
	    RECT 119.8000 133.1000 120.2000 133.2000 ;
	    RECT 118.2000 132.8000 120.2000 133.1000 ;
	    RECT 166.2000 133.1000 166.6000 133.2000 ;
	    RECT 176.6000 133.1000 177.0000 133.2000 ;
	    RECT 201.4000 133.1000 201.8000 133.2000 ;
	    RECT 207.0000 133.1000 207.4000 133.2000 ;
	    RECT 207.8000 133.1000 208.2000 133.2000 ;
	    RECT 166.2000 132.8000 208.2000 133.1000 ;
	    RECT 208.6000 133.1000 209.0000 133.2000 ;
	    RECT 211.8000 133.1000 212.2000 133.2000 ;
	    RECT 208.6000 132.8000 212.2000 133.1000 ;
	    RECT 213.4000 132.8000 213.8000 133.2000 ;
	    RECT 215.0000 133.1000 215.4000 133.2000 ;
	    RECT 219.0000 133.1000 219.4000 133.2000 ;
	    RECT 215.0000 132.8000 219.4000 133.1000 ;
	    RECT 222.2000 133.1000 222.6000 133.2000 ;
	    RECT 225.4000 133.1000 225.8000 133.2000 ;
	    RECT 222.2000 132.8000 225.8000 133.1000 ;
	    RECT 228.6000 133.1000 229.0000 133.2000 ;
	    RECT 231.0000 133.1000 231.4000 133.2000 ;
	    RECT 228.6000 132.8000 231.4000 133.1000 ;
	    RECT 237.4000 133.1000 237.8000 133.2000 ;
	    RECT 239.0000 133.1000 239.4000 133.2000 ;
	    RECT 254.2000 133.1000 254.6000 133.2000 ;
	    RECT 237.4000 132.8000 239.4000 133.1000 ;
	    RECT 252.6000 132.8000 254.6000 133.1000 ;
	    RECT 259.0000 133.1000 259.4000 133.2000 ;
	    RECT 260.6000 133.1000 261.0000 133.2000 ;
	    RECT 259.0000 132.8000 261.0000 133.1000 ;
	    RECT 39.0000 132.1000 39.4000 132.2000 ;
	    RECT 58.2000 132.1000 58.6000 132.2000 ;
	    RECT 39.0000 131.8000 58.6000 132.1000 ;
	    RECT 100.6000 132.1000 101.0000 132.2000 ;
	    RECT 103.8000 132.1000 104.2000 132.2000 ;
	    RECT 114.2000 132.1000 114.6000 132.2000 ;
	    RECT 118.2000 132.1000 118.6000 132.2000 ;
	    RECT 100.6000 131.8000 118.6000 132.1000 ;
	    RECT 127.8000 132.1000 128.2000 132.2000 ;
	    RECT 134.2000 132.1000 134.6000 132.2000 ;
	    RECT 127.8000 131.8000 134.6000 132.1000 ;
	    RECT 156.6000 132.1000 157.0000 132.2000 ;
	    RECT 159.0000 132.1000 159.4000 132.2000 ;
	    RECT 156.6000 131.8000 159.4000 132.1000 ;
	    RECT 205.4000 132.1000 205.8000 132.2000 ;
	    RECT 213.4000 132.1000 213.7000 132.8000 ;
	    RECT 252.6000 132.2000 252.9000 132.8000 ;
	    RECT 205.4000 131.8000 213.7000 132.1000 ;
	    RECT 225.4000 132.1000 225.8000 132.2000 ;
	    RECT 238.2000 132.1000 238.6000 132.2000 ;
	    RECT 225.4000 131.8000 238.6000 132.1000 ;
	    RECT 245.4000 132.1000 245.8000 132.2000 ;
	    RECT 250.2000 132.1000 250.6000 132.2000 ;
	    RECT 245.4000 131.8000 250.6000 132.1000 ;
	    RECT 252.6000 131.8000 253.0000 132.2000 ;
	    RECT 39.0000 131.2000 39.3000 131.8000 ;
	    RECT 19.8000 131.1000 20.2000 131.2000 ;
	    RECT 26.2000 131.1000 26.6000 131.2000 ;
	    RECT 19.8000 130.8000 26.6000 131.1000 ;
	    RECT 39.0000 130.8000 39.4000 131.2000 ;
	    RECT 88.6000 131.1000 89.0000 131.2000 ;
	    RECT 105.4000 131.1000 105.8000 131.2000 ;
	    RECT 88.6000 130.8000 105.8000 131.1000 ;
	    RECT 191.0000 131.1000 191.4000 131.2000 ;
	    RECT 191.8000 131.1000 192.2000 131.2000 ;
	    RECT 194.2000 131.1000 194.6000 131.2000 ;
	    RECT 191.0000 130.8000 194.6000 131.1000 ;
	    RECT 218.2000 131.1000 218.6000 131.2000 ;
	    RECT 230.2000 131.1000 230.6000 131.2000 ;
	    RECT 218.2000 130.8000 230.6000 131.1000 ;
	    RECT 231.8000 130.8000 232.2000 131.2000 ;
	    RECT 239.8000 131.1000 240.2000 131.2000 ;
	    RECT 255.0000 131.1000 255.4000 131.2000 ;
	    RECT 257.4000 131.1000 257.8000 131.2000 ;
	    RECT 239.8000 130.8000 257.8000 131.1000 ;
	    RECT 231.8000 130.2000 232.1000 130.8000 ;
	    RECT 22.2000 130.1000 22.6000 130.2000 ;
	    RECT 24.6000 130.1000 25.0000 130.2000 ;
	    RECT 22.2000 129.8000 25.0000 130.1000 ;
	    RECT 231.8000 129.8000 232.2000 130.2000 ;
	    RECT 243.0000 130.1000 243.4000 130.2000 ;
	    RECT 232.6000 129.8000 243.4000 130.1000 ;
	    RECT 257.4000 130.1000 257.8000 130.2000 ;
	    RECT 262.2000 130.1000 262.6000 130.2000 ;
	    RECT 257.4000 129.8000 262.6000 130.1000 ;
	    RECT 232.6000 129.2000 232.9000 129.8000 ;
	    RECT 1.4000 129.1000 1.8000 129.2000 ;
	    RECT 4.6000 129.1000 5.0000 129.2000 ;
	    RECT 7.0000 129.1000 7.4000 129.2000 ;
	    RECT 1.4000 128.8000 7.4000 129.1000 ;
	    RECT 23.8000 128.8000 24.2000 129.2000 ;
	    RECT 38.2000 128.8000 38.6000 129.2000 ;
	    RECT 42.2000 129.1000 42.6000 129.2000 ;
	    RECT 49.4000 129.1000 49.8000 129.2000 ;
	    RECT 62.2000 129.1000 62.6000 129.2000 ;
	    RECT 72.6000 129.1000 73.0000 129.2000 ;
	    RECT 42.2000 128.8000 73.0000 129.1000 ;
	    RECT 106.2000 129.1000 106.6000 129.2000 ;
	    RECT 111.8000 129.1000 112.2000 129.2000 ;
	    RECT 106.2000 128.8000 112.2000 129.1000 ;
	    RECT 113.4000 128.8000 113.8000 129.2000 ;
	    RECT 124.6000 129.1000 125.0000 129.2000 ;
	    RECT 128.6000 129.1000 129.0000 129.2000 ;
	    RECT 124.6000 128.8000 129.0000 129.1000 ;
	    RECT 193.4000 129.1000 193.8000 129.2000 ;
	    RECT 232.6000 129.1000 233.0000 129.2000 ;
	    RECT 193.4000 128.8000 233.0000 129.1000 ;
	    RECT 235.0000 129.1000 235.4000 129.2000 ;
	    RECT 243.0000 129.1000 243.4000 129.2000 ;
	    RECT 235.0000 128.8000 243.4000 129.1000 ;
	    RECT 253.4000 128.8000 253.8000 129.2000 ;
	    RECT 255.8000 128.8000 256.2000 129.2000 ;
	    RECT 259.8000 128.8000 260.2000 129.2000 ;
	    RECT 23.8000 128.1000 24.1000 128.8000 ;
	    RECT 26.2000 128.1000 26.6000 128.2000 ;
	    RECT 23.8000 127.8000 26.6000 128.1000 ;
	    RECT 28.6000 128.1000 29.0000 128.2000 ;
	    RECT 30.2000 128.1000 30.6000 128.2000 ;
	    RECT 28.6000 127.8000 30.6000 128.1000 ;
	    RECT 32.6000 128.1000 33.0000 128.2000 ;
	    RECT 34.2000 128.1000 34.6000 128.2000 ;
	    RECT 32.6000 127.8000 34.6000 128.1000 ;
	    RECT 35.0000 128.1000 35.4000 128.2000 ;
	    RECT 38.2000 128.1000 38.5000 128.8000 ;
	    RECT 113.4000 128.2000 113.7000 128.8000 ;
	    RECT 35.0000 127.8000 38.5000 128.1000 ;
	    RECT 43.8000 128.1000 44.2000 128.2000 ;
	    RECT 52.6000 128.1000 53.0000 128.2000 ;
	    RECT 53.4000 128.1000 53.8000 128.2000 ;
	    RECT 43.8000 127.8000 53.8000 128.1000 ;
	    RECT 63.0000 128.1000 63.4000 128.2000 ;
	    RECT 75.0000 128.1000 75.4000 128.2000 ;
	    RECT 63.0000 127.8000 75.4000 128.1000 ;
	    RECT 79.0000 127.8000 79.4000 128.2000 ;
	    RECT 99.8000 128.1000 100.2000 128.2000 ;
	    RECT 105.4000 128.1000 105.8000 128.2000 ;
	    RECT 99.8000 127.8000 105.8000 128.1000 ;
	    RECT 113.4000 127.8000 113.8000 128.2000 ;
	    RECT 114.2000 128.1000 114.6000 128.2000 ;
	    RECT 115.8000 128.1000 116.2000 128.2000 ;
	    RECT 114.2000 127.8000 116.2000 128.1000 ;
	    RECT 126.2000 127.8000 126.6000 128.2000 ;
	    RECT 130.2000 127.8000 130.6000 128.2000 ;
	    RECT 147.8000 128.1000 148.2000 128.2000 ;
	    RECT 150.2000 128.1000 150.6000 128.2000 ;
	    RECT 147.8000 127.8000 150.6000 128.1000 ;
	    RECT 152.6000 128.1000 153.0000 128.2000 ;
	    RECT 153.4000 128.1000 153.8000 128.2000 ;
	    RECT 152.6000 127.8000 153.8000 128.1000 ;
	    RECT 158.2000 128.1000 158.6000 128.2000 ;
	    RECT 159.0000 128.1000 159.4000 128.2000 ;
	    RECT 158.2000 127.8000 159.4000 128.1000 ;
	    RECT 174.2000 128.1000 174.6000 128.2000 ;
	    RECT 180.6000 128.1000 181.0000 128.2000 ;
	    RECT 191.8000 128.1000 192.2000 128.2000 ;
	    RECT 195.0000 128.1000 195.4000 128.2000 ;
	    RECT 207.8000 128.1000 208.2000 128.2000 ;
	    RECT 214.2000 128.1000 214.6000 128.2000 ;
	    RECT 174.2000 127.8000 214.6000 128.1000 ;
	    RECT 216.6000 128.1000 217.0000 128.2000 ;
	    RECT 217.4000 128.1000 217.8000 128.2000 ;
	    RECT 216.6000 127.8000 217.8000 128.1000 ;
	    RECT 223.8000 127.8000 224.2000 128.2000 ;
	    RECT 235.8000 128.1000 236.2000 128.2000 ;
	    RECT 247.0000 128.1000 247.4000 128.2000 ;
	    RECT 235.8000 127.8000 247.4000 128.1000 ;
	    RECT 253.4000 128.1000 253.7000 128.8000 ;
	    RECT 255.8000 128.1000 256.1000 128.8000 ;
	    RECT 253.4000 127.8000 256.1000 128.1000 ;
	    RECT 259.8000 128.1000 260.1000 128.8000 ;
	    RECT 263.0000 128.1000 263.4000 128.2000 ;
	    RECT 259.8000 127.8000 263.4000 128.1000 ;
	    RECT 30.2000 126.8000 30.6000 127.2000 ;
	    RECT 31.0000 127.1000 31.4000 127.2000 ;
	    RECT 35.8000 127.1000 36.2000 127.2000 ;
	    RECT 37.4000 127.1000 37.8000 127.2000 ;
	    RECT 42.2000 127.1000 42.6000 127.2000 ;
	    RECT 31.0000 126.8000 42.6000 127.1000 ;
	    RECT 64.6000 126.8000 65.0000 127.2000 ;
	    RECT 66.2000 126.8000 66.6000 127.2000 ;
	    RECT 75.0000 127.1000 75.4000 127.2000 ;
	    RECT 79.0000 127.1000 79.3000 127.8000 ;
	    RECT 93.4000 127.1000 93.8000 127.2000 ;
	    RECT 100.6000 127.1000 101.0000 127.2000 ;
	    RECT 75.0000 126.8000 79.3000 127.1000 ;
	    RECT 83.8000 126.8000 93.8000 127.1000 ;
	    RECT 99.0000 126.8000 101.0000 127.1000 ;
	    RECT 113.4000 127.1000 113.8000 127.2000 ;
	    RECT 119.8000 127.1000 120.2000 127.2000 ;
	    RECT 126.2000 127.1000 126.5000 127.8000 ;
	    RECT 113.4000 126.8000 126.5000 127.1000 ;
	    RECT 127.0000 127.1000 127.4000 127.2000 ;
	    RECT 130.2000 127.1000 130.5000 127.8000 ;
	    RECT 223.8000 127.2000 224.1000 127.8000 ;
	    RECT 127.0000 126.8000 130.5000 127.1000 ;
	    RECT 133.4000 127.1000 133.8000 127.2000 ;
	    RECT 140.6000 127.1000 141.0000 127.2000 ;
	    RECT 133.4000 126.8000 141.0000 127.1000 ;
	    RECT 146.2000 127.1000 146.6000 127.2000 ;
	    RECT 147.0000 127.1000 147.4000 127.2000 ;
	    RECT 146.2000 126.8000 147.4000 127.1000 ;
	    RECT 177.4000 127.1000 177.8000 127.2000 ;
	    RECT 183.0000 127.1000 183.4000 127.2000 ;
	    RECT 189.4000 127.1000 189.8000 127.2000 ;
	    RECT 208.6000 127.1000 209.0000 127.2000 ;
	    RECT 211.0000 127.1000 211.4000 127.2000 ;
	    RECT 177.4000 126.8000 211.4000 127.1000 ;
	    RECT 223.8000 126.8000 224.2000 127.2000 ;
	    RECT 227.0000 127.1000 227.4000 127.2000 ;
	    RECT 228.6000 127.1000 229.0000 127.2000 ;
	    RECT 227.0000 126.8000 229.0000 127.1000 ;
	    RECT 230.2000 127.1000 230.6000 127.2000 ;
	    RECT 233.4000 127.1000 233.8000 127.2000 ;
	    RECT 230.2000 126.8000 233.8000 127.1000 ;
	    RECT 262.2000 127.1000 262.6000 127.2000 ;
	    RECT 264.6000 127.1000 265.0000 127.2000 ;
	    RECT 262.2000 126.8000 265.0000 127.1000 ;
	    RECT 7.0000 126.1000 7.4000 126.2000 ;
	    RECT 8.6000 126.1000 9.0000 126.2000 ;
	    RECT 7.0000 125.8000 9.0000 126.1000 ;
	    RECT 16.6000 125.8000 17.0000 126.2000 ;
	    RECT 18.2000 126.1000 18.6000 126.2000 ;
	    RECT 19.0000 126.1000 19.4000 126.2000 ;
	    RECT 18.2000 125.8000 19.4000 126.1000 ;
	    RECT 30.2000 126.1000 30.5000 126.8000 ;
	    RECT 34.2000 126.1000 34.6000 126.2000 ;
	    RECT 54.2000 126.1000 54.6000 126.2000 ;
	    RECT 30.2000 125.8000 54.6000 126.1000 ;
	    RECT 55.8000 126.1000 56.2000 126.2000 ;
	    RECT 57.4000 126.1000 57.8000 126.2000 ;
	    RECT 55.8000 125.8000 57.8000 126.1000 ;
	    RECT 64.6000 126.1000 64.9000 126.8000 ;
	    RECT 66.2000 126.1000 66.5000 126.8000 ;
	    RECT 83.8000 126.2000 84.1000 126.8000 ;
	    RECT 99.0000 126.6000 99.4000 126.8000 ;
	    RECT 64.6000 125.8000 66.5000 126.1000 ;
	    RECT 76.6000 126.1000 77.0000 126.2000 ;
	    RECT 79.8000 126.1000 80.2000 126.2000 ;
	    RECT 76.6000 125.8000 80.2000 126.1000 ;
	    RECT 83.8000 125.8000 84.2000 126.2000 ;
	    RECT 111.0000 126.1000 111.4000 126.2000 ;
	    RECT 119.0000 126.1000 119.4000 126.2000 ;
	    RECT 125.4000 126.1000 125.8000 126.2000 ;
	    RECT 111.0000 125.8000 125.8000 126.1000 ;
	    RECT 138.2000 126.1000 138.6000 126.2000 ;
	    RECT 145.4000 126.1000 145.8000 126.2000 ;
	    RECT 147.0000 126.1000 147.4000 126.2000 ;
	    RECT 152.6000 126.1000 153.0000 126.2000 ;
	    RECT 138.2000 125.8000 153.0000 126.1000 ;
	    RECT 174.2000 126.1000 174.6000 126.2000 ;
	    RECT 179.0000 126.1000 179.4000 126.2000 ;
	    RECT 185.4000 126.1000 185.8000 126.2000 ;
	    RECT 174.2000 125.8000 185.8000 126.1000 ;
	    RECT 193.4000 126.1000 193.8000 126.2000 ;
	    RECT 197.4000 126.1000 197.8000 126.2000 ;
	    RECT 205.4000 126.1000 205.8000 126.2000 ;
	    RECT 193.4000 125.8000 197.8000 126.1000 ;
	    RECT 202.2000 125.8000 205.8000 126.1000 ;
	    RECT 208.6000 125.8000 209.0000 126.2000 ;
	    RECT 212.6000 126.1000 213.0000 126.2000 ;
	    RECT 215.8000 126.1000 216.2000 126.2000 ;
	    RECT 223.0000 126.1000 223.4000 126.2000 ;
	    RECT 225.4000 126.1000 225.8000 126.2000 ;
	    RECT 212.6000 125.8000 225.8000 126.1000 ;
	    RECT 227.8000 126.1000 228.2000 126.2000 ;
	    RECT 236.6000 126.1000 237.0000 126.2000 ;
	    RECT 227.8000 125.8000 237.0000 126.1000 ;
	    RECT 239.8000 126.1000 240.2000 126.2000 ;
	    RECT 240.6000 126.1000 241.0000 126.2000 ;
	    RECT 245.4000 126.1000 245.8000 126.2000 ;
	    RECT 239.8000 125.8000 245.8000 126.1000 ;
	    RECT 249.4000 126.1000 249.8000 126.2000 ;
	    RECT 266.2000 126.1000 266.6000 126.2000 ;
	    RECT 249.4000 125.8000 266.6000 126.1000 ;
	    RECT 16.6000 125.1000 16.9000 125.8000 ;
	    RECT 202.2000 125.2000 202.5000 125.8000 ;
	    RECT 21.4000 125.1000 21.8000 125.2000 ;
	    RECT 16.6000 124.8000 21.8000 125.1000 ;
	    RECT 27.0000 125.1000 27.4000 125.2000 ;
	    RECT 39.0000 125.1000 39.4000 125.2000 ;
	    RECT 47.0000 125.1000 47.4000 125.2000 ;
	    RECT 27.0000 124.8000 39.4000 125.1000 ;
	    RECT 41.4000 124.8000 47.4000 125.1000 ;
	    RECT 81.4000 124.8000 81.8000 125.2000 ;
	    RECT 97.4000 125.1000 97.8000 125.2000 ;
	    RECT 101.4000 125.1000 101.8000 125.2000 ;
	    RECT 97.4000 124.8000 101.8000 125.1000 ;
	    RECT 113.4000 125.1000 113.8000 125.2000 ;
	    RECT 114.2000 125.1000 114.6000 125.2000 ;
	    RECT 113.4000 124.8000 114.6000 125.1000 ;
	    RECT 117.4000 125.1000 117.8000 125.2000 ;
	    RECT 128.6000 125.1000 129.0000 125.2000 ;
	    RECT 139.0000 125.1000 139.4000 125.2000 ;
	    RECT 117.4000 124.8000 139.4000 125.1000 ;
	    RECT 151.0000 125.1000 151.4000 125.2000 ;
	    RECT 158.2000 125.1000 158.6000 125.2000 ;
	    RECT 151.0000 124.8000 158.6000 125.1000 ;
	    RECT 175.0000 125.1000 175.4000 125.2000 ;
	    RECT 185.4000 125.1000 185.8000 125.2000 ;
	    RECT 175.0000 124.8000 185.8000 125.1000 ;
	    RECT 202.2000 124.8000 202.6000 125.2000 ;
	    RECT 208.6000 125.1000 208.9000 125.8000 ;
	    RECT 214.2000 125.1000 214.6000 125.2000 ;
	    RECT 224.6000 125.1000 225.0000 125.2000 ;
	    RECT 226.2000 125.1000 226.6000 125.2000 ;
	    RECT 208.6000 124.8000 226.6000 125.1000 ;
	    RECT 238.2000 125.1000 238.6000 125.2000 ;
	    RECT 258.2000 125.1000 258.6000 125.2000 ;
	    RECT 238.2000 124.8000 243.3000 125.1000 ;
	    RECT 41.4000 124.2000 41.7000 124.8000 ;
	    RECT 23.8000 124.1000 24.2000 124.2000 ;
	    RECT 27.0000 124.1000 27.4000 124.2000 ;
	    RECT 23.8000 123.8000 27.4000 124.1000 ;
	    RECT 41.4000 123.8000 41.8000 124.2000 ;
	    RECT 48.6000 124.1000 49.0000 124.2000 ;
	    RECT 69.4000 124.1000 69.8000 124.2000 ;
	    RECT 81.4000 124.1000 81.7000 124.8000 ;
	    RECT 243.0000 124.2000 243.3000 124.8000 ;
	    RECT 243.8000 124.8000 258.6000 125.1000 ;
	    RECT 243.8000 124.2000 244.1000 124.8000 ;
	    RECT 48.6000 123.8000 81.7000 124.1000 ;
	    RECT 115.8000 124.1000 116.2000 124.2000 ;
	    RECT 121.4000 124.1000 121.8000 124.2000 ;
	    RECT 126.2000 124.1000 126.6000 124.2000 ;
	    RECT 140.6000 124.1000 141.0000 124.2000 ;
	    RECT 142.2000 124.1000 142.6000 124.2000 ;
	    RECT 156.6000 124.1000 157.0000 124.2000 ;
	    RECT 115.8000 123.8000 116.9000 124.1000 ;
	    RECT 121.4000 123.8000 157.0000 124.1000 ;
	    RECT 189.4000 124.1000 189.8000 124.2000 ;
	    RECT 192.6000 124.1000 193.0000 124.2000 ;
	    RECT 189.4000 123.8000 193.0000 124.1000 ;
	    RECT 207.0000 124.1000 207.4000 124.2000 ;
	    RECT 216.6000 124.1000 217.0000 124.2000 ;
	    RECT 207.0000 123.8000 217.0000 124.1000 ;
	    RECT 219.8000 124.1000 220.2000 124.2000 ;
	    RECT 221.4000 124.1000 221.8000 124.2000 ;
	    RECT 219.8000 123.8000 221.8000 124.1000 ;
	    RECT 222.2000 124.1000 222.6000 124.2000 ;
	    RECT 223.0000 124.1000 223.4000 124.2000 ;
	    RECT 222.2000 123.8000 223.4000 124.1000 ;
	    RECT 235.0000 124.1000 235.4000 124.2000 ;
	    RECT 235.8000 124.1000 236.2000 124.2000 ;
	    RECT 235.0000 123.8000 236.2000 124.1000 ;
	    RECT 240.6000 123.8000 241.0000 124.2000 ;
	    RECT 243.0000 123.8000 243.4000 124.2000 ;
	    RECT 243.8000 123.8000 244.2000 124.2000 ;
	    RECT 116.6000 123.2000 116.9000 123.8000 ;
	    RECT 18.2000 123.1000 18.6000 123.2000 ;
	    RECT 31.8000 123.1000 32.2000 123.2000 ;
	    RECT 18.2000 122.8000 32.2000 123.1000 ;
	    RECT 35.0000 123.1000 35.4000 123.2000 ;
	    RECT 65.4000 123.1000 65.8000 123.2000 ;
	    RECT 35.0000 122.8000 65.8000 123.1000 ;
	    RECT 96.6000 123.1000 97.0000 123.2000 ;
	    RECT 97.4000 123.1000 97.8000 123.2000 ;
	    RECT 113.4000 123.1000 113.8000 123.2000 ;
	    RECT 96.6000 122.8000 113.8000 123.1000 ;
	    RECT 116.6000 122.8000 117.0000 123.2000 ;
	    RECT 128.6000 123.1000 129.0000 123.2000 ;
	    RECT 139.8000 123.1000 140.2000 123.2000 ;
	    RECT 144.6000 123.1000 145.0000 123.2000 ;
	    RECT 148.6000 123.1000 149.0000 123.2000 ;
	    RECT 128.6000 122.8000 149.0000 123.1000 ;
	    RECT 178.2000 123.1000 178.6000 123.2000 ;
	    RECT 217.4000 123.1000 217.8000 123.2000 ;
	    RECT 238.2000 123.1000 238.6000 123.2000 ;
	    RECT 239.0000 123.1000 239.4000 123.2000 ;
	    RECT 178.2000 122.8000 239.4000 123.1000 ;
	    RECT 240.6000 123.1000 240.9000 123.8000 ;
	    RECT 251.0000 123.1000 251.4000 123.2000 ;
	    RECT 240.6000 122.8000 251.4000 123.1000 ;
	    RECT 43.0000 122.1000 43.4000 122.2000 ;
	    RECT 46.2000 122.1000 46.6000 122.2000 ;
	    RECT 60.6000 122.1000 61.0000 122.2000 ;
	    RECT 43.0000 121.8000 61.0000 122.1000 ;
	    RECT 82.2000 122.1000 82.6000 122.2000 ;
	    RECT 84.6000 122.1000 85.0000 122.2000 ;
	    RECT 91.8000 122.1000 92.2000 122.2000 ;
	    RECT 82.2000 121.8000 92.2000 122.1000 ;
	    RECT 213.4000 122.1000 213.8000 122.2000 ;
	    RECT 232.6000 122.1000 233.0000 122.2000 ;
	    RECT 213.4000 121.8000 233.0000 122.1000 ;
	    RECT 105.4000 121.1000 105.8000 121.2000 ;
	    RECT 121.4000 121.1000 121.8000 121.2000 ;
	    RECT 105.4000 120.8000 121.8000 121.1000 ;
	    RECT 210.2000 121.1000 210.6000 121.2000 ;
	    RECT 223.8000 121.1000 224.2000 121.2000 ;
	    RECT 210.2000 120.8000 224.2000 121.1000 ;
	    RECT 234.2000 121.1000 234.6000 121.2000 ;
	    RECT 259.0000 121.1000 259.4000 121.2000 ;
	    RECT 234.2000 120.8000 259.4000 121.1000 ;
	    RECT 95.0000 120.1000 95.4000 120.2000 ;
	    RECT 121.4000 120.1000 121.8000 120.2000 ;
	    RECT 95.0000 119.8000 121.8000 120.1000 ;
	    RECT 132.6000 120.1000 133.0000 120.2000 ;
	    RECT 141.4000 120.1000 141.8000 120.2000 ;
	    RECT 144.6000 120.1000 145.0000 120.2000 ;
	    RECT 132.6000 119.8000 145.0000 120.1000 ;
	    RECT 230.2000 120.1000 230.6000 120.2000 ;
	    RECT 243.0000 120.1000 243.4000 120.2000 ;
	    RECT 230.2000 119.8000 243.4000 120.1000 ;
	    RECT 159.8000 119.1000 160.2000 119.2000 ;
	    RECT 168.6000 119.1000 169.0000 119.2000 ;
	    RECT 159.8000 118.8000 169.0000 119.1000 ;
	    RECT 243.0000 119.1000 243.4000 119.2000 ;
	    RECT 255.0000 119.1000 255.4000 119.2000 ;
	    RECT 243.0000 118.8000 255.4000 119.1000 ;
	    RECT 30.2000 117.8000 30.6000 118.2000 ;
	    RECT 101.4000 118.1000 101.8000 118.2000 ;
	    RECT 135.8000 118.1000 136.2000 118.2000 ;
	    RECT 152.6000 118.1000 153.0000 118.2000 ;
	    RECT 155.0000 118.1000 155.4000 118.2000 ;
	    RECT 101.4000 117.8000 155.4000 118.1000 ;
	    RECT 173.4000 118.1000 173.8000 118.2000 ;
	    RECT 183.8000 118.1000 184.2000 118.2000 ;
	    RECT 229.4000 118.1000 229.8000 118.2000 ;
	    RECT 252.6000 118.1000 253.0000 118.2000 ;
	    RECT 173.4000 117.8000 253.0000 118.1000 ;
	    RECT 30.2000 117.1000 30.5000 117.8000 ;
	    RECT 35.0000 117.1000 35.4000 117.2000 ;
	    RECT 30.2000 116.8000 35.4000 117.1000 ;
	    RECT 42.2000 117.1000 42.6000 117.2000 ;
	    RECT 50.2000 117.1000 50.6000 117.2000 ;
	    RECT 55.8000 117.1000 56.2000 117.2000 ;
	    RECT 70.2000 117.1000 70.6000 117.2000 ;
	    RECT 42.2000 116.8000 70.6000 117.1000 ;
	    RECT 73.4000 117.1000 73.8000 117.2000 ;
	    RECT 75.0000 117.1000 75.4000 117.2000 ;
	    RECT 73.4000 116.8000 75.4000 117.1000 ;
	    RECT 106.2000 117.1000 106.6000 117.2000 ;
	    RECT 128.6000 117.1000 129.0000 117.2000 ;
	    RECT 106.2000 116.8000 129.0000 117.1000 ;
	    RECT 130.2000 117.1000 130.6000 117.2000 ;
	    RECT 131.0000 117.1000 131.4000 117.2000 ;
	    RECT 130.2000 116.8000 131.4000 117.1000 ;
	    RECT 134.2000 116.8000 134.6000 117.2000 ;
	    RECT 151.8000 116.8000 152.2000 117.2000 ;
	    RECT 181.4000 117.1000 181.8000 117.2000 ;
	    RECT 186.2000 117.1000 186.6000 117.2000 ;
	    RECT 181.4000 116.8000 186.6000 117.1000 ;
	    RECT 191.0000 117.1000 191.4000 117.2000 ;
	    RECT 194.2000 117.1000 194.6000 117.2000 ;
	    RECT 222.2000 117.1000 222.6000 117.2000 ;
	    RECT 235.0000 117.1000 235.4000 117.2000 ;
	    RECT 239.0000 117.1000 239.4000 117.2000 ;
	    RECT 191.0000 116.8000 239.4000 117.1000 ;
	    RECT 240.6000 117.1000 241.0000 117.2000 ;
	    RECT 255.8000 117.1000 256.2000 117.2000 ;
	    RECT 240.6000 116.8000 256.2000 117.1000 ;
	    RECT 29.4000 116.1000 29.8000 116.2000 ;
	    RECT 33.4000 116.1000 33.8000 116.2000 ;
	    RECT 29.4000 115.8000 33.8000 116.1000 ;
	    RECT 39.0000 115.8000 39.4000 116.2000 ;
	    RECT 83.0000 116.1000 83.4000 116.2000 ;
	    RECT 85.4000 116.1000 85.8000 116.2000 ;
	    RECT 90.2000 116.1000 90.6000 116.2000 ;
	    RECT 83.0000 115.8000 90.6000 116.1000 ;
	    RECT 106.2000 116.1000 106.6000 116.2000 ;
	    RECT 108.6000 116.1000 109.0000 116.2000 ;
	    RECT 106.2000 115.8000 109.0000 116.1000 ;
	    RECT 134.2000 116.1000 134.5000 116.8000 ;
	    RECT 135.8000 116.1000 136.2000 116.2000 ;
	    RECT 134.2000 115.8000 136.2000 116.1000 ;
	    RECT 149.4000 116.1000 149.8000 116.2000 ;
	    RECT 151.8000 116.1000 152.1000 116.8000 ;
	    RECT 153.4000 116.1000 153.8000 116.2000 ;
	    RECT 149.4000 115.8000 153.8000 116.1000 ;
	    RECT 167.8000 116.1000 168.2000 116.2000 ;
	    RECT 182.2000 116.1000 182.6000 116.2000 ;
	    RECT 191.8000 116.1000 192.2000 116.2000 ;
	    RECT 167.8000 115.8000 192.2000 116.1000 ;
	    RECT 194.2000 116.1000 194.6000 116.2000 ;
	    RECT 204.6000 116.1000 205.0000 116.2000 ;
	    RECT 229.4000 116.1000 229.8000 116.2000 ;
	    RECT 194.2000 115.8000 205.0000 116.1000 ;
	    RECT 218.2000 115.8000 229.8000 116.1000 ;
	    RECT 231.0000 116.1000 231.4000 116.2000 ;
	    RECT 236.6000 116.1000 237.0000 116.2000 ;
	    RECT 231.0000 115.8000 237.0000 116.1000 ;
	    RECT 242.2000 116.1000 242.6000 116.2000 ;
	    RECT 247.0000 116.1000 247.4000 116.2000 ;
	    RECT 242.2000 115.8000 247.4000 116.1000 ;
	    RECT 253.4000 115.8000 253.8000 116.2000 ;
	    RECT 254.2000 115.8000 254.6000 116.2000 ;
	    RECT 258.2000 116.1000 258.6000 116.2000 ;
	    RECT 267.0000 116.1000 267.4000 116.2000 ;
	    RECT 258.2000 115.8000 267.4000 116.1000 ;
	    RECT 20.6000 115.1000 21.0000 115.2000 ;
	    RECT 23.8000 115.1000 24.2000 115.2000 ;
	    RECT 20.6000 114.8000 24.2000 115.1000 ;
	    RECT 31.0000 114.8000 31.4000 115.2000 ;
	    RECT 39.0000 115.1000 39.3000 115.8000 ;
	    RECT 218.2000 115.2000 218.5000 115.8000 ;
	    RECT 34.2000 114.8000 39.3000 115.1000 ;
	    RECT 54.2000 115.1000 54.6000 115.2000 ;
	    RECT 59.8000 115.1000 60.2000 115.2000 ;
	    RECT 54.2000 114.8000 60.2000 115.1000 ;
	    RECT 75.0000 115.1000 75.4000 115.2000 ;
	    RECT 75.8000 115.1000 76.2000 115.2000 ;
	    RECT 75.0000 114.8000 76.2000 115.1000 ;
	    RECT 88.6000 115.1000 89.0000 115.2000 ;
	    RECT 99.8000 115.1000 100.2000 115.2000 ;
	    RECT 112.6000 115.1000 113.0000 115.2000 ;
	    RECT 117.4000 115.1000 117.8000 115.2000 ;
	    RECT 133.4000 115.1000 133.8000 115.2000 ;
	    RECT 88.6000 114.8000 93.0000 115.1000 ;
	    RECT 99.8000 114.8000 117.8000 115.1000 ;
	    RECT 130.2000 114.8000 133.8000 115.1000 ;
	    RECT 135.0000 115.1000 135.4000 115.2000 ;
	    RECT 150.2000 115.1000 150.6000 115.2000 ;
	    RECT 135.0000 114.8000 150.6000 115.1000 ;
	    RECT 169.4000 115.1000 169.8000 115.2000 ;
	    RECT 179.0000 115.1000 179.4000 115.2000 ;
	    RECT 169.4000 114.8000 179.4000 115.1000 ;
	    RECT 180.6000 115.1000 181.0000 115.2000 ;
	    RECT 181.4000 115.1000 181.8000 115.2000 ;
	    RECT 180.6000 114.8000 181.8000 115.1000 ;
	    RECT 195.8000 114.8000 196.2000 115.2000 ;
	    RECT 200.6000 114.8000 201.0000 115.2000 ;
	    RECT 207.8000 115.1000 208.2000 115.2000 ;
	    RECT 211.8000 115.1000 212.2000 115.2000 ;
	    RECT 207.8000 114.8000 212.2000 115.1000 ;
	    RECT 218.2000 114.8000 218.6000 115.2000 ;
	    RECT 224.6000 114.8000 225.0000 115.2000 ;
	    RECT 225.4000 114.8000 225.8000 115.2000 ;
	    RECT 230.2000 115.1000 230.6000 115.2000 ;
	    RECT 235.8000 115.1000 236.2000 115.2000 ;
	    RECT 241.4000 115.1000 241.8000 115.2000 ;
	    RECT 246.2000 115.1000 246.6000 115.2000 ;
	    RECT 230.2000 114.8000 246.6000 115.1000 ;
	    RECT 248.6000 115.1000 249.0000 115.2000 ;
	    RECT 253.4000 115.1000 253.7000 115.8000 ;
	    RECT 248.6000 114.8000 253.7000 115.1000 ;
	    RECT 254.2000 115.1000 254.5000 115.8000 ;
	    RECT 263.0000 115.1000 263.4000 115.2000 ;
	    RECT 254.2000 114.8000 263.4000 115.1000 ;
	    RECT 31.0000 114.2000 31.3000 114.8000 ;
	    RECT 34.2000 114.2000 34.5000 114.8000 ;
	    RECT 92.6000 114.7000 93.0000 114.8000 ;
	    RECT 130.2000 114.2000 130.5000 114.8000 ;
	    RECT 195.8000 114.2000 196.1000 114.8000 ;
	    RECT 200.6000 114.2000 200.9000 114.8000 ;
	    RECT 6.2000 114.1000 6.6000 114.2000 ;
	    RECT 11.0000 114.1000 11.4000 114.2000 ;
	    RECT 6.2000 113.8000 11.4000 114.1000 ;
	    RECT 17.4000 113.8000 17.8000 114.2000 ;
	    RECT 27.0000 114.1000 27.4000 114.2000 ;
	    RECT 28.6000 114.1000 29.0000 114.2000 ;
	    RECT 21.4000 113.8000 29.0000 114.1000 ;
	    RECT 31.0000 113.8000 31.4000 114.2000 ;
	    RECT 34.2000 113.8000 34.6000 114.2000 ;
	    RECT 35.8000 114.1000 36.2000 114.2000 ;
	    RECT 47.0000 114.1000 47.4000 114.2000 ;
	    RECT 35.8000 113.8000 47.4000 114.1000 ;
	    RECT 63.0000 114.1000 63.4000 114.2000 ;
	    RECT 93.4000 114.1000 93.8000 114.2000 ;
	    RECT 102.2000 114.1000 102.6000 114.2000 ;
	    RECT 63.0000 113.8000 102.6000 114.1000 ;
	    RECT 105.4000 114.1000 105.8000 114.2000 ;
	    RECT 107.8000 114.1000 108.2000 114.2000 ;
	    RECT 116.6000 114.1000 117.0000 114.2000 ;
	    RECT 105.4000 113.8000 117.0000 114.1000 ;
	    RECT 126.2000 113.8000 126.6000 114.2000 ;
	    RECT 130.2000 113.8000 130.6000 114.2000 ;
	    RECT 131.8000 114.1000 132.2000 114.2000 ;
	    RECT 134.2000 114.1000 134.6000 114.2000 ;
	    RECT 131.8000 113.8000 134.6000 114.1000 ;
	    RECT 135.8000 114.1000 136.2000 114.2000 ;
	    RECT 136.6000 114.1000 137.0000 114.2000 ;
	    RECT 135.8000 113.8000 137.0000 114.1000 ;
	    RECT 140.6000 114.1000 141.0000 114.2000 ;
	    RECT 144.6000 114.1000 145.0000 114.2000 ;
	    RECT 140.6000 113.8000 145.0000 114.1000 ;
	    RECT 149.4000 114.1000 149.8000 114.2000 ;
	    RECT 163.0000 114.1000 163.4000 114.2000 ;
	    RECT 149.4000 113.8000 163.4000 114.1000 ;
	    RECT 179.8000 114.1000 180.2000 114.2000 ;
	    RECT 183.8000 114.1000 184.2000 114.2000 ;
	    RECT 179.8000 113.8000 184.2000 114.1000 ;
	    RECT 195.8000 113.8000 196.2000 114.2000 ;
	    RECT 200.6000 113.8000 201.0000 114.2000 ;
	    RECT 207.0000 114.1000 207.4000 114.2000 ;
	    RECT 215.8000 114.1000 216.2000 114.2000 ;
	    RECT 221.4000 114.1000 221.8000 114.2000 ;
	    RECT 207.0000 113.8000 221.8000 114.1000 ;
	    RECT 223.0000 114.1000 223.4000 114.2000 ;
	    RECT 224.6000 114.1000 224.9000 114.8000 ;
	    RECT 223.0000 113.8000 224.9000 114.1000 ;
	    RECT 225.4000 114.1000 225.7000 114.8000 ;
	    RECT 228.6000 114.1000 229.0000 114.2000 ;
	    RECT 225.4000 113.8000 229.0000 114.1000 ;
	    RECT 230.2000 114.1000 230.6000 114.2000 ;
	    RECT 231.0000 114.1000 231.4000 114.2000 ;
	    RECT 230.2000 113.8000 231.4000 114.1000 ;
	    RECT 235.0000 114.1000 235.4000 114.2000 ;
	    RECT 247.8000 114.1000 248.2000 114.2000 ;
	    RECT 235.0000 113.8000 248.2000 114.1000 ;
	    RECT 250.2000 114.1000 250.6000 114.2000 ;
	    RECT 251.0000 114.1000 251.4000 114.2000 ;
	    RECT 250.2000 113.8000 251.4000 114.1000 ;
	    RECT 258.2000 114.1000 258.6000 114.2000 ;
	    RECT 259.8000 114.1000 260.2000 114.2000 ;
	    RECT 258.2000 113.8000 260.2000 114.1000 ;
	    RECT 262.2000 114.1000 262.6000 114.2000 ;
	    RECT 266.2000 114.1000 266.6000 114.2000 ;
	    RECT 262.2000 113.8000 266.6000 114.1000 ;
	    RECT 17.4000 113.2000 17.7000 113.8000 ;
	    RECT 21.4000 113.2000 21.7000 113.8000 ;
	    RECT 17.4000 112.8000 17.8000 113.2000 ;
	    RECT 21.4000 112.8000 21.8000 113.2000 ;
	    RECT 26.2000 113.1000 26.6000 113.2000 ;
	    RECT 27.0000 113.1000 27.4000 113.2000 ;
	    RECT 26.2000 112.8000 27.4000 113.1000 ;
	    RECT 63.8000 113.1000 64.2000 113.2000 ;
	    RECT 87.0000 113.1000 87.4000 113.2000 ;
	    RECT 63.8000 112.8000 87.4000 113.1000 ;
	    RECT 87.8000 113.1000 88.2000 113.2000 ;
	    RECT 98.2000 113.1000 98.6000 113.2000 ;
	    RECT 110.2000 113.1000 110.6000 113.2000 ;
	    RECT 113.4000 113.1000 113.8000 113.2000 ;
	    RECT 87.8000 112.8000 99.3000 113.1000 ;
	    RECT 110.2000 112.8000 113.8000 113.1000 ;
	    RECT 124.6000 113.1000 125.0000 113.2000 ;
	    RECT 126.2000 113.1000 126.5000 113.8000 ;
	    RECT 132.6000 113.1000 133.0000 113.2000 ;
	    RECT 124.6000 112.8000 133.0000 113.1000 ;
	    RECT 133.4000 113.1000 133.8000 113.2000 ;
	    RECT 136.6000 113.1000 137.0000 113.2000 ;
	    RECT 133.4000 112.8000 137.0000 113.1000 ;
	    RECT 139.8000 113.1000 140.2000 113.2000 ;
	    RECT 141.4000 113.1000 141.8000 113.2000 ;
	    RECT 139.8000 112.8000 141.8000 113.1000 ;
	    RECT 147.0000 113.1000 147.4000 113.2000 ;
	    RECT 150.2000 113.1000 150.6000 113.2000 ;
	    RECT 147.0000 112.8000 150.6000 113.1000 ;
	    RECT 155.0000 112.8000 155.4000 113.2000 ;
	    RECT 163.8000 113.1000 164.2000 113.2000 ;
	    RECT 178.2000 113.1000 178.6000 113.2000 ;
	    RECT 163.8000 112.8000 178.6000 113.1000 ;
	    RECT 191.8000 113.1000 192.2000 113.2000 ;
	    RECT 193.4000 113.1000 193.8000 113.2000 ;
	    RECT 191.8000 112.8000 193.8000 113.1000 ;
	    RECT 203.8000 113.1000 204.2000 113.2000 ;
	    RECT 208.6000 113.1000 209.0000 113.2000 ;
	    RECT 218.2000 113.1000 218.6000 113.2000 ;
	    RECT 203.8000 112.8000 218.6000 113.1000 ;
	    RECT 220.6000 113.1000 221.0000 113.2000 ;
	    RECT 226.2000 113.1000 226.6000 113.2000 ;
	    RECT 239.0000 113.1000 239.4000 113.2000 ;
	    RECT 245.4000 113.1000 245.8000 113.2000 ;
	    RECT 250.2000 113.1000 250.6000 113.2000 ;
	    RECT 220.6000 112.8000 250.6000 113.1000 ;
	    RECT 256.6000 113.1000 257.0000 113.2000 ;
	    RECT 257.4000 113.1000 257.8000 113.2000 ;
	    RECT 256.6000 112.8000 257.8000 113.1000 ;
	    RECT 13.4000 112.1000 13.8000 112.2000 ;
	    RECT 27.8000 112.1000 28.2000 112.2000 ;
	    RECT 13.4000 111.8000 28.2000 112.1000 ;
	    RECT 59.8000 112.1000 60.2000 112.2000 ;
	    RECT 63.0000 112.1000 63.4000 112.2000 ;
	    RECT 59.8000 111.8000 63.4000 112.1000 ;
	    RECT 81.4000 112.1000 81.8000 112.2000 ;
	    RECT 90.2000 112.1000 90.6000 112.2000 ;
	    RECT 81.4000 111.8000 90.6000 112.1000 ;
	    RECT 99.0000 112.1000 99.4000 112.2000 ;
	    RECT 99.8000 112.1000 100.2000 112.2000 ;
	    RECT 99.0000 111.8000 100.2000 112.1000 ;
	    RECT 100.6000 112.1000 101.0000 112.2000 ;
	    RECT 115.0000 112.1000 115.4000 112.2000 ;
	    RECT 100.6000 111.8000 115.4000 112.1000 ;
	    RECT 144.6000 112.1000 145.0000 112.2000 ;
	    RECT 155.0000 112.1000 155.3000 112.8000 ;
	    RECT 144.6000 111.8000 155.3000 112.1000 ;
	    RECT 165.4000 112.1000 165.8000 112.2000 ;
	    RECT 174.2000 112.1000 174.6000 112.2000 ;
	    RECT 165.4000 111.8000 174.6000 112.1000 ;
	    RECT 185.4000 112.1000 185.8000 112.2000 ;
	    RECT 189.4000 112.1000 189.8000 112.2000 ;
	    RECT 185.4000 111.8000 189.8000 112.1000 ;
	    RECT 204.6000 112.1000 205.0000 112.2000 ;
	    RECT 209.4000 112.1000 209.8000 112.2000 ;
	    RECT 204.6000 111.8000 209.8000 112.1000 ;
	    RECT 210.2000 112.1000 210.6000 112.2000 ;
	    RECT 242.2000 112.1000 242.6000 112.2000 ;
	    RECT 247.0000 112.1000 247.4000 112.2000 ;
	    RECT 210.2000 111.8000 232.9000 112.1000 ;
	    RECT 242.2000 111.8000 247.4000 112.1000 ;
	    RECT 36.6000 111.1000 37.0000 111.2000 ;
	    RECT 63.0000 111.1000 63.4000 111.2000 ;
	    RECT 63.8000 111.1000 64.2000 111.2000 ;
	    RECT 36.6000 110.8000 64.2000 111.1000 ;
	    RECT 83.0000 111.1000 83.4000 111.2000 ;
	    RECT 84.6000 111.1000 85.0000 111.2000 ;
	    RECT 83.0000 110.8000 85.0000 111.1000 ;
	    RECT 90.2000 111.1000 90.6000 111.2000 ;
	    RECT 100.6000 111.1000 101.0000 111.2000 ;
	    RECT 90.2000 110.8000 101.0000 111.1000 ;
	    RECT 148.6000 111.1000 149.0000 111.2000 ;
	    RECT 173.4000 111.1000 173.8000 111.2000 ;
	    RECT 148.6000 110.8000 173.8000 111.1000 ;
	    RECT 187.0000 111.1000 187.4000 111.2000 ;
	    RECT 189.4000 111.1000 189.8000 111.2000 ;
	    RECT 187.0000 110.8000 189.8000 111.1000 ;
	    RECT 197.4000 111.1000 197.8000 111.2000 ;
	    RECT 199.8000 111.1000 200.2000 111.2000 ;
	    RECT 197.4000 110.8000 200.2000 111.1000 ;
	    RECT 222.2000 111.1000 222.6000 111.2000 ;
	    RECT 231.8000 111.1000 232.2000 111.2000 ;
	    RECT 222.2000 110.8000 232.2000 111.1000 ;
	    RECT 232.6000 111.1000 232.9000 111.8000 ;
	    RECT 243.0000 111.1000 243.4000 111.2000 ;
	    RECT 232.6000 110.8000 243.4000 111.1000 ;
	    RECT 243.8000 110.8000 244.2000 111.2000 ;
	    RECT 243.8000 110.2000 244.1000 110.8000 ;
	    RECT 63.8000 110.1000 64.2000 110.2000 ;
	    RECT 66.2000 110.1000 66.6000 110.2000 ;
	    RECT 77.4000 110.1000 77.8000 110.2000 ;
	    RECT 87.0000 110.1000 87.4000 110.2000 ;
	    RECT 63.8000 109.8000 87.4000 110.1000 ;
	    RECT 101.4000 110.1000 101.8000 110.2000 ;
	    RECT 107.0000 110.1000 107.4000 110.2000 ;
	    RECT 101.4000 109.8000 107.4000 110.1000 ;
	    RECT 138.2000 110.1000 138.6000 110.2000 ;
	    RECT 143.0000 110.1000 143.4000 110.2000 ;
	    RECT 138.2000 109.8000 143.4000 110.1000 ;
	    RECT 153.4000 110.1000 153.8000 110.2000 ;
	    RECT 155.8000 110.1000 156.2000 110.2000 ;
	    RECT 171.0000 110.1000 171.4000 110.2000 ;
	    RECT 153.4000 109.8000 171.4000 110.1000 ;
	    RECT 176.6000 110.1000 177.0000 110.2000 ;
	    RECT 178.2000 110.1000 178.6000 110.2000 ;
	    RECT 176.6000 109.8000 178.6000 110.1000 ;
	    RECT 183.8000 110.1000 184.2000 110.2000 ;
	    RECT 200.6000 110.1000 201.0000 110.2000 ;
	    RECT 183.8000 109.8000 201.0000 110.1000 ;
	    RECT 201.4000 110.1000 201.8000 110.2000 ;
	    RECT 207.0000 110.1000 207.4000 110.2000 ;
	    RECT 234.2000 110.1000 234.6000 110.2000 ;
	    RECT 201.4000 109.8000 207.4000 110.1000 ;
	    RECT 212.6000 109.8000 234.6000 110.1000 ;
	    RECT 243.8000 109.8000 244.2000 110.2000 ;
	    RECT 11.0000 109.1000 11.4000 109.2000 ;
	    RECT 18.2000 109.1000 18.6000 109.2000 ;
	    RECT 3.0000 108.8000 18.6000 109.1000 ;
	    RECT 30.2000 108.8000 30.6000 109.2000 ;
	    RECT 42.2000 109.1000 42.6000 109.2000 ;
	    RECT 52.6000 109.1000 53.0000 109.2000 ;
	    RECT 55.8000 109.1000 56.2000 109.2000 ;
	    RECT 59.8000 109.1000 60.2000 109.2000 ;
	    RECT 65.4000 109.1000 65.8000 109.2000 ;
	    RECT 41.4000 108.8000 65.8000 109.1000 ;
	    RECT 87.0000 109.1000 87.4000 109.2000 ;
	    RECT 111.0000 109.1000 111.4000 109.2000 ;
	    RECT 120.6000 109.1000 121.0000 109.2000 ;
	    RECT 87.0000 108.8000 121.0000 109.1000 ;
	    RECT 125.4000 109.1000 125.8000 109.2000 ;
	    RECT 134.2000 109.1000 134.6000 109.2000 ;
	    RECT 147.0000 109.1000 147.4000 109.2000 ;
	    RECT 125.4000 108.8000 147.4000 109.1000 ;
	    RECT 163.0000 108.8000 163.4000 109.2000 ;
	    RECT 172.6000 109.1000 173.0000 109.2000 ;
	    RECT 177.4000 109.1000 177.8000 109.2000 ;
	    RECT 172.6000 108.8000 177.8000 109.1000 ;
	    RECT 179.0000 109.1000 179.4000 109.2000 ;
	    RECT 184.6000 109.1000 185.0000 109.2000 ;
	    RECT 191.0000 109.1000 191.4000 109.2000 ;
	    RECT 200.6000 109.1000 201.0000 109.2000 ;
	    RECT 201.4000 109.1000 201.8000 109.2000 ;
	    RECT 179.0000 108.8000 201.8000 109.1000 ;
	    RECT 208.6000 109.1000 209.0000 109.2000 ;
	    RECT 212.6000 109.1000 212.9000 109.8000 ;
	    RECT 208.6000 108.8000 212.9000 109.1000 ;
	    RECT 221.4000 108.8000 221.8000 109.2000 ;
	    RECT 223.8000 109.1000 224.2000 109.2000 ;
	    RECT 229.4000 109.1000 229.8000 109.2000 ;
	    RECT 223.8000 108.8000 229.8000 109.1000 ;
	    RECT 230.2000 108.8000 230.6000 109.2000 ;
	    RECT 248.6000 109.1000 249.0000 109.2000 ;
	    RECT 252.6000 109.1000 253.0000 109.2000 ;
	    RECT 248.6000 108.8000 253.0000 109.1000 ;
	    RECT 3.0000 108.2000 3.3000 108.8000 ;
	    RECT 3.0000 107.8000 3.4000 108.2000 ;
	    RECT 3.8000 108.1000 4.2000 108.2000 ;
	    RECT 5.4000 108.1000 5.8000 108.2000 ;
	    RECT 3.8000 107.8000 5.8000 108.1000 ;
	    RECT 30.2000 108.1000 30.5000 108.8000 ;
	    RECT 37.4000 108.1000 37.8000 108.2000 ;
	    RECT 30.2000 107.8000 37.8000 108.1000 ;
	    RECT 45.4000 108.1000 45.8000 108.2000 ;
	    RECT 48.6000 108.1000 49.0000 108.2000 ;
	    RECT 45.4000 107.8000 49.0000 108.1000 ;
	    RECT 51.8000 108.1000 52.2000 108.2000 ;
	    RECT 67.8000 108.1000 68.2000 108.2000 ;
	    RECT 51.8000 107.8000 68.2000 108.1000 ;
	    RECT 78.2000 108.1000 78.6000 108.2000 ;
	    RECT 83.8000 108.1000 84.2000 108.2000 ;
	    RECT 78.2000 107.8000 84.2000 108.1000 ;
	    RECT 95.0000 108.1000 95.4000 108.2000 ;
	    RECT 100.6000 108.1000 101.0000 108.2000 ;
	    RECT 103.0000 108.1000 103.4000 108.2000 ;
	    RECT 95.0000 107.8000 103.4000 108.1000 ;
	    RECT 105.4000 108.1000 105.8000 108.2000 ;
	    RECT 130.2000 108.1000 130.6000 108.2000 ;
	    RECT 137.4000 108.1000 137.8000 108.2000 ;
	    RECT 105.4000 107.8000 119.3000 108.1000 ;
	    RECT 130.2000 107.8000 137.8000 108.1000 ;
	    RECT 143.0000 108.1000 143.4000 108.2000 ;
	    RECT 147.8000 108.1000 148.2000 108.2000 ;
	    RECT 143.0000 107.8000 148.2000 108.1000 ;
	    RECT 158.2000 108.1000 158.6000 108.2000 ;
	    RECT 163.0000 108.1000 163.3000 108.8000 ;
	    RECT 158.2000 107.8000 163.3000 108.1000 ;
	    RECT 171.0000 108.1000 171.4000 108.2000 ;
	    RECT 174.2000 108.1000 174.6000 108.2000 ;
	    RECT 171.0000 107.8000 174.6000 108.1000 ;
	    RECT 192.6000 108.1000 193.0000 108.2000 ;
	    RECT 201.4000 108.1000 201.8000 108.2000 ;
	    RECT 192.6000 107.8000 201.8000 108.1000 ;
	    RECT 202.2000 107.8000 202.6000 108.2000 ;
	    RECT 203.0000 108.1000 203.4000 108.2000 ;
	    RECT 203.8000 108.1000 204.2000 108.2000 ;
	    RECT 205.4000 108.1000 205.8000 108.2000 ;
	    RECT 203.0000 107.8000 205.8000 108.1000 ;
	    RECT 215.8000 107.8000 216.2000 108.2000 ;
	    RECT 216.6000 108.1000 217.0000 108.2000 ;
	    RECT 221.4000 108.1000 221.7000 108.8000 ;
	    RECT 216.6000 107.8000 221.7000 108.1000 ;
	    RECT 230.2000 108.1000 230.5000 108.8000 ;
	    RECT 231.8000 108.1000 232.2000 108.2000 ;
	    RECT 234.2000 108.1000 234.6000 108.2000 ;
	    RECT 230.2000 107.8000 234.6000 108.1000 ;
	    RECT 119.0000 107.2000 119.3000 107.8000 ;
	    RECT 174.2000 107.2000 174.5000 107.8000 ;
	    RECT 1.4000 107.1000 1.8000 107.2000 ;
	    RECT 4.6000 107.1000 5.0000 107.2000 ;
	    RECT 1.4000 106.8000 5.0000 107.1000 ;
	    RECT 8.6000 107.1000 9.0000 107.2000 ;
	    RECT 11.0000 107.1000 11.4000 107.2000 ;
	    RECT 8.6000 106.8000 11.4000 107.1000 ;
	    RECT 30.2000 106.8000 30.6000 107.2000 ;
	    RECT 42.2000 107.1000 42.6000 107.2000 ;
	    RECT 45.4000 107.1000 45.8000 107.2000 ;
	    RECT 55.0000 107.1000 55.4000 107.2000 ;
	    RECT 58.2000 107.1000 58.6000 107.2000 ;
	    RECT 42.2000 106.8000 45.8000 107.1000 ;
	    RECT 54.2000 106.8000 58.6000 107.1000 ;
	    RECT 83.0000 107.1000 83.4000 107.2000 ;
	    RECT 88.6000 107.1000 89.0000 107.2000 ;
	    RECT 90.2000 107.1000 90.6000 107.2000 ;
	    RECT 83.0000 106.8000 90.6000 107.1000 ;
	    RECT 95.8000 107.1000 96.2000 107.2000 ;
	    RECT 97.4000 107.1000 97.8000 107.2000 ;
	    RECT 95.8000 106.8000 97.8000 107.1000 ;
	    RECT 99.0000 107.1000 99.4000 107.2000 ;
	    RECT 103.8000 107.1000 104.2000 107.2000 ;
	    RECT 107.0000 107.1000 107.4000 107.2000 ;
	    RECT 99.0000 106.8000 107.4000 107.1000 ;
	    RECT 107.8000 107.1000 108.2000 107.2000 ;
	    RECT 118.2000 107.1000 118.6000 107.2000 ;
	    RECT 107.8000 106.8000 118.6000 107.1000 ;
	    RECT 119.0000 106.8000 119.4000 107.2000 ;
	    RECT 123.8000 107.1000 124.2000 107.2000 ;
	    RECT 124.6000 107.1000 125.0000 107.2000 ;
	    RECT 123.8000 106.8000 125.0000 107.1000 ;
	    RECT 136.6000 106.8000 137.0000 107.2000 ;
	    RECT 163.0000 107.1000 163.4000 107.2000 ;
	    RECT 166.2000 107.1000 166.6000 107.2000 ;
	    RECT 167.0000 107.1000 167.4000 107.2000 ;
	    RECT 163.0000 106.8000 167.4000 107.1000 ;
	    RECT 170.2000 107.1000 170.6000 107.2000 ;
	    RECT 171.8000 107.1000 172.2000 107.2000 ;
	    RECT 170.2000 106.8000 172.2000 107.1000 ;
	    RECT 174.2000 106.8000 174.6000 107.2000 ;
	    RECT 177.4000 107.1000 177.8000 107.2000 ;
	    RECT 178.2000 107.1000 178.6000 107.2000 ;
	    RECT 177.4000 106.8000 178.6000 107.1000 ;
	    RECT 182.2000 107.1000 182.6000 107.2000 ;
	    RECT 183.0000 107.1000 183.4000 107.2000 ;
	    RECT 182.2000 106.8000 183.4000 107.1000 ;
	    RECT 191.0000 107.1000 191.4000 107.2000 ;
	    RECT 202.2000 107.1000 202.5000 107.8000 ;
	    RECT 204.6000 107.1000 205.0000 107.2000 ;
	    RECT 191.0000 106.8000 205.0000 107.1000 ;
	    RECT 207.0000 107.1000 207.4000 107.2000 ;
	    RECT 209.4000 107.1000 209.8000 107.2000 ;
	    RECT 207.0000 106.8000 209.8000 107.1000 ;
	    RECT 215.8000 107.1000 216.1000 107.8000 ;
	    RECT 218.2000 107.1000 218.6000 107.2000 ;
	    RECT 215.8000 106.8000 218.6000 107.1000 ;
	    RECT 222.2000 106.8000 222.6000 107.2000 ;
	    RECT 224.6000 107.1000 225.0000 107.2000 ;
	    RECT 227.0000 107.1000 227.4000 107.2000 ;
	    RECT 230.2000 107.1000 230.6000 107.2000 ;
	    RECT 224.6000 106.8000 230.6000 107.1000 ;
	    RECT 261.4000 107.1000 261.8000 107.2000 ;
	    RECT 266.2000 107.1000 266.6000 107.2000 ;
	    RECT 261.4000 106.8000 266.6000 107.1000 ;
	    RECT 6.2000 106.1000 6.6000 106.2000 ;
	    RECT 5.4000 105.8000 6.6000 106.1000 ;
	    RECT 9.4000 106.1000 9.8000 106.2000 ;
	    RECT 10.2000 106.1000 10.6000 106.2000 ;
	    RECT 9.4000 105.8000 10.6000 106.1000 ;
	    RECT 15.8000 105.8000 16.2000 106.2000 ;
	    RECT 21.4000 106.1000 21.8000 106.2000 ;
	    RECT 22.2000 106.1000 22.6000 106.2000 ;
	    RECT 21.4000 105.8000 22.6000 106.1000 ;
	    RECT 30.2000 106.1000 30.5000 106.8000 ;
	    RECT 35.0000 106.1000 35.4000 106.2000 ;
	    RECT 30.2000 105.8000 35.4000 106.1000 ;
	    RECT 41.4000 106.1000 41.8000 106.2000 ;
	    RECT 47.8000 106.1000 48.2000 106.2000 ;
	    RECT 77.4000 106.1000 77.8000 106.2000 ;
	    RECT 113.4000 106.1000 113.8000 106.2000 ;
	    RECT 41.4000 105.8000 48.2000 106.1000 ;
	    RECT 74.2000 105.8000 77.8000 106.1000 ;
	    RECT 80.6000 105.8000 113.8000 106.1000 ;
	    RECT 115.8000 106.1000 116.2000 106.2000 ;
	    RECT 122.2000 106.1000 122.6000 106.2000 ;
	    RECT 115.8000 105.8000 122.6000 106.1000 ;
	    RECT 129.4000 106.1000 129.8000 106.2000 ;
	    RECT 136.6000 106.1000 136.9000 106.8000 ;
	    RECT 129.4000 105.8000 136.9000 106.1000 ;
	    RECT 139.0000 106.1000 139.4000 106.3000 ;
	    RECT 222.2000 106.2000 222.5000 106.8000 ;
	    RECT 143.8000 106.1000 144.2000 106.2000 ;
	    RECT 139.0000 105.8000 144.2000 106.1000 ;
	    RECT 150.2000 106.1000 150.6000 106.2000 ;
	    RECT 162.2000 106.1000 162.6000 106.2000 ;
	    RECT 150.2000 105.8000 162.6000 106.1000 ;
	    RECT 165.4000 106.1000 165.8000 106.2000 ;
	    RECT 169.4000 106.1000 169.8000 106.2000 ;
	    RECT 170.2000 106.1000 170.6000 106.2000 ;
	    RECT 178.2000 106.1000 178.6000 106.2000 ;
	    RECT 165.4000 105.8000 178.6000 106.1000 ;
	    RECT 182.2000 106.1000 182.6000 106.2000 ;
	    RECT 184.6000 106.1000 185.0000 106.2000 ;
	    RECT 195.8000 106.1000 196.2000 106.2000 ;
	    RECT 206.2000 106.1000 206.6000 106.2000 ;
	    RECT 182.2000 105.8000 206.6000 106.1000 ;
	    RECT 211.8000 106.1000 212.2000 106.2000 ;
	    RECT 215.8000 106.1000 216.2000 106.2000 ;
	    RECT 219.8000 106.1000 220.2000 106.2000 ;
	    RECT 220.6000 106.1000 221.0000 106.2000 ;
	    RECT 211.8000 105.8000 218.5000 106.1000 ;
	    RECT 219.8000 105.8000 221.0000 106.1000 ;
	    RECT 222.2000 105.8000 222.6000 106.2000 ;
	    RECT 231.0000 106.1000 231.4000 106.2000 ;
	    RECT 231.8000 106.1000 232.2000 106.2000 ;
	    RECT 231.0000 105.8000 232.2000 106.1000 ;
	    RECT 233.4000 105.8000 233.8000 106.2000 ;
	    RECT 235.0000 106.1000 235.4000 106.2000 ;
	    RECT 247.0000 106.1000 247.4000 106.2000 ;
	    RECT 235.0000 105.8000 247.4000 106.1000 ;
	    RECT 247.8000 105.8000 248.2000 106.2000 ;
	    RECT 255.8000 106.1000 256.2000 106.2000 ;
	    RECT 264.6000 106.1000 265.0000 106.2000 ;
	    RECT 255.8000 105.8000 265.0000 106.1000 ;
	    RECT 3.8000 105.1000 4.2000 105.2000 ;
	    RECT 5.4000 105.1000 5.7000 105.8000 ;
	    RECT 3.8000 104.8000 5.7000 105.1000 ;
	    RECT 6.2000 105.1000 6.6000 105.2000 ;
	    RECT 15.8000 105.1000 16.1000 105.8000 ;
	    RECT 74.2000 105.2000 74.5000 105.8000 ;
	    RECT 80.6000 105.2000 80.9000 105.8000 ;
	    RECT 6.2000 104.8000 16.1000 105.1000 ;
	    RECT 51.0000 105.1000 51.4000 105.2000 ;
	    RECT 53.4000 105.1000 53.8000 105.2000 ;
	    RECT 51.0000 104.8000 53.8000 105.1000 ;
	    RECT 74.2000 104.8000 74.6000 105.2000 ;
	    RECT 80.6000 104.8000 81.0000 105.2000 ;
	    RECT 82.2000 105.1000 82.6000 105.2000 ;
	    RECT 89.4000 105.1000 89.8000 105.2000 ;
	    RECT 82.2000 104.8000 89.8000 105.1000 ;
	    RECT 91.0000 105.1000 91.4000 105.2000 ;
	    RECT 95.8000 105.1000 96.2000 105.2000 ;
	    RECT 91.0000 104.8000 96.2000 105.1000 ;
	    RECT 97.4000 105.1000 97.8000 105.2000 ;
	    RECT 100.6000 105.1000 101.0000 105.2000 ;
	    RECT 97.4000 104.8000 101.0000 105.1000 ;
	    RECT 111.8000 104.8000 112.2000 105.2000 ;
	    RECT 119.8000 105.1000 120.2000 105.2000 ;
	    RECT 121.4000 105.1000 121.8000 105.2000 ;
	    RECT 119.8000 104.8000 121.8000 105.1000 ;
	    RECT 141.4000 105.1000 141.8000 105.2000 ;
	    RECT 144.6000 105.1000 145.0000 105.2000 ;
	    RECT 141.4000 104.8000 145.0000 105.1000 ;
	    RECT 155.0000 105.1000 155.4000 105.2000 ;
	    RECT 163.8000 105.1000 164.2000 105.2000 ;
	    RECT 155.0000 104.8000 164.2000 105.1000 ;
	    RECT 167.8000 105.1000 168.2000 105.2000 ;
	    RECT 171.0000 105.1000 171.4000 105.2000 ;
	    RECT 167.8000 104.8000 171.4000 105.1000 ;
	    RECT 175.0000 104.8000 175.4000 105.2000 ;
	    RECT 181.4000 105.1000 181.8000 105.2000 ;
	    RECT 182.2000 105.1000 182.6000 105.2000 ;
	    RECT 193.4000 105.1000 193.8000 105.2000 ;
	    RECT 195.8000 105.1000 196.2000 105.2000 ;
	    RECT 181.4000 104.8000 183.3000 105.1000 ;
	    RECT 193.4000 104.8000 196.2000 105.1000 ;
	    RECT 200.6000 105.1000 201.0000 105.2000 ;
	    RECT 217.4000 105.1000 217.8000 105.2000 ;
	    RECT 200.6000 104.8000 217.8000 105.1000 ;
	    RECT 218.2000 105.1000 218.5000 105.8000 ;
	    RECT 233.4000 105.1000 233.7000 105.8000 ;
	    RECT 218.2000 104.8000 233.7000 105.1000 ;
	    RECT 247.8000 105.1000 248.1000 105.8000 ;
	    RECT 260.6000 105.1000 261.0000 105.2000 ;
	    RECT 247.8000 104.8000 261.0000 105.1000 ;
	    RECT 7.8000 104.1000 8.2000 104.2000 ;
	    RECT 12.6000 104.1000 13.0000 104.2000 ;
	    RECT 7.8000 103.8000 13.0000 104.1000 ;
	    RECT 13.4000 104.1000 13.8000 104.2000 ;
	    RECT 14.2000 104.1000 14.6000 104.2000 ;
	    RECT 13.4000 103.8000 14.6000 104.1000 ;
	    RECT 24.6000 104.1000 25.0000 104.2000 ;
	    RECT 33.4000 104.1000 33.8000 104.2000 ;
	    RECT 35.8000 104.1000 36.2000 104.2000 ;
	    RECT 24.6000 103.8000 36.2000 104.1000 ;
	    RECT 55.0000 104.1000 55.4000 104.2000 ;
	    RECT 61.4000 104.1000 61.8000 104.2000 ;
	    RECT 68.6000 104.1000 69.0000 104.2000 ;
	    RECT 80.6000 104.1000 80.9000 104.8000 ;
	    RECT 55.0000 103.8000 80.9000 104.1000 ;
	    RECT 84.6000 104.1000 85.0000 104.2000 ;
	    RECT 86.2000 104.1000 86.6000 104.2000 ;
	    RECT 84.6000 103.8000 86.6000 104.1000 ;
	    RECT 107.8000 104.1000 108.2000 104.2000 ;
	    RECT 111.8000 104.1000 112.1000 104.8000 ;
	    RECT 107.8000 103.8000 112.1000 104.1000 ;
	    RECT 116.6000 104.1000 117.0000 104.2000 ;
	    RECT 127.8000 104.1000 128.2000 104.2000 ;
	    RECT 116.6000 103.8000 128.2000 104.1000 ;
	    RECT 175.0000 104.1000 175.3000 104.8000 ;
	    RECT 175.8000 104.1000 176.2000 104.2000 ;
	    RECT 175.0000 103.8000 176.2000 104.1000 ;
	    RECT 187.8000 104.1000 188.2000 104.2000 ;
	    RECT 207.0000 104.1000 207.4000 104.2000 ;
	    RECT 187.8000 103.8000 207.4000 104.1000 ;
	    RECT 223.0000 104.1000 223.4000 104.2000 ;
	    RECT 223.8000 104.1000 224.2000 104.2000 ;
	    RECT 239.8000 104.1000 240.2000 104.2000 ;
	    RECT 255.0000 104.1000 255.4000 104.2000 ;
	    RECT 223.0000 103.8000 240.2000 104.1000 ;
	    RECT 249.4000 103.8000 255.4000 104.1000 ;
	    RECT 263.0000 104.1000 263.4000 104.2000 ;
	    RECT 267.0000 104.1000 267.4000 104.2000 ;
	    RECT 263.0000 103.8000 267.4000 104.1000 ;
	    RECT 249.4000 103.2000 249.7000 103.8000 ;
	    RECT 23.8000 103.1000 24.2000 103.2000 ;
	    RECT 31.8000 103.1000 32.2000 103.2000 ;
	    RECT 23.8000 102.8000 32.2000 103.1000 ;
	    RECT 115.0000 103.1000 115.4000 103.2000 ;
	    RECT 124.6000 103.1000 125.0000 103.2000 ;
	    RECT 115.0000 102.8000 125.0000 103.1000 ;
	    RECT 249.4000 102.8000 249.8000 103.2000 ;
	    RECT 58.2000 102.1000 58.6000 102.2000 ;
	    RECT 94.2000 102.1000 94.6000 102.2000 ;
	    RECT 58.2000 101.8000 94.6000 102.1000 ;
	    RECT 108.6000 102.1000 109.0000 102.2000 ;
	    RECT 118.2000 102.1000 118.6000 102.2000 ;
	    RECT 108.6000 101.8000 118.6000 102.1000 ;
	    RECT 243.8000 101.8000 244.2000 102.2000 ;
	    RECT 247.8000 102.1000 248.2000 102.2000 ;
	    RECT 258.2000 102.1000 258.6000 102.2000 ;
	    RECT 247.8000 101.8000 258.6000 102.1000 ;
	    RECT 243.8000 101.2000 244.1000 101.8000 ;
	    RECT 83.8000 101.1000 84.2000 101.2000 ;
	    RECT 102.2000 101.1000 102.6000 101.2000 ;
	    RECT 83.8000 100.8000 102.6000 101.1000 ;
	    RECT 243.8000 100.8000 244.2000 101.2000 ;
	    RECT 98.2000 99.8000 98.6000 100.2000 ;
	    RECT 189.4000 100.1000 189.8000 100.2000 ;
	    RECT 230.2000 100.1000 230.6000 100.2000 ;
	    RECT 235.8000 100.1000 236.2000 100.2000 ;
	    RECT 247.0000 100.1000 247.4000 100.2000 ;
	    RECT 189.4000 99.8000 247.4000 100.1000 ;
	    RECT 98.2000 99.2000 98.5000 99.8000 ;
	    RECT 63.8000 99.1000 64.2000 99.2000 ;
	    RECT 75.0000 99.1000 75.4000 99.2000 ;
	    RECT 63.8000 98.8000 75.4000 99.1000 ;
	    RECT 98.2000 98.8000 98.6000 99.2000 ;
	    RECT 200.6000 99.1000 201.0000 99.2000 ;
	    RECT 203.8000 99.1000 204.2000 99.2000 ;
	    RECT 200.6000 98.8000 204.2000 99.1000 ;
	    RECT 66.2000 98.1000 66.6000 98.2000 ;
	    RECT 77.4000 98.1000 77.8000 98.2000 ;
	    RECT 98.2000 98.1000 98.6000 98.2000 ;
	    RECT 100.6000 98.1000 101.0000 98.2000 ;
	    RECT 66.2000 97.8000 101.0000 98.1000 ;
	    RECT 103.8000 97.8000 104.2000 98.2000 ;
	    RECT 161.4000 97.8000 161.8000 98.2000 ;
	    RECT 177.4000 98.1000 177.8000 98.2000 ;
	    RECT 182.2000 98.1000 182.6000 98.2000 ;
	    RECT 186.2000 98.1000 186.6000 98.2000 ;
	    RECT 191.8000 98.1000 192.2000 98.2000 ;
	    RECT 177.4000 97.8000 192.2000 98.1000 ;
	    RECT 223.8000 98.1000 224.2000 98.2000 ;
	    RECT 266.2000 98.1000 266.6000 98.2000 ;
	    RECT 223.8000 97.8000 266.6000 98.1000 ;
	    RECT 103.8000 97.2000 104.1000 97.8000 ;
	    RECT 36.6000 96.8000 37.0000 97.2000 ;
	    RECT 74.2000 97.1000 74.6000 97.2000 ;
	    RECT 81.4000 97.1000 81.8000 97.2000 ;
	    RECT 84.6000 97.1000 85.0000 97.2000 ;
	    RECT 74.2000 96.8000 87.3000 97.1000 ;
	    RECT 103.8000 96.8000 104.2000 97.2000 ;
	    RECT 142.2000 97.1000 142.6000 97.2000 ;
	    RECT 145.4000 97.1000 145.8000 97.2000 ;
	    RECT 146.2000 97.1000 146.6000 97.2000 ;
	    RECT 142.2000 96.8000 146.6000 97.1000 ;
	    RECT 161.4000 97.1000 161.7000 97.8000 ;
	    RECT 164.6000 97.1000 165.0000 97.2000 ;
	    RECT 175.0000 97.1000 175.4000 97.2000 ;
	    RECT 161.4000 96.8000 175.4000 97.1000 ;
	    RECT 185.4000 96.8000 185.8000 97.2000 ;
	    RECT 187.0000 96.8000 187.4000 97.2000 ;
	    RECT 205.4000 97.1000 205.8000 97.2000 ;
	    RECT 206.2000 97.1000 206.6000 97.2000 ;
	    RECT 211.0000 97.1000 211.4000 97.2000 ;
	    RECT 205.4000 96.8000 211.4000 97.1000 ;
	    RECT 231.0000 96.8000 231.4000 97.2000 ;
	    RECT 239.0000 97.1000 239.4000 97.2000 ;
	    RECT 246.2000 97.1000 246.6000 97.2000 ;
	    RECT 239.0000 96.8000 246.6000 97.1000 ;
	    RECT 250.2000 97.1000 250.6000 97.2000 ;
	    RECT 264.6000 97.1000 265.0000 97.2000 ;
	    RECT 250.2000 96.8000 265.0000 97.1000 ;
	    RECT 1.4000 96.1000 1.8000 96.2000 ;
	    RECT 11.0000 96.1000 11.4000 96.2000 ;
	    RECT 1.4000 95.8000 11.4000 96.1000 ;
	    RECT 23.0000 96.1000 23.4000 96.2000 ;
	    RECT 28.6000 96.1000 29.0000 96.2000 ;
	    RECT 23.0000 95.8000 29.0000 96.1000 ;
	    RECT 36.6000 96.1000 36.9000 96.8000 ;
	    RECT 87.0000 96.2000 87.3000 96.8000 ;
	    RECT 43.0000 96.1000 43.4000 96.2000 ;
	    RECT 36.6000 95.8000 43.4000 96.1000 ;
	    RECT 47.0000 96.1000 47.4000 96.2000 ;
	    RECT 50.2000 96.1000 50.6000 96.2000 ;
	    RECT 47.0000 95.8000 50.6000 96.1000 ;
	    RECT 61.4000 96.1000 61.8000 96.2000 ;
	    RECT 72.6000 96.1000 73.0000 96.2000 ;
	    RECT 61.4000 95.8000 73.0000 96.1000 ;
	    RECT 87.0000 95.8000 87.4000 96.2000 ;
	    RECT 95.0000 95.8000 95.4000 96.2000 ;
	    RECT 97.4000 95.8000 97.8000 96.2000 ;
	    RECT 139.8000 96.1000 140.2000 96.2000 ;
	    RECT 140.6000 96.1000 141.0000 96.2000 ;
	    RECT 139.8000 95.8000 141.0000 96.1000 ;
	    RECT 168.6000 96.1000 169.0000 96.2000 ;
	    RECT 169.4000 96.1000 169.8000 96.2000 ;
	    RECT 168.6000 95.8000 169.8000 96.1000 ;
	    RECT 185.4000 96.1000 185.7000 96.8000 ;
	    RECT 187.0000 96.1000 187.3000 96.8000 ;
	    RECT 185.4000 95.8000 187.3000 96.1000 ;
	    RECT 204.6000 96.1000 205.0000 96.2000 ;
	    RECT 209.4000 96.1000 209.8000 96.2000 ;
	    RECT 225.4000 96.1000 225.8000 96.2000 ;
	    RECT 204.6000 95.8000 225.8000 96.1000 ;
	    RECT 227.8000 96.1000 228.2000 96.2000 ;
	    RECT 231.0000 96.1000 231.3000 96.8000 ;
	    RECT 227.8000 95.8000 231.3000 96.1000 ;
	    RECT 235.0000 96.1000 235.4000 96.2000 ;
	    RECT 235.8000 96.1000 236.2000 96.2000 ;
	    RECT 235.0000 95.8000 236.2000 96.1000 ;
	    RECT 240.6000 96.1000 241.0000 96.2000 ;
	    RECT 249.4000 96.1000 249.8000 96.2000 ;
	    RECT 240.6000 95.8000 249.8000 96.1000 ;
	    RECT 95.0000 95.2000 95.3000 95.8000 ;
	    RECT 11.8000 95.1000 12.2000 95.2000 ;
	    RECT 14.2000 95.1000 14.6000 95.2000 ;
	    RECT 9.4000 94.8000 14.6000 95.1000 ;
	    RECT 24.6000 95.1000 25.0000 95.2000 ;
	    RECT 25.4000 95.1000 25.8000 95.2000 ;
	    RECT 24.6000 94.8000 25.8000 95.1000 ;
	    RECT 40.6000 95.1000 41.0000 95.2000 ;
	    RECT 48.6000 95.1000 49.0000 95.2000 ;
	    RECT 49.4000 95.1000 49.8000 95.2000 ;
	    RECT 40.6000 94.8000 49.8000 95.1000 ;
	    RECT 50.2000 94.8000 50.6000 95.2000 ;
	    RECT 51.0000 95.1000 51.4000 95.2000 ;
	    RECT 72.6000 95.1000 73.0000 95.2000 ;
	    RECT 75.0000 95.1000 75.4000 95.2000 ;
	    RECT 51.0000 94.8000 65.8000 95.1000 ;
	    RECT 72.6000 94.8000 75.4000 95.1000 ;
	    RECT 88.6000 94.8000 89.0000 95.2000 ;
	    RECT 95.0000 94.8000 95.4000 95.2000 ;
	    RECT 97.4000 95.1000 97.7000 95.8000 ;
	    RECT 101.4000 95.1000 101.8000 95.2000 ;
	    RECT 97.4000 94.8000 101.8000 95.1000 ;
	    RECT 111.0000 95.1000 111.4000 95.2000 ;
	    RECT 124.6000 95.1000 125.0000 95.2000 ;
	    RECT 111.0000 94.8000 117.7000 95.1000 ;
	    RECT 9.4000 94.2000 9.7000 94.8000 ;
	    RECT 50.2000 94.2000 50.5000 94.8000 ;
	    RECT 65.4000 94.7000 65.8000 94.8000 ;
	    RECT 88.6000 94.2000 88.9000 94.8000 ;
	    RECT 117.4000 94.2000 117.7000 94.8000 ;
	    RECT 120.6000 94.8000 125.0000 95.1000 ;
	    RECT 158.2000 95.1000 158.6000 95.2000 ;
	    RECT 163.8000 95.1000 164.2000 95.2000 ;
	    RECT 158.2000 94.8000 164.2000 95.1000 ;
	    RECT 168.6000 95.1000 169.0000 95.2000 ;
	    RECT 171.8000 95.1000 172.2000 95.2000 ;
	    RECT 168.6000 94.8000 172.2000 95.1000 ;
	    RECT 183.0000 95.1000 183.4000 95.2000 ;
	    RECT 190.2000 95.1000 190.6000 95.2000 ;
	    RECT 207.0000 95.1000 207.4000 95.2000 ;
	    RECT 183.0000 94.8000 207.4000 95.1000 ;
	    RECT 215.8000 94.8000 216.2000 95.2000 ;
	    RECT 222.2000 95.1000 222.6000 95.2000 ;
	    RECT 239.8000 95.1000 240.2000 95.2000 ;
	    RECT 240.6000 95.1000 241.0000 95.2000 ;
	    RECT 222.2000 94.8000 241.0000 95.1000 ;
	    RECT 241.4000 95.1000 241.8000 95.2000 ;
	    RECT 253.4000 95.1000 253.8000 95.2000 ;
	    RECT 241.4000 94.8000 253.8000 95.1000 ;
	    RECT 120.6000 94.2000 120.9000 94.8000 ;
	    RECT 215.8000 94.2000 216.1000 94.8000 ;
	    RECT 9.4000 93.8000 9.8000 94.2000 ;
	    RECT 22.2000 94.1000 22.6000 94.2000 ;
	    RECT 24.6000 94.1000 25.0000 94.2000 ;
	    RECT 26.2000 94.1000 26.6000 94.2000 ;
	    RECT 22.2000 93.8000 23.3000 94.1000 ;
	    RECT 24.6000 93.8000 26.6000 94.1000 ;
	    RECT 35.8000 94.1000 36.2000 94.2000 ;
	    RECT 36.6000 94.1000 37.0000 94.2000 ;
	    RECT 35.8000 93.8000 37.0000 94.1000 ;
	    RECT 47.0000 93.8000 47.4000 94.2000 ;
	    RECT 50.2000 93.8000 50.6000 94.2000 ;
	    RECT 52.6000 94.1000 53.0000 94.2000 ;
	    RECT 53.4000 94.1000 53.8000 94.2000 ;
	    RECT 79.0000 94.1000 79.4000 94.2000 ;
	    RECT 52.6000 93.8000 79.4000 94.1000 ;
	    RECT 88.6000 93.8000 89.0000 94.2000 ;
	    RECT 93.4000 93.8000 93.8000 94.2000 ;
	    RECT 99.8000 94.1000 100.2000 94.2000 ;
	    RECT 106.2000 94.1000 106.6000 94.2000 ;
	    RECT 99.8000 93.8000 106.6000 94.1000 ;
	    RECT 109.4000 94.1000 109.8000 94.2000 ;
	    RECT 113.4000 94.1000 113.8000 94.2000 ;
	    RECT 109.4000 93.8000 113.8000 94.1000 ;
	    RECT 117.4000 93.8000 117.8000 94.2000 ;
	    RECT 120.6000 93.8000 121.0000 94.2000 ;
	    RECT 138.2000 93.8000 138.6000 94.2000 ;
	    RECT 139.8000 94.1000 140.2000 94.2000 ;
	    RECT 152.6000 94.1000 153.0000 94.2000 ;
	    RECT 166.2000 94.1000 166.6000 94.2000 ;
	    RECT 169.4000 94.1000 169.8000 94.2000 ;
	    RECT 139.8000 93.8000 144.1000 94.1000 ;
	    RECT 152.6000 93.8000 155.3000 94.1000 ;
	    RECT 166.2000 93.8000 169.8000 94.1000 ;
	    RECT 177.4000 94.1000 177.8000 94.2000 ;
	    RECT 189.4000 94.1000 189.8000 94.2000 ;
	    RECT 177.4000 93.8000 189.8000 94.1000 ;
	    RECT 200.6000 93.8000 201.0000 94.2000 ;
	    RECT 206.2000 94.1000 206.6000 94.2000 ;
	    RECT 209.4000 94.1000 209.8000 94.2000 ;
	    RECT 206.2000 93.8000 209.8000 94.1000 ;
	    RECT 215.8000 93.8000 216.2000 94.2000 ;
	    RECT 233.4000 94.1000 233.8000 94.2000 ;
	    RECT 235.0000 94.1000 235.4000 94.2000 ;
	    RECT 237.4000 94.1000 237.8000 94.2000 ;
	    RECT 233.4000 93.8000 237.8000 94.1000 ;
	    RECT 239.0000 94.1000 239.4000 94.2000 ;
	    RECT 248.6000 94.1000 249.0000 94.2000 ;
	    RECT 239.0000 93.8000 249.0000 94.1000 ;
	    RECT 23.0000 93.2000 23.3000 93.8000 ;
	    RECT 7.8000 93.1000 8.2000 93.2000 ;
	    RECT 13.4000 93.1000 13.8000 93.2000 ;
	    RECT 7.8000 92.8000 13.8000 93.1000 ;
	    RECT 23.0000 92.8000 23.4000 93.2000 ;
	    RECT 43.8000 93.1000 44.2000 93.2000 ;
	    RECT 47.0000 93.1000 47.3000 93.8000 ;
	    RECT 43.8000 92.8000 47.3000 93.1000 ;
	    RECT 47.8000 93.1000 48.2000 93.2000 ;
	    RECT 55.0000 93.1000 55.4000 93.2000 ;
	    RECT 55.8000 93.1000 56.2000 93.2000 ;
	    RECT 47.8000 92.8000 56.2000 93.1000 ;
	    RECT 59.8000 93.1000 60.2000 93.2000 ;
	    RECT 60.6000 93.1000 61.0000 93.2000 ;
	    RECT 59.8000 92.8000 61.0000 93.1000 ;
	    RECT 81.4000 93.1000 81.8000 93.2000 ;
	    RECT 84.6000 93.1000 85.0000 93.2000 ;
	    RECT 93.4000 93.1000 93.7000 93.8000 ;
	    RECT 138.2000 93.2000 138.5000 93.8000 ;
	    RECT 143.8000 93.2000 144.1000 93.8000 ;
	    RECT 155.0000 93.2000 155.3000 93.8000 ;
	    RECT 200.6000 93.2000 200.9000 93.8000 ;
	    RECT 81.4000 92.8000 93.7000 93.1000 ;
	    RECT 96.6000 93.1000 97.0000 93.2000 ;
	    RECT 98.2000 93.1000 98.6000 93.2000 ;
	    RECT 96.6000 92.8000 98.6000 93.1000 ;
	    RECT 138.2000 92.8000 138.6000 93.2000 ;
	    RECT 142.2000 93.1000 142.6000 93.2000 ;
	    RECT 143.0000 93.1000 143.4000 93.2000 ;
	    RECT 142.2000 92.8000 143.4000 93.1000 ;
	    RECT 143.8000 92.8000 144.2000 93.2000 ;
	    RECT 155.0000 92.8000 155.4000 93.2000 ;
	    RECT 157.4000 93.1000 157.8000 93.2000 ;
	    RECT 162.2000 93.1000 162.6000 93.2000 ;
	    RECT 164.6000 93.1000 165.0000 93.2000 ;
	    RECT 172.6000 93.1000 173.0000 93.2000 ;
	    RECT 179.8000 93.1000 180.2000 93.2000 ;
	    RECT 157.4000 92.8000 180.2000 93.1000 ;
	    RECT 181.4000 93.1000 181.8000 93.2000 ;
	    RECT 186.2000 93.1000 186.6000 93.2000 ;
	    RECT 181.4000 92.8000 186.6000 93.1000 ;
	    RECT 200.6000 92.8000 201.0000 93.2000 ;
	    RECT 201.4000 92.8000 201.8000 93.2000 ;
	    RECT 202.2000 93.1000 202.6000 93.2000 ;
	    RECT 213.4000 93.1000 213.8000 93.2000 ;
	    RECT 202.2000 92.8000 213.8000 93.1000 ;
	    RECT 236.6000 92.8000 237.0000 93.2000 ;
	    RECT 238.2000 93.1000 238.6000 93.2000 ;
	    RECT 241.4000 93.1000 241.8000 93.2000 ;
	    RECT 238.2000 92.8000 241.8000 93.1000 ;
	    RECT 254.2000 93.1000 254.6000 93.2000 ;
	    RECT 255.0000 93.1000 255.4000 93.2000 ;
	    RECT 254.2000 92.8000 255.4000 93.1000 ;
	    RECT 38.2000 92.1000 38.6000 92.2000 ;
	    RECT 42.2000 92.1000 42.6000 92.2000 ;
	    RECT 44.6000 92.1000 45.0000 92.2000 ;
	    RECT 46.2000 92.1000 46.6000 92.2000 ;
	    RECT 54.2000 92.1000 54.6000 92.2000 ;
	    RECT 38.2000 91.8000 54.6000 92.1000 ;
	    RECT 128.6000 92.1000 129.0000 92.2000 ;
	    RECT 131.8000 92.1000 132.2000 92.2000 ;
	    RECT 128.6000 91.8000 132.2000 92.1000 ;
	    RECT 168.6000 92.1000 169.0000 92.2000 ;
	    RECT 169.4000 92.1000 169.8000 92.2000 ;
	    RECT 168.6000 91.8000 169.8000 92.1000 ;
	    RECT 195.0000 92.1000 195.4000 92.2000 ;
	    RECT 201.4000 92.1000 201.7000 92.8000 ;
	    RECT 195.0000 91.8000 201.7000 92.1000 ;
	    RECT 215.0000 92.1000 215.4000 92.2000 ;
	    RECT 218.2000 92.1000 218.6000 92.2000 ;
	    RECT 215.0000 91.8000 218.6000 92.1000 ;
	    RECT 231.0000 92.1000 231.4000 92.2000 ;
	    RECT 236.6000 92.1000 236.9000 92.8000 ;
	    RECT 231.0000 91.8000 236.9000 92.1000 ;
	    RECT 238.2000 92.1000 238.6000 92.2000 ;
	    RECT 259.0000 92.1000 259.4000 92.2000 ;
	    RECT 238.2000 91.8000 259.4000 92.1000 ;
	    RECT 91.8000 91.1000 92.2000 91.2000 ;
	    RECT 105.4000 91.1000 105.8000 91.2000 ;
	    RECT 91.8000 90.8000 105.8000 91.1000 ;
	    RECT 179.8000 91.1000 180.2000 91.2000 ;
	    RECT 183.8000 91.1000 184.2000 91.2000 ;
	    RECT 179.8000 90.8000 184.2000 91.1000 ;
	    RECT 185.4000 91.1000 185.8000 91.2000 ;
	    RECT 188.6000 91.1000 189.0000 91.2000 ;
	    RECT 185.4000 90.8000 189.0000 91.1000 ;
	    RECT 196.6000 91.1000 197.0000 91.2000 ;
	    RECT 209.4000 91.1000 209.8000 91.2000 ;
	    RECT 196.6000 90.8000 209.8000 91.1000 ;
	    RECT 231.8000 91.1000 232.2000 91.2000 ;
	    RECT 237.4000 91.1000 237.8000 91.2000 ;
	    RECT 231.8000 90.8000 237.8000 91.1000 ;
	    RECT 251.0000 91.1000 251.4000 91.2000 ;
	    RECT 265.4000 91.1000 265.8000 91.2000 ;
	    RECT 251.0000 90.8000 265.8000 91.1000 ;
	    RECT 30.2000 89.8000 30.6000 90.2000 ;
	    RECT 57.4000 90.1000 57.8000 90.2000 ;
	    RECT 76.6000 90.1000 77.0000 90.2000 ;
	    RECT 57.4000 89.8000 77.0000 90.1000 ;
	    RECT 86.2000 90.1000 86.6000 90.2000 ;
	    RECT 87.8000 90.1000 88.2000 90.2000 ;
	    RECT 86.2000 89.8000 88.2000 90.1000 ;
	    RECT 88.6000 89.8000 89.0000 90.2000 ;
	    RECT 100.6000 90.1000 101.0000 90.2000 ;
	    RECT 103.0000 90.1000 103.4000 90.2000 ;
	    RECT 100.6000 89.8000 103.4000 90.1000 ;
	    RECT 120.6000 90.1000 121.0000 90.2000 ;
	    RECT 126.2000 90.1000 126.6000 90.2000 ;
	    RECT 120.6000 89.8000 126.6000 90.1000 ;
	    RECT 172.6000 90.1000 173.0000 90.2000 ;
	    RECT 175.8000 90.1000 176.2000 90.2000 ;
	    RECT 172.6000 89.8000 176.2000 90.1000 ;
	    RECT 187.0000 90.1000 187.4000 90.2000 ;
	    RECT 193.4000 90.1000 193.8000 90.2000 ;
	    RECT 200.6000 90.1000 201.0000 90.2000 ;
	    RECT 187.0000 89.8000 201.0000 90.1000 ;
	    RECT 215.0000 90.1000 215.4000 90.2000 ;
	    RECT 229.4000 90.1000 229.8000 90.2000 ;
	    RECT 243.0000 90.1000 243.4000 90.2000 ;
	    RECT 215.0000 89.8000 243.4000 90.1000 ;
	    RECT 259.0000 90.1000 259.4000 90.2000 ;
	    RECT 268.6000 90.1000 269.0000 90.2000 ;
	    RECT 259.0000 89.8000 269.0000 90.1000 ;
	    RECT 30.2000 89.2000 30.5000 89.8000 ;
	    RECT 13.4000 89.1000 13.8000 89.2000 ;
	    RECT 19.0000 89.1000 19.4000 89.2000 ;
	    RECT 13.4000 88.8000 19.4000 89.1000 ;
	    RECT 27.0000 88.8000 27.4000 89.2000 ;
	    RECT 30.2000 88.8000 30.6000 89.2000 ;
	    RECT 47.8000 89.1000 48.2000 89.2000 ;
	    RECT 53.4000 89.1000 53.8000 89.2000 ;
	    RECT 47.8000 88.8000 53.8000 89.1000 ;
	    RECT 57.4000 88.8000 57.8000 89.2000 ;
	    RECT 75.8000 89.1000 76.2000 89.2000 ;
	    RECT 81.4000 89.1000 81.8000 89.2000 ;
	    RECT 75.8000 88.8000 81.8000 89.1000 ;
	    RECT 82.2000 89.1000 82.6000 89.2000 ;
	    RECT 88.6000 89.1000 88.9000 89.8000 ;
	    RECT 82.2000 88.8000 88.9000 89.1000 ;
	    RECT 93.4000 89.1000 93.8000 89.2000 ;
	    RECT 107.8000 89.1000 108.2000 89.2000 ;
	    RECT 114.2000 89.1000 114.6000 89.2000 ;
	    RECT 93.4000 88.8000 114.6000 89.1000 ;
	    RECT 130.2000 88.8000 130.6000 89.2000 ;
	    RECT 146.2000 89.1000 146.6000 89.2000 ;
	    RECT 159.0000 89.1000 159.4000 89.2000 ;
	    RECT 159.8000 89.1000 160.2000 89.2000 ;
	    RECT 146.2000 88.8000 160.2000 89.1000 ;
	    RECT 165.4000 89.1000 165.8000 89.2000 ;
	    RECT 165.4000 88.8000 182.5000 89.1000 ;
	    RECT 27.0000 88.2000 27.3000 88.8000 ;
	    RECT 27.0000 87.8000 27.4000 88.2000 ;
	    RECT 51.8000 88.1000 52.2000 88.2000 ;
	    RECT 57.4000 88.1000 57.7000 88.8000 ;
	    RECT 51.8000 87.8000 57.7000 88.1000 ;
	    RECT 67.8000 88.1000 68.2000 88.2000 ;
	    RECT 71.0000 88.1000 71.4000 88.2000 ;
	    RECT 75.0000 88.1000 75.4000 88.2000 ;
	    RECT 84.6000 88.1000 85.0000 88.2000 ;
	    RECT 96.6000 88.1000 97.0000 88.2000 ;
	    RECT 104.6000 88.1000 105.0000 88.2000 ;
	    RECT 67.8000 87.8000 105.0000 88.1000 ;
	    RECT 127.0000 88.1000 127.4000 88.2000 ;
	    RECT 130.2000 88.1000 130.5000 88.8000 ;
	    RECT 182.2000 88.2000 182.5000 88.8000 ;
	    RECT 183.0000 88.8000 183.4000 89.2000 ;
	    RECT 187.8000 89.1000 188.2000 89.2000 ;
	    RECT 188.6000 89.1000 189.0000 89.2000 ;
	    RECT 187.8000 88.8000 189.0000 89.1000 ;
	    RECT 190.2000 89.1000 190.6000 89.2000 ;
	    RECT 191.0000 89.1000 191.4000 89.2000 ;
	    RECT 226.2000 89.1000 226.6000 89.2000 ;
	    RECT 243.0000 89.1000 243.4000 89.2000 ;
	    RECT 190.2000 88.8000 191.4000 89.1000 ;
	    RECT 198.2000 88.8000 243.4000 89.1000 ;
	    RECT 245.4000 89.1000 245.8000 89.2000 ;
	    RECT 251.0000 89.1000 251.4000 89.2000 ;
	    RECT 251.8000 89.1000 252.2000 89.2000 ;
	    RECT 245.4000 88.8000 252.2000 89.1000 ;
	    RECT 252.6000 89.1000 253.0000 89.2000 ;
	    RECT 260.6000 89.1000 261.0000 89.2000 ;
	    RECT 252.6000 88.8000 261.0000 89.1000 ;
	    RECT 127.0000 87.8000 130.5000 88.1000 ;
	    RECT 145.4000 88.1000 145.8000 88.2000 ;
	    RECT 155.8000 88.1000 156.2000 88.2000 ;
	    RECT 145.4000 87.8000 156.2000 88.1000 ;
	    RECT 159.0000 88.1000 159.4000 88.2000 ;
	    RECT 162.2000 88.1000 162.6000 88.2000 ;
	    RECT 159.0000 87.8000 162.6000 88.1000 ;
	    RECT 164.6000 88.1000 165.0000 88.2000 ;
	    RECT 167.0000 88.1000 167.4000 88.2000 ;
	    RECT 164.6000 87.8000 167.4000 88.1000 ;
	    RECT 171.8000 88.1000 172.2000 88.2000 ;
	    RECT 181.4000 88.1000 181.8000 88.2000 ;
	    RECT 171.8000 87.8000 181.8000 88.1000 ;
	    RECT 182.2000 87.8000 182.6000 88.2000 ;
	    RECT 183.0000 88.1000 183.3000 88.8000 ;
	    RECT 198.2000 88.2000 198.5000 88.8000 ;
	    RECT 195.8000 88.1000 196.2000 88.2000 ;
	    RECT 197.4000 88.1000 197.8000 88.2000 ;
	    RECT 183.0000 87.8000 197.8000 88.1000 ;
	    RECT 198.2000 87.8000 198.6000 88.2000 ;
	    RECT 199.0000 88.1000 199.4000 88.2000 ;
	    RECT 206.2000 88.1000 206.6000 88.2000 ;
	    RECT 215.0000 88.1000 215.4000 88.2000 ;
	    RECT 199.0000 87.8000 215.4000 88.1000 ;
	    RECT 219.8000 88.1000 220.2000 88.2000 ;
	    RECT 225.4000 88.1000 225.8000 88.2000 ;
	    RECT 227.0000 88.1000 227.4000 88.2000 ;
	    RECT 219.8000 87.8000 224.9000 88.1000 ;
	    RECT 225.4000 87.8000 227.4000 88.1000 ;
	    RECT 231.8000 87.8000 232.2000 88.2000 ;
	    RECT 224.6000 87.2000 224.9000 87.8000 ;
	    RECT 44.6000 86.8000 45.0000 87.2000 ;
	    RECT 49.4000 87.1000 49.8000 87.2000 ;
	    RECT 55.8000 87.1000 56.2000 87.2000 ;
	    RECT 57.4000 87.1000 57.8000 87.2000 ;
	    RECT 49.4000 86.8000 57.8000 87.1000 ;
	    RECT 73.4000 86.8000 73.8000 87.2000 ;
	    RECT 90.2000 87.1000 90.6000 87.2000 ;
	    RECT 99.0000 87.1000 99.4000 87.2000 ;
	    RECT 90.2000 86.8000 99.4000 87.1000 ;
	    RECT 102.2000 87.1000 102.6000 87.2000 ;
	    RECT 108.6000 87.1000 109.0000 87.2000 ;
	    RECT 102.2000 86.8000 109.0000 87.1000 ;
	    RECT 112.6000 86.8000 113.0000 87.2000 ;
	    RECT 127.0000 86.8000 127.4000 87.2000 ;
	    RECT 152.6000 86.8000 153.0000 87.2000 ;
	    RECT 161.4000 87.1000 161.8000 87.2000 ;
	    RECT 164.6000 87.1000 165.0000 87.2000 ;
	    RECT 161.4000 86.8000 165.0000 87.1000 ;
	    RECT 170.2000 87.1000 170.6000 87.2000 ;
	    RECT 184.6000 87.1000 185.0000 87.2000 ;
	    RECT 170.2000 86.8000 185.0000 87.1000 ;
	    RECT 185.4000 87.1000 185.8000 87.2000 ;
	    RECT 191.8000 87.1000 192.2000 87.2000 ;
	    RECT 185.4000 86.8000 192.2000 87.1000 ;
	    RECT 194.2000 87.1000 194.6000 87.2000 ;
	    RECT 202.2000 87.1000 202.6000 87.2000 ;
	    RECT 194.2000 86.8000 202.6000 87.1000 ;
	    RECT 206.2000 87.1000 206.6000 87.2000 ;
	    RECT 207.0000 87.1000 207.4000 87.2000 ;
	    RECT 206.2000 86.8000 207.4000 87.1000 ;
	    RECT 221.4000 87.1000 221.8000 87.2000 ;
	    RECT 223.0000 87.1000 223.4000 87.2000 ;
	    RECT 221.4000 86.8000 223.4000 87.1000 ;
	    RECT 224.6000 86.8000 225.0000 87.2000 ;
	    RECT 225.4000 87.1000 225.8000 87.2000 ;
	    RECT 227.8000 87.1000 228.2000 87.2000 ;
	    RECT 225.4000 86.8000 228.2000 87.1000 ;
	    RECT 231.8000 87.1000 232.1000 87.8000 ;
	    RECT 233.4000 87.1000 233.8000 87.2000 ;
	    RECT 231.8000 86.8000 233.8000 87.1000 ;
	    RECT 255.0000 87.1000 255.4000 87.2000 ;
	    RECT 255.8000 87.1000 256.2000 87.2000 ;
	    RECT 255.0000 86.8000 256.2000 87.1000 ;
	    RECT 44.6000 86.1000 44.9000 86.8000 ;
	    RECT 59.8000 86.1000 60.2000 86.2000 ;
	    RECT 44.6000 85.8000 60.2000 86.1000 ;
	    RECT 73.4000 86.1000 73.7000 86.8000 ;
	    RECT 76.6000 86.1000 77.0000 86.2000 ;
	    RECT 102.2000 86.1000 102.6000 86.2000 ;
	    RECT 111.8000 86.1000 112.2000 86.2000 ;
	    RECT 73.4000 85.8000 77.0000 86.1000 ;
	    RECT 101.4000 85.8000 112.2000 86.1000 ;
	    RECT 112.6000 86.1000 112.9000 86.8000 ;
	    RECT 115.0000 86.1000 115.4000 86.2000 ;
	    RECT 112.6000 85.8000 115.4000 86.1000 ;
	    RECT 127.0000 86.1000 127.3000 86.8000 ;
	    RECT 130.2000 86.1000 130.6000 86.2000 ;
	    RECT 127.0000 85.8000 130.6000 86.1000 ;
	    RECT 152.6000 86.1000 152.9000 86.8000 ;
	    RECT 170.2000 86.2000 170.5000 86.8000 ;
	    RECT 160.6000 86.1000 161.0000 86.2000 ;
	    RECT 152.6000 85.8000 161.0000 86.1000 ;
	    RECT 170.2000 85.8000 170.6000 86.2000 ;
	    RECT 181.4000 86.1000 181.8000 86.2000 ;
	    RECT 195.0000 86.1000 195.4000 86.2000 ;
	    RECT 195.8000 86.1000 196.2000 86.2000 ;
	    RECT 181.4000 85.8000 196.2000 86.1000 ;
	    RECT 207.8000 86.1000 208.2000 86.2000 ;
	    RECT 212.6000 86.1000 213.0000 86.2000 ;
	    RECT 207.8000 85.8000 213.0000 86.1000 ;
	    RECT 218.2000 86.1000 218.6000 86.2000 ;
	    RECT 222.2000 86.1000 222.6000 86.2000 ;
	    RECT 218.2000 85.8000 222.6000 86.1000 ;
	    RECT 223.8000 86.1000 224.2000 86.2000 ;
	    RECT 234.2000 86.1000 234.6000 86.2000 ;
	    RECT 223.8000 85.8000 234.6000 86.1000 ;
	    RECT 239.0000 86.1000 239.4000 86.2000 ;
	    RECT 244.6000 86.1000 245.0000 86.2000 ;
	    RECT 239.0000 85.8000 245.0000 86.1000 ;
	    RECT 253.4000 86.1000 253.8000 86.2000 ;
	    RECT 256.6000 86.1000 257.0000 86.2000 ;
	    RECT 253.4000 85.8000 257.0000 86.1000 ;
	    RECT 1.4000 85.1000 1.8000 85.2000 ;
	    RECT 4.6000 85.1000 5.0000 85.2000 ;
	    RECT 1.4000 84.8000 5.0000 85.1000 ;
	    RECT 54.2000 85.1000 54.6000 85.2000 ;
	    RECT 58.2000 85.1000 58.6000 85.2000 ;
	    RECT 54.2000 84.8000 58.6000 85.1000 ;
	    RECT 63.0000 85.1000 63.4000 85.2000 ;
	    RECT 75.0000 85.1000 75.4000 85.2000 ;
	    RECT 63.0000 84.8000 75.4000 85.1000 ;
	    RECT 100.6000 85.1000 101.0000 85.2000 ;
	    RECT 116.6000 85.1000 117.0000 85.2000 ;
	    RECT 123.8000 85.1000 124.2000 85.2000 ;
	    RECT 100.6000 84.8000 124.2000 85.1000 ;
	    RECT 159.0000 85.1000 159.4000 85.2000 ;
	    RECT 179.8000 85.1000 180.2000 85.2000 ;
	    RECT 159.0000 84.8000 180.2000 85.1000 ;
	    RECT 184.6000 85.1000 185.0000 85.2000 ;
	    RECT 195.8000 85.1000 196.2000 85.2000 ;
	    RECT 184.6000 84.8000 196.2000 85.1000 ;
	    RECT 199.8000 84.8000 204.9000 85.1000 ;
	    RECT 199.8000 84.2000 200.1000 84.8000 ;
	    RECT 204.6000 84.2000 204.9000 84.8000 ;
	    RECT 205.4000 84.8000 205.8000 85.2000 ;
	    RECT 207.8000 85.1000 208.2000 85.2000 ;
	    RECT 208.6000 85.1000 209.0000 85.2000 ;
	    RECT 207.8000 84.8000 209.0000 85.1000 ;
	    RECT 219.8000 85.1000 220.2000 85.2000 ;
	    RECT 231.8000 85.1000 232.2000 85.2000 ;
	    RECT 251.8000 85.1000 252.2000 85.2000 ;
	    RECT 219.8000 84.8000 232.2000 85.1000 ;
	    RECT 245.4000 84.8000 252.2000 85.1000 ;
	    RECT 256.6000 85.1000 257.0000 85.2000 ;
	    RECT 257.4000 85.1000 257.8000 85.2000 ;
	    RECT 256.6000 84.8000 257.8000 85.1000 ;
	    RECT 205.4000 84.2000 205.7000 84.8000 ;
	    RECT 245.4000 84.2000 245.7000 84.8000 ;
	    RECT 49.4000 84.1000 49.8000 84.2000 ;
	    RECT 50.2000 84.1000 50.6000 84.2000 ;
	    RECT 49.4000 83.8000 50.6000 84.1000 ;
	    RECT 65.4000 84.1000 65.8000 84.2000 ;
	    RECT 72.6000 84.1000 73.0000 84.2000 ;
	    RECT 65.4000 83.8000 73.0000 84.1000 ;
	    RECT 141.4000 84.1000 141.8000 84.2000 ;
	    RECT 152.6000 84.1000 153.0000 84.2000 ;
	    RECT 141.4000 83.8000 153.0000 84.1000 ;
	    RECT 178.2000 84.1000 178.6000 84.2000 ;
	    RECT 194.2000 84.1000 194.6000 84.2000 ;
	    RECT 178.2000 83.8000 194.6000 84.1000 ;
	    RECT 195.8000 84.1000 196.2000 84.2000 ;
	    RECT 199.0000 84.1000 199.4000 84.2000 ;
	    RECT 195.8000 83.8000 199.4000 84.1000 ;
	    RECT 199.8000 83.8000 200.2000 84.2000 ;
	    RECT 204.6000 83.8000 205.0000 84.2000 ;
	    RECT 205.4000 83.8000 205.8000 84.2000 ;
	    RECT 234.2000 84.1000 234.6000 84.2000 ;
	    RECT 235.0000 84.1000 235.4000 84.2000 ;
	    RECT 234.2000 83.8000 235.4000 84.1000 ;
	    RECT 245.4000 83.8000 245.8000 84.2000 ;
	    RECT 65.4000 83.2000 65.7000 83.8000 ;
	    RECT 47.8000 83.1000 48.2000 83.2000 ;
	    RECT 56.6000 83.1000 57.0000 83.2000 ;
	    RECT 47.8000 82.8000 57.0000 83.1000 ;
	    RECT 65.4000 82.8000 65.8000 83.2000 ;
	    RECT 115.0000 83.1000 115.4000 83.2000 ;
	    RECT 117.4000 83.1000 117.8000 83.2000 ;
	    RECT 137.4000 83.1000 137.8000 83.2000 ;
	    RECT 115.0000 82.8000 137.8000 83.1000 ;
	    RECT 203.8000 83.1000 204.2000 83.2000 ;
	    RECT 219.8000 83.1000 220.2000 83.2000 ;
	    RECT 203.8000 82.8000 220.2000 83.1000 ;
	    RECT 254.2000 83.1000 254.6000 83.2000 ;
	    RECT 262.2000 83.1000 262.6000 83.2000 ;
	    RECT 254.2000 82.8000 262.6000 83.1000 ;
	    RECT 62.2000 82.1000 62.6000 82.2000 ;
	    RECT 74.2000 82.1000 74.6000 82.2000 ;
	    RECT 62.2000 81.8000 74.6000 82.1000 ;
	    RECT 131.8000 82.1000 132.2000 82.2000 ;
	    RECT 135.8000 82.1000 136.2000 82.2000 ;
	    RECT 140.6000 82.1000 141.0000 82.2000 ;
	    RECT 131.8000 81.8000 141.0000 82.1000 ;
	    RECT 195.0000 82.1000 195.4000 82.2000 ;
	    RECT 218.2000 82.1000 218.6000 82.2000 ;
	    RECT 195.0000 81.8000 218.6000 82.1000 ;
	    RECT 188.6000 81.1000 189.0000 81.2000 ;
	    RECT 199.0000 81.1000 199.4000 81.2000 ;
	    RECT 208.6000 81.1000 209.0000 81.2000 ;
	    RECT 188.6000 80.8000 209.0000 81.1000 ;
	    RECT 98.2000 80.1000 98.6000 80.2000 ;
	    RECT 101.4000 80.1000 101.8000 80.2000 ;
	    RECT 98.2000 79.8000 101.8000 80.1000 ;
	    RECT 179.8000 80.1000 180.2000 80.2000 ;
	    RECT 204.6000 80.1000 205.0000 80.2000 ;
	    RECT 179.8000 79.8000 205.0000 80.1000 ;
	    RECT 248.6000 80.1000 249.0000 80.2000 ;
	    RECT 256.6000 80.1000 257.0000 80.2000 ;
	    RECT 248.6000 79.8000 257.0000 80.1000 ;
	    RECT 46.2000 79.1000 46.6000 79.2000 ;
	    RECT 52.6000 79.1000 53.0000 79.2000 ;
	    RECT 46.2000 78.8000 53.0000 79.1000 ;
	    RECT 55.8000 79.1000 56.2000 79.2000 ;
	    RECT 57.4000 79.1000 57.8000 79.2000 ;
	    RECT 55.8000 78.8000 57.8000 79.1000 ;
	    RECT 242.2000 79.1000 242.6000 79.2000 ;
	    RECT 252.6000 79.1000 253.0000 79.2000 ;
	    RECT 242.2000 78.8000 253.0000 79.1000 ;
	    RECT 268.6000 78.8000 269.0000 79.2000 ;
	    RECT 7.8000 78.1000 8.2000 78.2000 ;
	    RECT 8.6000 78.1000 9.0000 78.2000 ;
	    RECT 7.8000 77.8000 9.0000 78.1000 ;
	    RECT 10.2000 77.8000 10.6000 78.2000 ;
	    RECT 17.4000 78.1000 17.8000 78.2000 ;
	    RECT 18.2000 78.1000 18.6000 78.2000 ;
	    RECT 17.4000 77.8000 18.6000 78.1000 ;
	    RECT 30.2000 77.8000 30.6000 78.2000 ;
	    RECT 244.6000 78.1000 245.0000 78.2000 ;
	    RECT 257.4000 78.1000 257.8000 78.2000 ;
	    RECT 244.6000 77.8000 257.8000 78.1000 ;
	    RECT 259.8000 78.1000 260.2000 78.2000 ;
	    RECT 268.6000 78.1000 268.9000 78.8000 ;
	    RECT 259.8000 77.8000 268.9000 78.1000 ;
	    RECT 5.4000 77.1000 5.8000 77.2000 ;
	    RECT 10.2000 77.1000 10.5000 77.8000 ;
	    RECT 30.2000 77.2000 30.5000 77.8000 ;
	    RECT 5.4000 76.8000 10.5000 77.1000 ;
	    RECT 12.6000 77.1000 13.0000 77.2000 ;
	    RECT 17.4000 77.1000 17.8000 77.2000 ;
	    RECT 12.6000 76.8000 17.8000 77.1000 ;
	    RECT 27.0000 76.8000 27.4000 77.2000 ;
	    RECT 30.2000 76.8000 30.6000 77.2000 ;
	    RECT 31.0000 76.8000 31.4000 77.2000 ;
	    RECT 44.6000 76.8000 45.0000 77.2000 ;
	    RECT 55.8000 77.1000 56.2000 77.2000 ;
	    RECT 60.6000 77.1000 61.0000 77.2000 ;
	    RECT 72.6000 77.1000 73.0000 77.2000 ;
	    RECT 55.8000 76.8000 73.0000 77.1000 ;
	    RECT 75.8000 77.1000 76.2000 77.2000 ;
	    RECT 79.8000 77.1000 80.2000 77.2000 ;
	    RECT 95.0000 77.1000 95.4000 77.2000 ;
	    RECT 75.8000 76.8000 95.4000 77.1000 ;
	    RECT 181.4000 77.1000 181.8000 77.2000 ;
	    RECT 183.0000 77.1000 183.4000 77.2000 ;
	    RECT 181.4000 76.8000 183.4000 77.1000 ;
	    RECT 185.4000 77.1000 185.8000 77.2000 ;
	    RECT 191.0000 77.1000 191.4000 77.2000 ;
	    RECT 185.4000 76.8000 191.4000 77.1000 ;
	    RECT 194.2000 76.8000 194.6000 77.2000 ;
	    RECT 201.4000 76.8000 201.8000 77.2000 ;
	    RECT 205.4000 77.1000 205.8000 77.2000 ;
	    RECT 222.2000 77.1000 222.6000 77.2000 ;
	    RECT 205.4000 76.8000 222.6000 77.1000 ;
	    RECT 223.8000 77.1000 224.2000 77.2000 ;
	    RECT 229.4000 77.1000 229.8000 77.2000 ;
	    RECT 223.8000 76.8000 229.8000 77.1000 ;
	    RECT 247.8000 77.1000 248.2000 77.2000 ;
	    RECT 256.6000 77.1000 257.0000 77.2000 ;
	    RECT 260.6000 77.1000 261.0000 77.2000 ;
	    RECT 247.8000 76.8000 261.0000 77.1000 ;
	    RECT 16.6000 76.1000 17.0000 76.2000 ;
	    RECT 20.6000 76.1000 21.0000 76.2000 ;
	    RECT 16.6000 75.8000 21.0000 76.1000 ;
	    RECT 23.0000 76.1000 23.4000 76.2000 ;
	    RECT 23.8000 76.1000 24.2000 76.2000 ;
	    RECT 25.4000 76.1000 25.8000 76.2000 ;
	    RECT 23.0000 75.8000 25.8000 76.1000 ;
	    RECT 27.0000 76.1000 27.3000 76.8000 ;
	    RECT 31.0000 76.1000 31.3000 76.8000 ;
	    RECT 27.0000 75.8000 31.3000 76.1000 ;
	    RECT 44.6000 76.1000 44.9000 76.8000 ;
	    RECT 51.0000 76.1000 51.4000 76.2000 ;
	    RECT 44.6000 75.8000 51.4000 76.1000 ;
	    RECT 65.4000 76.1000 65.8000 76.2000 ;
	    RECT 71.8000 76.1000 72.2000 76.2000 ;
	    RECT 65.4000 75.8000 72.2000 76.1000 ;
	    RECT 108.6000 75.8000 109.0000 76.2000 ;
	    RECT 159.0000 76.1000 159.4000 76.2000 ;
	    RECT 161.4000 76.1000 161.8000 76.2000 ;
	    RECT 159.0000 75.8000 161.8000 76.1000 ;
	    RECT 167.0000 76.1000 167.4000 76.2000 ;
	    RECT 185.4000 76.1000 185.7000 76.8000 ;
	    RECT 167.0000 75.8000 185.7000 76.1000 ;
	    RECT 194.2000 76.2000 194.5000 76.8000 ;
	    RECT 194.2000 75.8000 194.6000 76.2000 ;
	    RECT 201.4000 76.1000 201.7000 76.8000 ;
	    RECT 207.8000 76.1000 208.2000 76.2000 ;
	    RECT 201.4000 75.8000 208.2000 76.1000 ;
	    RECT 209.4000 76.1000 209.8000 76.2000 ;
	    RECT 228.6000 76.1000 229.0000 76.2000 ;
	    RECT 238.2000 76.1000 238.6000 76.2000 ;
	    RECT 240.6000 76.1000 241.0000 76.2000 ;
	    RECT 243.8000 76.1000 244.2000 76.2000 ;
	    RECT 255.0000 76.1000 255.4000 76.2000 ;
	    RECT 209.4000 75.8000 255.4000 76.1000 ;
	    RECT 259.0000 75.8000 259.4000 76.2000 ;
	    RECT 265.4000 76.1000 265.8000 76.2000 ;
	    RECT 267.0000 76.1000 267.4000 76.2000 ;
	    RECT 265.4000 75.8000 267.4000 76.1000 ;
	    RECT 4.6000 75.1000 5.0000 75.2000 ;
	    RECT 5.4000 75.1000 5.8000 75.2000 ;
	    RECT 3.8000 74.8000 5.8000 75.1000 ;
	    RECT 6.2000 74.8000 6.6000 75.2000 ;
	    RECT 9.4000 75.1000 9.8000 75.2000 ;
	    RECT 10.2000 75.1000 10.6000 75.2000 ;
	    RECT 9.4000 74.8000 10.6000 75.1000 ;
	    RECT 27.0000 74.8000 27.4000 75.2000 ;
	    RECT 27.8000 75.1000 28.2000 75.2000 ;
	    RECT 28.6000 75.1000 29.0000 75.2000 ;
	    RECT 27.8000 74.8000 29.0000 75.1000 ;
	    RECT 45.4000 75.1000 45.8000 75.2000 ;
	    RECT 47.0000 75.1000 47.4000 75.2000 ;
	    RECT 45.4000 74.8000 47.4000 75.1000 ;
	    RECT 49.4000 74.8000 49.8000 75.2000 ;
	    RECT 69.4000 75.1000 69.8000 75.2000 ;
	    RECT 65.4000 74.8000 69.8000 75.1000 ;
	    RECT 72.6000 75.1000 73.0000 75.2000 ;
	    RECT 76.6000 75.1000 77.0000 75.2000 ;
	    RECT 72.6000 74.8000 77.0000 75.1000 ;
	    RECT 78.2000 75.1000 78.6000 75.2000 ;
	    RECT 89.4000 75.1000 89.8000 75.2000 ;
	    RECT 95.0000 75.1000 95.4000 75.2000 ;
	    RECT 78.2000 74.8000 95.4000 75.1000 ;
	    RECT 97.4000 75.1000 97.8000 75.2000 ;
	    RECT 108.6000 75.1000 108.9000 75.8000 ;
	    RECT 259.0000 75.2000 259.3000 75.8000 ;
	    RECT 97.4000 74.8000 108.9000 75.1000 ;
	    RECT 111.0000 75.1000 111.4000 75.2000 ;
	    RECT 118.2000 75.1000 118.6000 75.2000 ;
	    RECT 111.0000 74.8000 118.6000 75.1000 ;
	    RECT 119.8000 75.1000 120.2000 75.2000 ;
	    RECT 136.6000 75.1000 137.0000 75.2000 ;
	    RECT 119.8000 74.8000 121.7000 75.1000 ;
	    RECT 2.2000 74.1000 2.6000 74.2000 ;
	    RECT 6.2000 74.1000 6.5000 74.8000 ;
	    RECT 27.0000 74.2000 27.3000 74.8000 ;
	    RECT 49.4000 74.2000 49.7000 74.8000 ;
	    RECT 65.4000 74.7000 65.8000 74.8000 ;
	    RECT 121.4000 74.2000 121.7000 74.8000 ;
	    RECT 124.6000 74.8000 137.0000 75.1000 ;
	    RECT 144.6000 74.8000 145.0000 75.2000 ;
	    RECT 155.8000 75.1000 156.2000 75.2000 ;
	    RECT 160.6000 75.1000 161.0000 75.2000 ;
	    RECT 162.2000 75.1000 162.6000 75.2000 ;
	    RECT 163.8000 75.1000 164.2000 75.2000 ;
	    RECT 155.8000 74.8000 164.2000 75.1000 ;
	    RECT 168.6000 75.1000 169.0000 75.2000 ;
	    RECT 181.4000 75.1000 181.8000 75.2000 ;
	    RECT 168.6000 74.8000 181.8000 75.1000 ;
	    RECT 184.6000 75.1000 185.0000 75.2000 ;
	    RECT 191.8000 75.1000 192.2000 75.2000 ;
	    RECT 184.6000 74.8000 192.2000 75.1000 ;
	    RECT 193.4000 74.8000 193.8000 75.2000 ;
	    RECT 195.8000 75.1000 196.2000 75.2000 ;
	    RECT 199.8000 75.1000 200.2000 75.2000 ;
	    RECT 195.8000 74.8000 200.2000 75.1000 ;
	    RECT 205.4000 75.1000 205.8000 75.2000 ;
	    RECT 226.2000 75.1000 226.6000 75.2000 ;
	    RECT 229.4000 75.1000 229.8000 75.2000 ;
	    RECT 205.4000 74.8000 213.8000 75.1000 ;
	    RECT 226.2000 74.8000 229.8000 75.1000 ;
	    RECT 232.6000 75.1000 233.0000 75.2000 ;
	    RECT 234.2000 75.1000 234.6000 75.2000 ;
	    RECT 232.6000 74.8000 234.6000 75.1000 ;
	    RECT 236.6000 75.1000 237.0000 75.2000 ;
	    RECT 239.0000 75.1000 239.4000 75.2000 ;
	    RECT 236.6000 74.8000 240.1000 75.1000 ;
	    RECT 259.0000 74.8000 259.4000 75.2000 ;
	    RECT 124.6000 74.2000 124.9000 74.8000 ;
	    RECT 2.2000 73.8000 6.5000 74.1000 ;
	    RECT 17.4000 74.1000 17.8000 74.2000 ;
	    RECT 24.6000 74.1000 25.0000 74.2000 ;
	    RECT 17.4000 73.8000 25.0000 74.1000 ;
	    RECT 27.0000 73.8000 27.4000 74.2000 ;
	    RECT 42.2000 74.1000 42.6000 74.2000 ;
	    RECT 44.6000 74.1000 45.0000 74.2000 ;
	    RECT 42.2000 73.8000 45.0000 74.1000 ;
	    RECT 49.4000 73.8000 49.8000 74.2000 ;
	    RECT 54.2000 74.1000 54.6000 74.2000 ;
	    RECT 70.2000 74.1000 70.6000 74.2000 ;
	    RECT 54.2000 73.8000 70.6000 74.1000 ;
	    RECT 71.8000 74.1000 72.2000 74.2000 ;
	    RECT 90.2000 74.1000 90.6000 74.2000 ;
	    RECT 91.8000 74.1000 92.2000 74.2000 ;
	    RECT 71.8000 73.8000 92.2000 74.1000 ;
	    RECT 95.0000 74.1000 95.4000 74.2000 ;
	    RECT 100.6000 74.1000 101.0000 74.2000 ;
	    RECT 95.0000 73.8000 101.0000 74.1000 ;
	    RECT 102.2000 73.8000 102.6000 74.2000 ;
	    RECT 103.8000 73.8000 104.2000 74.2000 ;
	    RECT 121.4000 73.8000 121.8000 74.2000 ;
	    RECT 124.6000 73.8000 125.0000 74.2000 ;
	    RECT 136.6000 74.1000 136.9000 74.8000 ;
	    RECT 144.6000 74.1000 144.9000 74.8000 ;
	    RECT 136.6000 73.8000 144.9000 74.1000 ;
	    RECT 164.6000 74.1000 165.0000 74.2000 ;
	    RECT 173.4000 74.1000 173.8000 74.2000 ;
	    RECT 164.6000 73.8000 173.8000 74.1000 ;
	    RECT 178.2000 73.8000 178.6000 74.2000 ;
	    RECT 184.6000 74.1000 185.0000 74.2000 ;
	    RECT 186.2000 74.1000 186.6000 74.2000 ;
	    RECT 184.6000 73.8000 186.6000 74.1000 ;
	    RECT 188.6000 74.1000 189.0000 74.2000 ;
	    RECT 189.4000 74.1000 189.8000 74.2000 ;
	    RECT 188.6000 73.8000 189.8000 74.1000 ;
	    RECT 193.4000 74.1000 193.7000 74.8000 ;
	    RECT 213.4000 74.7000 213.8000 74.8000 ;
	    RECT 195.8000 74.1000 196.2000 74.2000 ;
	    RECT 193.4000 73.8000 196.2000 74.1000 ;
	    RECT 202.2000 74.1000 202.6000 74.2000 ;
	    RECT 206.2000 74.1000 206.6000 74.2000 ;
	    RECT 202.2000 73.8000 206.6000 74.1000 ;
	    RECT 207.0000 74.1000 207.4000 74.2000 ;
	    RECT 207.8000 74.1000 208.2000 74.2000 ;
	    RECT 207.0000 73.8000 208.2000 74.1000 ;
	    RECT 209.4000 74.1000 209.8000 74.2000 ;
	    RECT 217.4000 74.1000 217.8000 74.2000 ;
	    RECT 223.0000 74.1000 223.4000 74.2000 ;
	    RECT 209.4000 73.8000 211.3000 74.1000 ;
	    RECT 217.4000 73.8000 223.4000 74.1000 ;
	    RECT 227.0000 74.1000 227.4000 74.2000 ;
	    RECT 230.2000 74.1000 230.6000 74.2000 ;
	    RECT 227.0000 73.8000 230.6000 74.1000 ;
	    RECT 237.4000 74.1000 237.8000 74.2000 ;
	    RECT 239.8000 74.1000 240.2000 74.2000 ;
	    RECT 240.6000 74.1000 241.0000 74.2000 ;
	    RECT 237.4000 73.8000 241.0000 74.1000 ;
	    RECT 102.2000 73.2000 102.5000 73.8000 ;
	    RECT 103.8000 73.2000 104.1000 73.8000 ;
	    RECT 14.2000 73.1000 14.6000 73.2000 ;
	    RECT 22.2000 73.1000 22.6000 73.2000 ;
	    RECT 24.6000 73.1000 25.0000 73.2000 ;
	    RECT 14.2000 72.8000 25.0000 73.1000 ;
	    RECT 26.2000 73.1000 26.6000 73.2000 ;
	    RECT 27.8000 73.1000 28.2000 73.2000 ;
	    RECT 26.2000 72.8000 28.2000 73.1000 ;
	    RECT 46.2000 73.1000 46.6000 73.2000 ;
	    RECT 47.8000 73.1000 48.2000 73.2000 ;
	    RECT 46.2000 72.8000 48.2000 73.1000 ;
	    RECT 59.8000 73.1000 60.2000 73.2000 ;
	    RECT 69.4000 73.1000 69.8000 73.2000 ;
	    RECT 59.8000 72.8000 69.8000 73.1000 ;
	    RECT 74.2000 73.1000 74.6000 73.2000 ;
	    RECT 83.8000 73.1000 84.2000 73.2000 ;
	    RECT 74.2000 72.8000 84.2000 73.1000 ;
	    RECT 95.8000 73.1000 96.2000 73.2000 ;
	    RECT 96.6000 73.1000 97.0000 73.2000 ;
	    RECT 95.8000 72.8000 97.0000 73.1000 ;
	    RECT 102.2000 72.8000 102.6000 73.2000 ;
	    RECT 103.8000 72.8000 104.2000 73.2000 ;
	    RECT 104.6000 73.1000 105.0000 73.2000 ;
	    RECT 143.8000 73.1000 144.2000 73.2000 ;
	    RECT 166.2000 73.1000 166.6000 73.2000 ;
	    RECT 104.6000 72.8000 166.6000 73.1000 ;
	    RECT 171.0000 73.1000 171.4000 73.2000 ;
	    RECT 178.2000 73.1000 178.5000 73.8000 ;
	    RECT 211.0000 73.2000 211.3000 73.8000 ;
	    RECT 171.0000 72.8000 178.5000 73.1000 ;
	    RECT 179.0000 73.1000 179.4000 73.2000 ;
	    RECT 179.8000 73.1000 180.2000 73.2000 ;
	    RECT 179.0000 72.8000 180.2000 73.1000 ;
	    RECT 187.0000 72.8000 187.4000 73.2000 ;
	    RECT 203.0000 73.1000 203.4000 73.2000 ;
	    RECT 204.6000 73.1000 205.0000 73.2000 ;
	    RECT 203.0000 72.8000 205.0000 73.1000 ;
	    RECT 211.0000 72.8000 211.4000 73.2000 ;
	    RECT 215.8000 73.1000 216.2000 73.2000 ;
	    RECT 227.8000 73.1000 228.2000 73.2000 ;
	    RECT 243.0000 73.1000 243.4000 73.2000 ;
	    RECT 215.8000 72.8000 243.4000 73.1000 ;
	    RECT 255.8000 73.1000 256.2000 73.2000 ;
	    RECT 259.0000 73.1000 259.4000 73.2000 ;
	    RECT 255.8000 72.8000 259.4000 73.1000 ;
	    RECT 263.0000 73.1000 263.4000 73.2000 ;
	    RECT 263.8000 73.1000 264.2000 73.2000 ;
	    RECT 263.0000 72.8000 264.2000 73.1000 ;
	    RECT 13.4000 72.1000 13.8000 72.2000 ;
	    RECT 14.2000 72.1000 14.6000 72.2000 ;
	    RECT 13.4000 71.8000 14.6000 72.1000 ;
	    RECT 17.4000 71.8000 17.8000 72.2000 ;
	    RECT 22.2000 72.1000 22.6000 72.2000 ;
	    RECT 23.0000 72.1000 23.4000 72.2000 ;
	    RECT 22.2000 71.8000 23.4000 72.1000 ;
	    RECT 23.8000 72.1000 24.2000 72.2000 ;
	    RECT 31.8000 72.1000 32.2000 72.2000 ;
	    RECT 23.8000 71.8000 32.2000 72.1000 ;
	    RECT 33.4000 72.1000 33.8000 72.2000 ;
	    RECT 38.2000 72.1000 38.6000 72.2000 ;
	    RECT 33.4000 71.8000 38.6000 72.1000 ;
	    RECT 49.4000 72.1000 49.8000 72.2000 ;
	    RECT 51.8000 72.1000 52.2000 72.2000 ;
	    RECT 49.4000 71.8000 52.2000 72.1000 ;
	    RECT 70.2000 72.1000 70.6000 72.2000 ;
	    RECT 75.8000 72.1000 76.2000 72.2000 ;
	    RECT 70.2000 71.8000 76.2000 72.1000 ;
	    RECT 79.0000 71.8000 79.4000 72.2000 ;
	    RECT 88.6000 72.1000 89.0000 72.2000 ;
	    RECT 94.2000 72.1000 94.6000 72.2000 ;
	    RECT 107.0000 72.1000 107.4000 72.2000 ;
	    RECT 115.8000 72.1000 116.2000 72.2000 ;
	    RECT 88.6000 71.8000 116.2000 72.1000 ;
	    RECT 129.4000 72.1000 129.8000 72.2000 ;
	    RECT 139.0000 72.1000 139.4000 72.2000 ;
	    RECT 129.4000 71.8000 139.4000 72.1000 ;
	    RECT 175.0000 72.1000 175.4000 72.2000 ;
	    RECT 175.8000 72.1000 176.2000 72.2000 ;
	    RECT 175.0000 71.8000 176.2000 72.1000 ;
	    RECT 177.4000 72.1000 177.8000 72.2000 ;
	    RECT 187.0000 72.1000 187.3000 72.8000 ;
	    RECT 177.4000 71.8000 187.3000 72.1000 ;
	    RECT 202.2000 72.1000 202.6000 72.2000 ;
	    RECT 209.4000 72.1000 209.8000 72.2000 ;
	    RECT 202.2000 71.8000 209.8000 72.1000 ;
	    RECT 219.8000 72.1000 220.2000 72.2000 ;
	    RECT 220.6000 72.1000 221.0000 72.2000 ;
	    RECT 219.8000 71.8000 221.0000 72.1000 ;
	    RECT 221.4000 72.1000 221.8000 72.2000 ;
	    RECT 229.4000 72.1000 229.8000 72.2000 ;
	    RECT 221.4000 71.8000 229.8000 72.1000 ;
	    RECT 230.2000 72.1000 230.6000 72.2000 ;
	    RECT 239.0000 72.1000 239.4000 72.2000 ;
	    RECT 230.2000 71.8000 239.4000 72.1000 ;
	    RECT 240.6000 72.1000 241.0000 72.2000 ;
	    RECT 243.0000 72.1000 243.4000 72.2000 ;
	    RECT 240.6000 71.8000 243.4000 72.1000 ;
	    RECT 243.8000 72.1000 244.2000 72.2000 ;
	    RECT 248.6000 72.1000 249.0000 72.2000 ;
	    RECT 243.8000 71.8000 249.0000 72.1000 ;
	    RECT 267.0000 72.1000 267.4000 72.2000 ;
	    RECT 268.6000 72.1000 269.0000 72.2000 ;
	    RECT 267.0000 71.8000 269.0000 72.1000 ;
	    RECT 17.4000 71.2000 17.7000 71.8000 ;
	    RECT 79.0000 71.2000 79.3000 71.8000 ;
	    RECT 17.4000 70.8000 17.8000 71.2000 ;
	    RECT 22.2000 71.1000 22.6000 71.2000 ;
	    RECT 23.0000 71.1000 23.4000 71.2000 ;
	    RECT 22.2000 70.8000 23.4000 71.1000 ;
	    RECT 31.0000 70.8000 31.4000 71.2000 ;
	    RECT 37.4000 71.1000 37.8000 71.2000 ;
	    RECT 43.0000 71.1000 43.4000 71.2000 ;
	    RECT 37.4000 70.8000 43.4000 71.1000 ;
	    RECT 55.8000 71.1000 56.2000 71.2000 ;
	    RECT 62.2000 71.1000 62.6000 71.2000 ;
	    RECT 67.8000 71.1000 68.2000 71.2000 ;
	    RECT 73.4000 71.1000 73.8000 71.2000 ;
	    RECT 55.8000 70.8000 73.8000 71.1000 ;
	    RECT 79.0000 70.8000 79.4000 71.2000 ;
	    RECT 83.8000 71.1000 84.2000 71.2000 ;
	    RECT 98.2000 71.1000 98.6000 71.2000 ;
	    RECT 83.8000 70.8000 98.6000 71.1000 ;
	    RECT 120.6000 71.1000 121.0000 71.2000 ;
	    RECT 125.4000 71.1000 125.8000 71.2000 ;
	    RECT 120.6000 70.8000 125.8000 71.1000 ;
	    RECT 135.0000 71.1000 135.4000 71.2000 ;
	    RECT 143.8000 71.1000 144.2000 71.2000 ;
	    RECT 135.0000 70.8000 144.2000 71.1000 ;
	    RECT 182.2000 71.1000 182.6000 71.2000 ;
	    RECT 195.8000 71.1000 196.2000 71.2000 ;
	    RECT 182.2000 70.8000 196.2000 71.1000 ;
	    RECT 203.8000 71.1000 204.2000 71.2000 ;
	    RECT 205.4000 71.1000 205.8000 71.2000 ;
	    RECT 203.8000 70.8000 205.8000 71.1000 ;
	    RECT 223.8000 71.1000 224.2000 71.2000 ;
	    RECT 227.0000 71.1000 227.4000 71.2000 ;
	    RECT 223.8000 70.8000 227.4000 71.1000 ;
	    RECT 228.6000 71.1000 229.0000 71.2000 ;
	    RECT 234.2000 71.1000 234.6000 71.2000 ;
	    RECT 228.6000 70.8000 234.6000 71.1000 ;
	    RECT 265.4000 71.1000 265.8000 71.2000 ;
	    RECT 267.8000 71.1000 268.2000 71.2000 ;
	    RECT 265.4000 70.8000 268.2000 71.1000 ;
	    RECT 31.0000 70.2000 31.3000 70.8000 ;
	    RECT 31.0000 69.8000 31.4000 70.2000 ;
	    RECT 56.6000 70.1000 57.0000 70.2000 ;
	    RECT 71.8000 70.1000 72.2000 70.2000 ;
	    RECT 56.6000 69.8000 72.2000 70.1000 ;
	    RECT 89.4000 70.1000 89.8000 70.2000 ;
	    RECT 99.0000 70.1000 99.4000 70.2000 ;
	    RECT 89.4000 69.8000 99.4000 70.1000 ;
	    RECT 117.4000 70.1000 117.8000 70.2000 ;
	    RECT 123.0000 70.1000 123.4000 70.2000 ;
	    RECT 117.4000 69.8000 123.4000 70.1000 ;
	    RECT 191.0000 70.1000 191.4000 70.2000 ;
	    RECT 202.2000 70.1000 202.6000 70.2000 ;
	    RECT 191.0000 69.8000 202.6000 70.1000 ;
	    RECT 206.2000 70.1000 206.6000 70.2000 ;
	    RECT 219.8000 70.1000 220.2000 70.2000 ;
	    RECT 237.4000 70.1000 237.8000 70.2000 ;
	    RECT 243.8000 70.1000 244.2000 70.2000 ;
	    RECT 206.2000 69.8000 209.7000 70.1000 ;
	    RECT 219.8000 69.8000 244.2000 70.1000 ;
	    RECT 18.2000 68.8000 18.6000 69.2000 ;
	    RECT 24.6000 68.8000 25.0000 69.2000 ;
	    RECT 25.4000 69.1000 25.8000 69.2000 ;
	    RECT 27.0000 69.1000 27.4000 69.2000 ;
	    RECT 29.4000 69.1000 29.8000 69.2000 ;
	    RECT 25.4000 68.8000 29.8000 69.1000 ;
	    RECT 43.0000 69.1000 43.4000 69.2000 ;
	    RECT 47.8000 69.1000 48.2000 69.2000 ;
	    RECT 43.0000 68.8000 48.2000 69.1000 ;
	    RECT 75.0000 69.1000 75.4000 69.2000 ;
	    RECT 75.8000 69.1000 76.2000 69.2000 ;
	    RECT 84.6000 69.1000 85.0000 69.2000 ;
	    RECT 96.6000 69.1000 97.0000 69.2000 ;
	    RECT 75.0000 68.8000 97.0000 69.1000 ;
	    RECT 107.8000 69.1000 108.2000 69.2000 ;
	    RECT 135.0000 69.1000 135.4000 69.2000 ;
	    RECT 138.2000 69.1000 138.6000 69.2000 ;
	    RECT 107.8000 68.8000 138.6000 69.1000 ;
	    RECT 139.8000 69.1000 140.2000 69.2000 ;
	    RECT 144.6000 69.1000 145.0000 69.2000 ;
	    RECT 151.0000 69.1000 151.4000 69.2000 ;
	    RECT 139.8000 68.8000 151.4000 69.1000 ;
	    RECT 194.2000 69.1000 194.6000 69.2000 ;
	    RECT 204.6000 69.1000 205.0000 69.2000 ;
	    RECT 194.2000 68.8000 205.0000 69.1000 ;
	    RECT 205.4000 69.1000 205.8000 69.2000 ;
	    RECT 208.6000 69.1000 209.0000 69.2000 ;
	    RECT 205.4000 68.8000 209.0000 69.1000 ;
	    RECT 209.4000 69.1000 209.7000 69.8000 ;
	    RECT 224.6000 69.1000 225.0000 69.2000 ;
	    RECT 209.4000 68.8000 225.0000 69.1000 ;
	    RECT 227.0000 69.1000 227.4000 69.2000 ;
	    RECT 232.6000 69.1000 233.0000 69.2000 ;
	    RECT 227.0000 68.8000 233.0000 69.1000 ;
	    RECT 18.2000 68.2000 18.5000 68.8000 ;
	    RECT 18.2000 67.8000 18.6000 68.2000 ;
	    RECT 23.0000 68.1000 23.4000 68.2000 ;
	    RECT 24.6000 68.1000 24.9000 68.8000 ;
	    RECT 23.0000 67.8000 24.9000 68.1000 ;
	    RECT 28.6000 67.8000 29.0000 68.2000 ;
	    RECT 36.6000 67.8000 37.0000 68.2000 ;
	    RECT 39.0000 68.1000 39.4000 68.2000 ;
	    RECT 41.4000 68.1000 41.8000 68.2000 ;
	    RECT 45.4000 68.1000 45.8000 68.2000 ;
	    RECT 55.0000 68.1000 55.4000 68.2000 ;
	    RECT 93.4000 68.1000 93.8000 68.2000 ;
	    RECT 125.4000 68.1000 125.8000 68.2000 ;
	    RECT 127.8000 68.1000 128.2000 68.2000 ;
	    RECT 39.0000 67.8000 128.2000 68.1000 ;
	    RECT 135.0000 68.1000 135.4000 68.2000 ;
	    RECT 165.4000 68.1000 165.8000 68.2000 ;
	    RECT 135.0000 67.8000 165.8000 68.1000 ;
	    RECT 173.4000 68.1000 173.8000 68.2000 ;
	    RECT 176.6000 68.1000 177.0000 68.2000 ;
	    RECT 173.4000 67.8000 177.0000 68.1000 ;
	    RECT 200.6000 68.1000 201.0000 68.2000 ;
	    RECT 219.8000 68.1000 220.2000 68.2000 ;
	    RECT 242.2000 68.1000 242.6000 68.2000 ;
	    RECT 249.4000 68.1000 249.8000 68.2000 ;
	    RECT 200.6000 67.8000 249.8000 68.1000 ;
	    RECT 255.0000 68.1000 255.4000 68.2000 ;
	    RECT 257.4000 68.1000 257.8000 68.2000 ;
	    RECT 255.0000 67.8000 257.8000 68.1000 ;
	    RECT 8.6000 67.1000 9.0000 67.2000 ;
	    RECT 9.4000 67.1000 9.8000 67.2000 ;
	    RECT 8.6000 66.8000 9.8000 67.1000 ;
	    RECT 15.0000 67.1000 15.4000 67.2000 ;
	    RECT 18.2000 67.1000 18.6000 67.2000 ;
	    RECT 15.0000 66.8000 18.6000 67.1000 ;
	    RECT 22.2000 66.8000 22.6000 67.2000 ;
	    RECT 28.6000 67.1000 28.9000 67.8000 ;
	    RECT 31.0000 67.1000 31.4000 67.2000 ;
	    RECT 28.6000 66.8000 31.4000 67.1000 ;
	    RECT 34.2000 67.1000 34.6000 67.2000 ;
	    RECT 36.6000 67.1000 36.9000 67.8000 ;
	    RECT 34.2000 66.8000 36.9000 67.1000 ;
	    RECT 42.2000 67.1000 42.6000 67.2000 ;
	    RECT 47.8000 67.1000 48.2000 67.2000 ;
	    RECT 42.2000 66.8000 48.2000 67.1000 ;
	    RECT 53.4000 67.1000 53.8000 67.2000 ;
	    RECT 59.8000 67.1000 60.2000 67.2000 ;
	    RECT 53.4000 66.8000 60.2000 67.1000 ;
	    RECT 61.4000 67.1000 61.8000 67.2000 ;
	    RECT 66.2000 67.1000 66.6000 67.2000 ;
	    RECT 61.4000 66.8000 66.6000 67.1000 ;
	    RECT 69.4000 67.1000 69.8000 67.2000 ;
	    RECT 79.8000 67.1000 80.2000 67.2000 ;
	    RECT 85.4000 67.1000 85.8000 67.2000 ;
	    RECT 101.4000 67.1000 101.8000 67.2000 ;
	    RECT 69.4000 66.8000 101.8000 67.1000 ;
	    RECT 111.8000 67.1000 112.2000 67.2000 ;
	    RECT 119.0000 67.1000 119.4000 67.2000 ;
	    RECT 111.8000 66.8000 119.4000 67.1000 ;
	    RECT 123.8000 67.1000 124.2000 67.2000 ;
	    RECT 127.0000 67.1000 127.4000 67.2000 ;
	    RECT 133.4000 67.1000 133.8000 67.2000 ;
	    RECT 140.6000 67.1000 141.0000 67.2000 ;
	    RECT 144.6000 67.1000 145.0000 67.2000 ;
	    RECT 123.8000 66.8000 145.0000 67.1000 ;
	    RECT 152.6000 67.1000 153.0000 67.2000 ;
	    RECT 155.0000 67.1000 155.4000 67.2000 ;
	    RECT 152.6000 66.8000 155.4000 67.1000 ;
	    RECT 175.8000 67.1000 176.2000 67.2000 ;
	    RECT 179.0000 67.1000 179.4000 67.2000 ;
	    RECT 183.8000 67.1000 184.2000 67.2000 ;
	    RECT 175.8000 66.8000 184.2000 67.1000 ;
	    RECT 186.2000 67.1000 186.6000 67.2000 ;
	    RECT 190.2000 67.1000 190.6000 67.2000 ;
	    RECT 186.2000 66.8000 190.6000 67.1000 ;
	    RECT 191.8000 67.1000 192.2000 67.2000 ;
	    RECT 193.4000 67.1000 193.8000 67.2000 ;
	    RECT 214.2000 67.1000 214.6000 67.2000 ;
	    RECT 191.8000 66.8000 214.6000 67.1000 ;
	    RECT 215.0000 67.1000 215.4000 67.2000 ;
	    RECT 223.0000 67.1000 223.4000 67.2000 ;
	    RECT 215.0000 66.8000 223.4000 67.1000 ;
	    RECT 233.4000 67.1000 233.8000 67.2000 ;
	    RECT 235.8000 67.1000 236.2000 67.2000 ;
	    RECT 233.4000 66.8000 236.2000 67.1000 ;
	    RECT 238.2000 67.1000 238.6000 67.2000 ;
	    RECT 245.4000 67.1000 245.8000 67.2000 ;
	    RECT 247.8000 67.1000 248.2000 67.2000 ;
	    RECT 238.2000 66.8000 245.8000 67.1000 ;
	    RECT 246.2000 66.8000 248.2000 67.1000 ;
	    RECT 251.0000 66.8000 251.4000 67.2000 ;
	    RECT 257.4000 67.1000 257.7000 67.8000 ;
	    RECT 263.0000 67.1000 263.4000 67.2000 ;
	    RECT 257.4000 66.8000 263.4000 67.1000 ;
	    RECT 266.2000 66.8000 266.6000 67.2000 ;
	    RECT 22.2000 66.2000 22.5000 66.8000 ;
	    RECT 3.8000 65.8000 4.2000 66.2000 ;
	    RECT 4.6000 66.1000 5.0000 66.2000 ;
	    RECT 8.6000 66.1000 9.0000 66.2000 ;
	    RECT 4.6000 65.8000 9.0000 66.1000 ;
	    RECT 19.8000 66.1000 20.2000 66.2000 ;
	    RECT 20.6000 66.1000 21.0000 66.2000 ;
	    RECT 19.8000 65.8000 21.0000 66.1000 ;
	    RECT 22.2000 65.8000 22.6000 66.2000 ;
	    RECT 25.4000 66.1000 25.8000 66.2000 ;
	    RECT 28.6000 66.1000 29.0000 66.2000 ;
	    RECT 25.4000 65.8000 29.0000 66.1000 ;
	    RECT 35.8000 66.1000 36.2000 66.2000 ;
	    RECT 38.2000 66.1000 38.6000 66.2000 ;
	    RECT 51.0000 66.1000 51.4000 66.2000 ;
	    RECT 60.6000 66.1000 61.0000 66.2000 ;
	    RECT 68.6000 66.1000 69.0000 66.2000 ;
	    RECT 79.0000 66.1000 79.4000 66.2000 ;
	    RECT 82.2000 66.1000 82.6000 66.2000 ;
	    RECT 35.8000 65.8000 82.6000 66.1000 ;
	    RECT 88.6000 66.1000 89.0000 66.2000 ;
	    RECT 90.2000 66.1000 90.6000 66.2000 ;
	    RECT 88.6000 65.8000 90.6000 66.1000 ;
	    RECT 97.4000 66.1000 97.8000 66.2000 ;
	    RECT 98.2000 66.1000 98.6000 66.2000 ;
	    RECT 97.4000 65.8000 98.6000 66.1000 ;
	    RECT 99.8000 66.1000 100.2000 66.2000 ;
	    RECT 105.4000 66.1000 105.8000 66.2000 ;
	    RECT 112.6000 66.1000 113.0000 66.2000 ;
	    RECT 120.6000 66.1000 121.0000 66.2000 ;
	    RECT 99.8000 65.8000 113.0000 66.1000 ;
	    RECT 118.2000 65.8000 121.0000 66.1000 ;
	    RECT 127.0000 66.1000 127.4000 66.2000 ;
	    RECT 139.8000 66.1000 140.2000 66.2000 ;
	    RECT 145.4000 66.1000 145.8000 66.2000 ;
	    RECT 127.0000 65.8000 145.8000 66.1000 ;
	    RECT 151.0000 66.1000 151.4000 66.2000 ;
	    RECT 180.6000 66.1000 181.0000 66.2000 ;
	    RECT 186.2000 66.1000 186.6000 66.2000 ;
	    RECT 188.6000 66.1000 189.0000 66.2000 ;
	    RECT 191.8000 66.1000 192.2000 66.2000 ;
	    RECT 151.0000 65.8000 156.1000 66.1000 ;
	    RECT 180.6000 65.8000 192.2000 66.1000 ;
	    RECT 199.0000 66.1000 199.4000 66.2000 ;
	    RECT 211.8000 66.1000 212.2000 66.2000 ;
	    RECT 199.0000 65.8000 212.2000 66.1000 ;
	    RECT 213.4000 66.1000 213.8000 66.2000 ;
	    RECT 215.8000 66.1000 216.2000 66.2000 ;
	    RECT 219.8000 66.1000 220.2000 66.2000 ;
	    RECT 213.4000 65.8000 220.2000 66.1000 ;
	    RECT 228.6000 65.8000 229.0000 66.2000 ;
	    RECT 229.4000 65.8000 229.8000 66.2000 ;
	    RECT 237.4000 66.1000 237.8000 66.2000 ;
	    RECT 238.2000 66.1000 238.6000 66.2000 ;
	    RECT 237.4000 65.8000 238.6000 66.1000 ;
	    RECT 241.4000 66.1000 241.8000 66.2000 ;
	    RECT 246.2000 66.1000 246.5000 66.8000 ;
	    RECT 241.4000 65.8000 246.5000 66.1000 ;
	    RECT 247.8000 66.1000 248.2000 66.2000 ;
	    RECT 248.6000 66.1000 249.0000 66.2000 ;
	    RECT 247.8000 65.8000 249.0000 66.1000 ;
	    RECT 251.0000 66.1000 251.3000 66.8000 ;
	    RECT 266.2000 66.2000 266.5000 66.8000 ;
	    RECT 266.2000 66.1000 266.6000 66.2000 ;
	    RECT 251.0000 65.8000 266.6000 66.1000 ;
	    RECT 2.2000 65.1000 2.6000 65.2000 ;
	    RECT 3.8000 65.1000 4.1000 65.8000 ;
	    RECT 118.2000 65.2000 118.5000 65.8000 ;
	    RECT 155.8000 65.2000 156.1000 65.8000 ;
	    RECT 228.6000 65.2000 228.9000 65.8000 ;
	    RECT 229.4000 65.2000 229.7000 65.8000 ;
	    RECT 2.2000 64.8000 4.1000 65.1000 ;
	    RECT 7.8000 65.1000 8.2000 65.2000 ;
	    RECT 9.4000 65.1000 9.8000 65.2000 ;
	    RECT 15.8000 65.1000 16.2000 65.2000 ;
	    RECT 7.8000 64.8000 16.2000 65.1000 ;
	    RECT 19.8000 65.1000 20.2000 65.2000 ;
	    RECT 26.2000 65.1000 26.6000 65.2000 ;
	    RECT 19.8000 64.8000 26.6000 65.1000 ;
	    RECT 31.8000 64.8000 32.2000 65.2000 ;
	    RECT 35.8000 65.1000 36.2000 65.2000 ;
	    RECT 42.2000 65.1000 42.6000 65.2000 ;
	    RECT 35.8000 64.8000 42.6000 65.1000 ;
	    RECT 44.6000 65.1000 45.0000 65.2000 ;
	    RECT 45.4000 65.1000 45.8000 65.2000 ;
	    RECT 44.6000 64.8000 45.8000 65.1000 ;
	    RECT 64.6000 65.1000 65.0000 65.2000 ;
	    RECT 65.4000 65.1000 65.8000 65.2000 ;
	    RECT 89.4000 65.1000 89.8000 65.2000 ;
	    RECT 64.6000 64.8000 89.8000 65.1000 ;
	    RECT 92.6000 64.8000 93.0000 65.2000 ;
	    RECT 104.6000 65.1000 105.0000 65.2000 ;
	    RECT 107.8000 65.1000 108.2000 65.2000 ;
	    RECT 104.6000 64.8000 108.2000 65.1000 ;
	    RECT 114.2000 64.8000 114.6000 65.2000 ;
	    RECT 118.2000 64.8000 118.6000 65.2000 ;
	    RECT 147.8000 64.8000 148.2000 65.2000 ;
	    RECT 155.8000 64.8000 156.2000 65.2000 ;
	    RECT 228.6000 64.8000 229.0000 65.2000 ;
	    RECT 229.4000 64.8000 229.8000 65.2000 ;
	    RECT 236.6000 65.1000 237.0000 65.2000 ;
	    RECT 250.2000 65.1000 250.6000 65.2000 ;
	    RECT 252.6000 65.1000 253.0000 65.2000 ;
	    RECT 236.6000 64.8000 253.0000 65.1000 ;
	    RECT 31.8000 64.2000 32.1000 64.8000 ;
	    RECT 8.6000 63.8000 9.0000 64.2000 ;
	    RECT 11.8000 64.1000 12.2000 64.2000 ;
	    RECT 19.0000 64.1000 19.4000 64.2000 ;
	    RECT 11.8000 63.8000 19.4000 64.1000 ;
	    RECT 31.8000 63.8000 32.2000 64.2000 ;
	    RECT 39.8000 64.1000 40.2000 64.2000 ;
	    RECT 43.8000 64.1000 44.2000 64.2000 ;
	    RECT 39.8000 63.8000 44.2000 64.1000 ;
	    RECT 59.8000 64.1000 60.2000 64.2000 ;
	    RECT 63.8000 64.1000 64.2000 64.2000 ;
	    RECT 59.8000 63.8000 64.2000 64.1000 ;
	    RECT 71.0000 64.1000 71.4000 64.2000 ;
	    RECT 71.8000 64.1000 72.2000 64.2000 ;
	    RECT 71.0000 63.8000 72.2000 64.1000 ;
	    RECT 82.2000 64.1000 82.6000 64.2000 ;
	    RECT 88.6000 64.1000 89.0000 64.2000 ;
	    RECT 82.2000 63.8000 89.0000 64.1000 ;
	    RECT 91.0000 64.1000 91.4000 64.2000 ;
	    RECT 92.6000 64.1000 92.9000 64.8000 ;
	    RECT 91.0000 63.8000 92.9000 64.1000 ;
	    RECT 105.4000 63.8000 105.8000 64.2000 ;
	    RECT 114.2000 64.1000 114.5000 64.8000 ;
	    RECT 123.8000 64.1000 124.2000 64.2000 ;
	    RECT 127.0000 64.1000 127.4000 64.2000 ;
	    RECT 114.2000 63.8000 127.4000 64.1000 ;
	    RECT 129.4000 64.1000 129.8000 64.2000 ;
	    RECT 147.8000 64.1000 148.1000 64.8000 ;
	    RECT 151.0000 64.1000 151.4000 64.2000 ;
	    RECT 129.4000 63.8000 151.4000 64.1000 ;
	    RECT 211.8000 64.1000 212.2000 64.2000 ;
	    RECT 215.0000 64.1000 215.4000 64.2000 ;
	    RECT 211.8000 63.8000 215.4000 64.1000 ;
	    RECT 235.8000 64.1000 236.2000 64.2000 ;
	    RECT 251.8000 64.1000 252.2000 64.2000 ;
	    RECT 235.8000 63.8000 252.2000 64.1000 ;
	    RECT 8.6000 63.2000 8.9000 63.8000 ;
	    RECT 8.6000 62.8000 9.0000 63.2000 ;
	    RECT 71.8000 63.1000 72.2000 63.2000 ;
	    RECT 75.0000 63.1000 75.4000 63.2000 ;
	    RECT 71.0000 62.8000 75.4000 63.1000 ;
	    RECT 78.2000 63.1000 78.6000 63.2000 ;
	    RECT 84.6000 63.1000 85.0000 63.2000 ;
	    RECT 78.2000 62.8000 85.0000 63.1000 ;
	    RECT 105.4000 63.1000 105.7000 63.8000 ;
	    RECT 111.0000 63.1000 111.4000 63.2000 ;
	    RECT 117.4000 63.1000 117.8000 63.2000 ;
	    RECT 248.6000 63.1000 249.0000 63.2000 ;
	    RECT 105.4000 62.8000 117.8000 63.1000 ;
	    RECT 244.6000 62.8000 249.0000 63.1000 ;
	    RECT 244.6000 62.2000 244.9000 62.8000 ;
	    RECT 48.6000 62.1000 49.0000 62.2000 ;
	    RECT 99.0000 62.1000 99.4000 62.2000 ;
	    RECT 48.6000 61.8000 99.4000 62.1000 ;
	    RECT 116.6000 62.1000 117.0000 62.2000 ;
	    RECT 130.2000 62.1000 130.6000 62.2000 ;
	    RECT 116.6000 61.8000 130.6000 62.1000 ;
	    RECT 135.0000 62.1000 135.4000 62.2000 ;
	    RECT 142.2000 62.1000 142.6000 62.2000 ;
	    RECT 159.0000 62.1000 159.4000 62.2000 ;
	    RECT 135.0000 61.8000 159.4000 62.1000 ;
	    RECT 229.4000 62.1000 229.8000 62.2000 ;
	    RECT 231.0000 62.1000 231.4000 62.2000 ;
	    RECT 235.8000 62.1000 236.2000 62.2000 ;
	    RECT 229.4000 61.8000 236.2000 62.1000 ;
	    RECT 244.6000 61.8000 245.0000 62.2000 ;
	    RECT 63.0000 61.1000 63.4000 61.2000 ;
	    RECT 71.8000 61.1000 72.2000 61.2000 ;
	    RECT 63.0000 60.8000 72.2000 61.1000 ;
	    RECT 95.0000 61.1000 95.4000 61.2000 ;
	    RECT 127.8000 61.1000 128.2000 61.2000 ;
	    RECT 95.0000 60.8000 128.2000 61.1000 ;
	    RECT 98.2000 60.1000 98.6000 60.2000 ;
	    RECT 131.8000 60.1000 132.2000 60.2000 ;
	    RECT 98.2000 59.8000 132.2000 60.1000 ;
	    RECT 163.0000 60.1000 163.4000 60.2000 ;
	    RECT 181.4000 60.1000 181.8000 60.2000 ;
	    RECT 163.0000 59.8000 181.8000 60.1000 ;
	    RECT 192.6000 59.8000 193.0000 60.2000 ;
	    RECT 33.4000 59.1000 33.8000 59.2000 ;
	    RECT 43.8000 59.1000 44.2000 59.2000 ;
	    RECT 49.4000 59.1000 49.8000 59.2000 ;
	    RECT 54.2000 59.1000 54.6000 59.2000 ;
	    RECT 33.4000 58.8000 54.6000 59.1000 ;
	    RECT 65.4000 59.1000 65.8000 59.2000 ;
	    RECT 80.6000 59.1000 81.0000 59.2000 ;
	    RECT 90.2000 59.1000 90.6000 59.2000 ;
	    RECT 65.4000 58.8000 90.6000 59.1000 ;
	    RECT 110.2000 59.1000 110.6000 59.2000 ;
	    RECT 122.2000 59.1000 122.6000 59.2000 ;
	    RECT 110.2000 58.8000 122.6000 59.1000 ;
	    RECT 142.2000 59.1000 142.6000 59.2000 ;
	    RECT 143.8000 59.1000 144.2000 59.2000 ;
	    RECT 142.2000 58.8000 144.2000 59.1000 ;
	    RECT 159.0000 59.1000 159.4000 59.2000 ;
	    RECT 165.4000 59.1000 165.8000 59.2000 ;
	    RECT 167.8000 59.1000 168.2000 59.2000 ;
	    RECT 159.0000 58.8000 168.2000 59.1000 ;
	    RECT 192.6000 59.1000 192.9000 59.8000 ;
	    RECT 194.2000 59.1000 194.6000 59.2000 ;
	    RECT 192.6000 58.8000 194.6000 59.1000 ;
	    RECT 235.0000 59.1000 235.4000 59.2000 ;
	    RECT 239.8000 59.1000 240.2000 59.2000 ;
	    RECT 235.0000 58.8000 240.2000 59.1000 ;
	    RECT 29.4000 58.1000 29.8000 58.2000 ;
	    RECT 104.6000 58.1000 105.0000 58.2000 ;
	    RECT 29.4000 57.8000 105.0000 58.1000 ;
	    RECT 108.6000 58.1000 109.0000 58.2000 ;
	    RECT 112.6000 58.1000 113.0000 58.2000 ;
	    RECT 108.6000 57.8000 113.0000 58.1000 ;
	    RECT 123.0000 58.1000 123.4000 58.2000 ;
	    RECT 145.4000 58.1000 145.8000 58.2000 ;
	    RECT 123.0000 57.8000 145.8000 58.1000 ;
	    RECT 3.8000 56.8000 4.2000 57.2000 ;
	    RECT 30.2000 56.8000 30.6000 57.2000 ;
	    RECT 52.6000 56.8000 53.0000 57.2000 ;
	    RECT 66.2000 57.1000 66.6000 57.2000 ;
	    RECT 69.4000 57.1000 69.8000 57.2000 ;
	    RECT 66.2000 56.8000 69.8000 57.1000 ;
	    RECT 103.0000 57.1000 103.4000 57.2000 ;
	    RECT 106.2000 57.1000 106.6000 57.2000 ;
	    RECT 103.0000 56.8000 106.6000 57.1000 ;
	    RECT 120.6000 57.1000 121.0000 57.2000 ;
	    RECT 123.8000 57.1000 124.2000 57.2000 ;
	    RECT 120.6000 56.8000 124.2000 57.1000 ;
	    RECT 127.8000 57.1000 128.2000 57.2000 ;
	    RECT 132.6000 57.1000 133.0000 57.2000 ;
	    RECT 127.8000 56.8000 133.0000 57.1000 ;
	    RECT 144.6000 57.1000 145.0000 57.2000 ;
	    RECT 147.8000 57.1000 148.2000 57.2000 ;
	    RECT 144.6000 56.8000 148.2000 57.1000 ;
	    RECT 175.8000 57.1000 176.2000 57.2000 ;
	    RECT 180.6000 57.1000 181.0000 57.2000 ;
	    RECT 175.8000 56.8000 181.0000 57.1000 ;
	    RECT 183.0000 57.1000 183.4000 57.2000 ;
	    RECT 191.0000 57.1000 191.4000 57.2000 ;
	    RECT 183.0000 56.8000 191.4000 57.1000 ;
	    RECT 240.6000 57.1000 241.0000 57.2000 ;
	    RECT 243.0000 57.1000 243.4000 57.2000 ;
	    RECT 240.6000 56.8000 243.4000 57.1000 ;
	    RECT 261.4000 56.8000 261.8000 57.2000 ;
	    RECT 3.8000 56.1000 4.1000 56.8000 ;
	    RECT 11.0000 56.1000 11.4000 56.2000 ;
	    RECT 3.8000 55.8000 11.4000 56.1000 ;
	    RECT 13.4000 55.8000 13.8000 56.2000 ;
	    RECT 20.6000 56.1000 21.0000 56.2000 ;
	    RECT 30.2000 56.1000 30.5000 56.8000 ;
	    RECT 20.6000 55.8000 30.5000 56.1000 ;
	    RECT 49.4000 56.1000 49.8000 56.2000 ;
	    RECT 52.6000 56.1000 52.9000 56.8000 ;
	    RECT 49.4000 55.8000 52.9000 56.1000 ;
	    RECT 79.8000 55.8000 80.2000 56.2000 ;
	    RECT 99.0000 56.1000 99.4000 56.2000 ;
	    RECT 103.0000 56.1000 103.4000 56.2000 ;
	    RECT 99.0000 55.8000 103.4000 56.1000 ;
	    RECT 123.0000 56.1000 123.4000 56.2000 ;
	    RECT 130.2000 56.1000 130.6000 56.2000 ;
	    RECT 146.2000 56.1000 146.6000 56.2000 ;
	    RECT 148.6000 56.1000 149.0000 56.2000 ;
	    RECT 154.2000 56.1000 154.6000 56.2000 ;
	    RECT 123.0000 55.8000 154.6000 56.1000 ;
	    RECT 172.6000 56.1000 173.0000 56.2000 ;
	    RECT 179.0000 56.1000 179.4000 56.2000 ;
	    RECT 172.6000 55.8000 179.4000 56.1000 ;
	    RECT 186.2000 55.8000 186.6000 56.2000 ;
	    RECT 259.8000 56.1000 260.2000 56.2000 ;
	    RECT 261.4000 56.1000 261.7000 56.8000 ;
	    RECT 259.8000 55.8000 261.7000 56.1000 ;
	    RECT 11.0000 55.1000 11.4000 55.2000 ;
	    RECT 13.4000 55.1000 13.7000 55.8000 ;
	    RECT 11.0000 54.8000 13.7000 55.1000 ;
	    RECT 16.6000 55.1000 17.0000 55.2000 ;
	    RECT 17.4000 55.1000 17.8000 55.2000 ;
	    RECT 22.2000 55.1000 22.6000 55.2000 ;
	    RECT 16.6000 54.8000 22.6000 55.1000 ;
	    RECT 32.6000 54.8000 33.0000 55.2000 ;
	    RECT 38.2000 55.1000 38.6000 55.2000 ;
	    RECT 39.8000 55.1000 40.2000 55.2000 ;
	    RECT 38.2000 54.8000 40.2000 55.1000 ;
	    RECT 51.0000 54.8000 51.4000 55.2000 ;
	    RECT 67.8000 55.1000 68.2000 55.2000 ;
	    RECT 63.0000 54.8000 68.2000 55.1000 ;
	    RECT 68.6000 55.1000 69.0000 55.2000 ;
	    RECT 73.4000 55.1000 73.8000 55.2000 ;
	    RECT 77.4000 55.1000 77.8000 55.2000 ;
	    RECT 79.8000 55.1000 80.1000 55.8000 ;
	    RECT 68.6000 54.8000 74.5000 55.1000 ;
	    RECT 77.4000 54.8000 80.1000 55.1000 ;
	    RECT 91.0000 54.8000 91.4000 55.2000 ;
	    RECT 100.6000 55.1000 101.0000 55.2000 ;
	    RECT 102.2000 55.1000 102.6000 55.2000 ;
	    RECT 123.8000 55.1000 124.2000 55.2000 ;
	    RECT 100.6000 54.8000 102.6000 55.1000 ;
	    RECT 115.0000 54.8000 120.1000 55.1000 ;
	    RECT 32.6000 54.2000 32.9000 54.8000 ;
	    RECT 32.6000 53.8000 33.0000 54.2000 ;
	    RECT 36.6000 54.1000 37.0000 54.2000 ;
	    RECT 37.4000 54.1000 37.8000 54.2000 ;
	    RECT 36.6000 53.8000 37.8000 54.1000 ;
	    RECT 51.0000 54.1000 51.3000 54.8000 ;
	    RECT 63.0000 54.7000 63.4000 54.8000 ;
	    RECT 53.4000 54.1000 53.8000 54.2000 ;
	    RECT 62.2000 54.1000 62.6000 54.2000 ;
	    RECT 51.0000 53.8000 62.6000 54.1000 ;
	    RECT 67.0000 54.1000 67.4000 54.2000 ;
	    RECT 79.0000 54.1000 79.4000 54.2000 ;
	    RECT 67.0000 53.8000 79.4000 54.1000 ;
	    RECT 91.0000 54.1000 91.3000 54.8000 ;
	    RECT 115.0000 54.7000 115.4000 54.8000 ;
	    RECT 119.8000 54.2000 120.1000 54.8000 ;
	    RECT 121.4000 54.8000 124.2000 55.1000 ;
	    RECT 125.4000 55.1000 125.8000 55.2000 ;
	    RECT 128.6000 55.1000 129.0000 55.2000 ;
	    RECT 130.2000 55.1000 130.6000 55.2000 ;
	    RECT 132.6000 55.1000 133.0000 55.2000 ;
	    RECT 125.4000 54.8000 130.6000 55.1000 ;
	    RECT 131.8000 54.8000 133.0000 55.1000 ;
	    RECT 134.2000 55.1000 134.6000 55.2000 ;
	    RECT 143.8000 55.1000 144.2000 55.2000 ;
	    RECT 162.2000 55.1000 162.6000 55.2000 ;
	    RECT 134.2000 54.8000 138.6000 55.1000 ;
	    RECT 121.4000 54.2000 121.7000 54.8000 ;
	    RECT 112.6000 54.1000 113.0000 54.2000 ;
	    RECT 91.0000 53.8000 113.0000 54.1000 ;
	    RECT 119.8000 53.8000 120.2000 54.2000 ;
	    RECT 121.4000 53.8000 121.8000 54.2000 ;
	    RECT 127.0000 54.1000 127.4000 54.2000 ;
	    RECT 127.8000 54.1000 128.2000 54.2000 ;
	    RECT 131.8000 54.1000 132.1000 54.8000 ;
	    RECT 138.2000 54.7000 138.6000 54.8000 ;
	    RECT 140.6000 54.8000 162.6000 55.1000 ;
	    RECT 167.0000 55.1000 167.4000 55.2000 ;
	    RECT 177.4000 55.1000 177.8000 55.2000 ;
	    RECT 178.2000 55.1000 178.6000 55.2000 ;
	    RECT 167.0000 54.8000 178.6000 55.1000 ;
	    RECT 181.4000 55.1000 181.8000 55.2000 ;
	    RECT 186.2000 55.1000 186.5000 55.8000 ;
	    RECT 181.4000 54.8000 186.5000 55.1000 ;
	    RECT 204.6000 55.1000 205.0000 55.2000 ;
	    RECT 206.2000 55.1000 206.6000 55.2000 ;
	    RECT 204.6000 54.8000 206.6000 55.1000 ;
	    RECT 210.2000 54.8000 210.6000 55.2000 ;
	    RECT 218.2000 55.1000 218.6000 55.2000 ;
	    RECT 228.6000 55.1000 229.0000 55.2000 ;
	    RECT 231.0000 55.1000 231.4000 55.2000 ;
	    RECT 218.2000 54.8000 231.4000 55.1000 ;
	    RECT 233.4000 55.1000 233.8000 55.2000 ;
	    RECT 260.6000 55.1000 261.0000 55.2000 ;
	    RECT 233.4000 54.8000 261.0000 55.1000 ;
	    RECT 140.6000 54.2000 140.9000 54.8000 ;
	    RECT 127.0000 53.8000 132.1000 54.1000 ;
	    RECT 132.6000 54.1000 133.0000 54.2000 ;
	    RECT 133.4000 54.1000 133.8000 54.2000 ;
	    RECT 132.6000 53.8000 133.8000 54.1000 ;
	    RECT 140.6000 53.8000 141.0000 54.2000 ;
	    RECT 166.2000 54.1000 166.6000 54.2000 ;
	    RECT 170.2000 54.1000 170.6000 54.2000 ;
	    RECT 166.2000 53.8000 170.6000 54.1000 ;
	    RECT 173.4000 54.1000 173.8000 54.2000 ;
	    RECT 174.2000 54.1000 174.6000 54.2000 ;
	    RECT 173.4000 53.8000 174.6000 54.1000 ;
	    RECT 180.6000 54.1000 181.0000 54.2000 ;
	    RECT 181.4000 54.1000 181.8000 54.2000 ;
	    RECT 205.4000 54.1000 205.8000 54.2000 ;
	    RECT 210.2000 54.1000 210.5000 54.8000 ;
	    RECT 180.6000 53.8000 181.8000 54.1000 ;
	    RECT 204.6000 53.8000 210.5000 54.1000 ;
	    RECT 216.6000 54.1000 217.0000 54.2000 ;
	    RECT 244.6000 54.1000 245.0000 54.2000 ;
	    RECT 257.4000 54.1000 257.8000 54.2000 ;
	    RECT 216.6000 53.8000 257.8000 54.1000 ;
	    RECT 258.2000 53.8000 258.6000 54.2000 ;
	    RECT 259.8000 54.1000 260.2000 54.2000 ;
	    RECT 266.2000 54.1000 266.6000 54.2000 ;
	    RECT 259.8000 53.8000 266.6000 54.1000 ;
	    RECT 35.0000 53.1000 35.4000 53.2000 ;
	    RECT 38.2000 53.1000 38.6000 53.2000 ;
	    RECT 35.0000 52.8000 38.6000 53.1000 ;
	    RECT 39.0000 52.8000 39.4000 53.2000 ;
	    RECT 81.4000 53.1000 81.8000 53.2000 ;
	    RECT 82.2000 53.1000 82.6000 53.2000 ;
	    RECT 124.6000 53.1000 125.0000 53.2000 ;
	    RECT 127.8000 53.1000 128.2000 53.2000 ;
	    RECT 129.4000 53.1000 129.8000 53.2000 ;
	    RECT 81.4000 52.8000 93.7000 53.1000 ;
	    RECT 124.6000 52.8000 129.8000 53.1000 ;
	    RECT 131.8000 53.1000 132.2000 53.2000 ;
	    RECT 133.4000 53.1000 133.8000 53.2000 ;
	    RECT 131.8000 52.8000 133.8000 53.1000 ;
	    RECT 156.6000 53.1000 157.0000 53.2000 ;
	    RECT 158.2000 53.1000 158.6000 53.2000 ;
	    RECT 156.6000 52.8000 158.6000 53.1000 ;
	    RECT 175.8000 53.1000 176.2000 53.2000 ;
	    RECT 176.6000 53.1000 177.0000 53.2000 ;
	    RECT 211.8000 53.1000 212.2000 53.2000 ;
	    RECT 175.8000 52.8000 177.0000 53.1000 ;
	    RECT 205.4000 52.8000 212.2000 53.1000 ;
	    RECT 239.0000 53.1000 239.4000 53.2000 ;
	    RECT 251.0000 53.1000 251.4000 53.2000 ;
	    RECT 258.2000 53.1000 258.5000 53.8000 ;
	    RECT 239.0000 52.8000 244.1000 53.1000 ;
	    RECT 251.0000 52.8000 258.5000 53.1000 ;
	    RECT 260.6000 53.1000 261.0000 53.2000 ;
	    RECT 267.0000 53.1000 267.4000 53.2000 ;
	    RECT 260.6000 52.8000 267.4000 53.1000 ;
	    RECT 20.6000 52.1000 21.0000 52.2000 ;
	    RECT 25.4000 52.1000 25.8000 52.2000 ;
	    RECT 20.6000 51.8000 25.8000 52.1000 ;
	    RECT 31.8000 52.1000 32.2000 52.2000 ;
	    RECT 39.0000 52.1000 39.3000 52.8000 ;
	    RECT 93.4000 52.2000 93.7000 52.8000 ;
	    RECT 205.4000 52.2000 205.7000 52.8000 ;
	    RECT 243.8000 52.2000 244.1000 52.8000 ;
	    RECT 31.8000 51.8000 39.3000 52.1000 ;
	    RECT 61.4000 52.1000 61.8000 52.2000 ;
	    RECT 69.4000 52.1000 69.8000 52.2000 ;
	    RECT 61.4000 51.8000 69.8000 52.1000 ;
	    RECT 93.4000 51.8000 93.8000 52.2000 ;
	    RECT 173.4000 52.1000 173.8000 52.2000 ;
	    RECT 176.6000 52.1000 177.0000 52.2000 ;
	    RECT 180.6000 52.1000 181.0000 52.2000 ;
	    RECT 173.4000 51.8000 181.0000 52.1000 ;
	    RECT 205.4000 51.8000 205.8000 52.2000 ;
	    RECT 219.0000 52.1000 219.4000 52.2000 ;
	    RECT 230.2000 52.1000 230.6000 52.2000 ;
	    RECT 219.0000 51.8000 230.6000 52.1000 ;
	    RECT 243.8000 51.8000 244.2000 52.2000 ;
	    RECT 251.8000 52.1000 252.2000 52.2000 ;
	    RECT 255.0000 52.1000 255.4000 52.2000 ;
	    RECT 251.8000 51.8000 255.4000 52.1000 ;
	    RECT 57.4000 51.1000 57.8000 51.2000 ;
	    RECT 69.4000 51.1000 69.8000 51.2000 ;
	    RECT 71.8000 51.1000 72.2000 51.2000 ;
	    RECT 57.4000 50.8000 72.2000 51.1000 ;
	    RECT 89.4000 51.1000 89.8000 51.2000 ;
	    RECT 94.2000 51.1000 94.6000 51.2000 ;
	    RECT 89.4000 50.8000 94.6000 51.1000 ;
	    RECT 170.2000 51.1000 170.6000 51.2000 ;
	    RECT 187.8000 51.1000 188.2000 51.2000 ;
	    RECT 170.2000 50.8000 188.2000 51.1000 ;
	    RECT 189.4000 51.1000 189.8000 51.2000 ;
	    RECT 195.8000 51.1000 196.2000 51.2000 ;
	    RECT 198.2000 51.1000 198.6000 51.2000 ;
	    RECT 189.4000 50.8000 198.6000 51.1000 ;
	    RECT 199.8000 51.1000 200.2000 51.2000 ;
	    RECT 207.0000 51.1000 207.4000 51.2000 ;
	    RECT 199.8000 50.8000 207.4000 51.1000 ;
	    RECT 227.0000 51.1000 227.4000 51.2000 ;
	    RECT 229.4000 51.1000 229.8000 51.2000 ;
	    RECT 227.0000 50.8000 229.8000 51.1000 ;
	    RECT 255.0000 51.1000 255.4000 51.2000 ;
	    RECT 259.8000 51.1000 260.2000 51.2000 ;
	    RECT 255.0000 50.8000 260.2000 51.1000 ;
	    RECT 40.6000 50.1000 41.0000 50.2000 ;
	    RECT 42.2000 50.1000 42.6000 50.2000 ;
	    RECT 40.6000 49.8000 42.6000 50.1000 ;
	    RECT 66.2000 50.1000 66.6000 50.2000 ;
	    RECT 71.8000 50.1000 72.2000 50.2000 ;
	    RECT 66.2000 49.8000 72.2000 50.1000 ;
	    RECT 79.0000 50.1000 79.4000 50.2000 ;
	    RECT 157.4000 50.1000 157.8000 50.2000 ;
	    RECT 159.8000 50.1000 160.2000 50.2000 ;
	    RECT 79.0000 49.8000 92.1000 50.1000 ;
	    RECT 157.4000 49.8000 160.2000 50.1000 ;
	    RECT 227.8000 49.8000 228.2000 50.2000 ;
	    RECT 265.4000 50.1000 265.8000 50.2000 ;
	    RECT 267.8000 50.1000 268.2000 50.2000 ;
	    RECT 265.4000 49.8000 268.2000 50.1000 ;
	    RECT 91.8000 49.2000 92.1000 49.8000 ;
	    RECT 227.8000 49.2000 228.1000 49.8000 ;
	    RECT 3.0000 49.1000 3.4000 49.2000 ;
	    RECT 8.6000 49.1000 9.0000 49.2000 ;
	    RECT 3.0000 48.8000 9.0000 49.1000 ;
	    RECT 43.8000 49.1000 44.2000 49.2000 ;
	    RECT 47.0000 49.1000 47.4000 49.2000 ;
	    RECT 54.2000 49.1000 54.6000 49.2000 ;
	    RECT 43.8000 48.8000 54.6000 49.1000 ;
	    RECT 57.4000 49.1000 57.8000 49.2000 ;
	    RECT 63.8000 49.1000 64.2000 49.2000 ;
	    RECT 57.4000 48.8000 64.2000 49.1000 ;
	    RECT 82.2000 49.1000 82.6000 49.2000 ;
	    RECT 87.8000 49.1000 88.2000 49.2000 ;
	    RECT 82.2000 48.8000 88.2000 49.1000 ;
	    RECT 91.8000 49.1000 92.2000 49.2000 ;
	    RECT 96.6000 49.1000 97.0000 49.2000 ;
	    RECT 101.4000 49.1000 101.8000 49.2000 ;
	    RECT 91.8000 48.8000 101.8000 49.1000 ;
	    RECT 121.4000 49.1000 121.8000 49.2000 ;
	    RECT 122.2000 49.1000 122.6000 49.2000 ;
	    RECT 121.4000 48.8000 122.6000 49.1000 ;
	    RECT 175.8000 48.8000 176.2000 49.2000 ;
	    RECT 227.8000 49.1000 228.2000 49.2000 ;
	    RECT 233.4000 49.1000 233.8000 49.2000 ;
	    RECT 255.0000 49.1000 255.4000 49.2000 ;
	    RECT 227.8000 48.8000 233.8000 49.1000 ;
	    RECT 251.0000 48.8000 255.4000 49.1000 ;
	    RECT 255.8000 49.1000 256.2000 49.2000 ;
	    RECT 263.8000 49.1000 264.2000 49.2000 ;
	    RECT 255.8000 48.8000 264.2000 49.1000 ;
	    RECT 29.4000 48.1000 29.8000 48.2000 ;
	    RECT 30.2000 48.1000 30.6000 48.2000 ;
	    RECT 29.4000 47.8000 30.6000 48.1000 ;
	    RECT 36.6000 48.1000 37.0000 48.2000 ;
	    RECT 37.4000 48.1000 37.8000 48.2000 ;
	    RECT 36.6000 47.8000 37.8000 48.1000 ;
	    RECT 55.8000 48.1000 56.2000 48.2000 ;
	    RECT 57.4000 48.1000 57.7000 48.8000 ;
	    RECT 55.8000 47.8000 57.7000 48.1000 ;
	    RECT 69.4000 48.1000 69.8000 48.2000 ;
	    RECT 70.2000 48.1000 70.6000 48.2000 ;
	    RECT 69.4000 47.8000 70.6000 48.1000 ;
	    RECT 83.0000 48.1000 83.4000 48.2000 ;
	    RECT 89.4000 48.1000 89.8000 48.2000 ;
	    RECT 83.0000 47.8000 89.8000 48.1000 ;
	    RECT 90.2000 48.1000 90.6000 48.2000 ;
	    RECT 92.6000 48.1000 93.0000 48.2000 ;
	    RECT 90.2000 47.8000 93.0000 48.1000 ;
	    RECT 95.8000 48.1000 96.2000 48.2000 ;
	    RECT 99.0000 48.1000 99.4000 48.2000 ;
	    RECT 108.6000 48.1000 109.0000 48.2000 ;
	    RECT 119.0000 48.1000 119.4000 48.2000 ;
	    RECT 95.8000 47.8000 119.4000 48.1000 ;
	    RECT 123.8000 48.1000 124.2000 48.2000 ;
	    RECT 127.0000 48.1000 127.4000 48.2000 ;
	    RECT 123.8000 47.8000 127.4000 48.1000 ;
	    RECT 171.8000 48.1000 172.2000 48.2000 ;
	    RECT 175.8000 48.1000 176.1000 48.8000 ;
	    RECT 251.0000 48.2000 251.3000 48.8000 ;
	    RECT 187.0000 48.1000 187.4000 48.2000 ;
	    RECT 194.2000 48.1000 194.6000 48.2000 ;
	    RECT 206.2000 48.1000 206.6000 48.2000 ;
	    RECT 171.8000 47.8000 206.6000 48.1000 ;
	    RECT 245.4000 48.1000 245.8000 48.2000 ;
	    RECT 250.2000 48.1000 250.6000 48.2000 ;
	    RECT 245.4000 47.8000 250.6000 48.1000 ;
	    RECT 251.0000 47.8000 251.4000 48.2000 ;
	    RECT 253.4000 48.1000 253.8000 48.2000 ;
	    RECT 256.6000 48.1000 257.0000 48.2000 ;
	    RECT 269.4000 48.1000 269.8000 48.2000 ;
	    RECT 253.4000 47.8000 269.8000 48.1000 ;
	    RECT 27.8000 47.1000 28.2000 47.2000 ;
	    RECT 29.4000 47.1000 29.7000 47.8000 ;
	    RECT 27.8000 46.8000 29.7000 47.1000 ;
	    RECT 49.4000 46.8000 49.8000 47.2000 ;
	    RECT 52.6000 46.8000 53.0000 47.2000 ;
	    RECT 63.0000 47.1000 63.4000 47.2000 ;
	    RECT 65.4000 47.1000 65.8000 47.2000 ;
	    RECT 63.0000 46.8000 65.8000 47.1000 ;
	    RECT 75.0000 47.1000 75.4000 47.2000 ;
	    RECT 78.2000 47.1000 78.6000 47.2000 ;
	    RECT 91.0000 47.1000 91.4000 47.2000 ;
	    RECT 103.0000 47.1000 103.4000 47.2000 ;
	    RECT 105.4000 47.1000 105.8000 47.2000 ;
	    RECT 75.0000 46.8000 105.8000 47.1000 ;
	    RECT 119.8000 46.8000 120.2000 47.2000 ;
	    RECT 127.8000 47.1000 128.2000 47.2000 ;
	    RECT 130.2000 47.1000 130.6000 47.2000 ;
	    RECT 127.8000 46.8000 130.6000 47.1000 ;
	    RECT 199.0000 47.1000 199.4000 47.2000 ;
	    RECT 201.4000 47.1000 201.8000 47.2000 ;
	    RECT 199.0000 46.8000 201.8000 47.1000 ;
	    RECT 212.6000 46.8000 213.0000 47.2000 ;
	    RECT 243.0000 47.1000 243.4000 47.2000 ;
	    RECT 253.4000 47.1000 253.8000 47.2000 ;
	    RECT 243.0000 46.8000 253.8000 47.1000 ;
	    RECT 7.0000 46.1000 7.4000 46.2000 ;
	    RECT 10.2000 46.1000 10.6000 46.2000 ;
	    RECT 7.0000 45.8000 10.6000 46.1000 ;
	    RECT 17.4000 46.1000 17.8000 46.2000 ;
	    RECT 19.8000 46.1000 20.2000 46.2000 ;
	    RECT 17.4000 45.8000 20.2000 46.1000 ;
	    RECT 49.4000 46.1000 49.7000 46.8000 ;
	    RECT 52.6000 46.1000 52.9000 46.8000 ;
	    RECT 49.4000 45.8000 52.9000 46.1000 ;
	    RECT 63.0000 46.1000 63.4000 46.2000 ;
	    RECT 64.6000 46.1000 65.0000 46.2000 ;
	    RECT 69.4000 46.1000 69.8000 46.2000 ;
	    RECT 72.6000 46.1000 73.0000 46.2000 ;
	    RECT 63.0000 45.8000 73.0000 46.1000 ;
	    RECT 75.0000 46.1000 75.4000 46.2000 ;
	    RECT 83.8000 46.1000 84.2000 46.2000 ;
	    RECT 91.8000 46.1000 92.2000 46.2000 ;
	    RECT 75.0000 45.8000 82.5000 46.1000 ;
	    RECT 83.8000 45.8000 92.2000 46.1000 ;
	    RECT 93.4000 46.1000 93.8000 46.2000 ;
	    RECT 111.0000 46.1000 111.4000 46.2000 ;
	    RECT 93.4000 45.8000 111.4000 46.1000 ;
	    RECT 119.8000 46.1000 120.1000 46.8000 ;
	    RECT 126.2000 46.1000 126.6000 46.2000 ;
	    RECT 119.8000 45.8000 126.6000 46.1000 ;
	    RECT 128.6000 46.1000 129.0000 46.2000 ;
	    RECT 131.0000 46.1000 131.4000 46.2000 ;
	    RECT 171.8000 46.1000 172.2000 46.3000 ;
	    RECT 174.2000 46.1000 174.6000 46.2000 ;
	    RECT 201.4000 46.1000 201.7000 46.8000 ;
	    RECT 203.0000 46.1000 203.4000 46.2000 ;
	    RECT 128.6000 45.8000 131.4000 46.1000 ;
	    RECT 133.4000 45.8000 144.1000 46.1000 ;
	    RECT 171.8000 45.8000 174.6000 46.1000 ;
	    RECT 189.4000 45.8000 192.9000 46.1000 ;
	    RECT 201.4000 45.8000 203.4000 46.1000 ;
	    RECT 209.4000 46.1000 209.8000 46.2000 ;
	    RECT 212.6000 46.1000 212.9000 46.8000 ;
	    RECT 248.6000 46.2000 248.9000 46.8000 ;
	    RECT 209.4000 45.8000 212.9000 46.1000 ;
	    RECT 215.0000 46.1000 215.4000 46.2000 ;
	    RECT 225.4000 46.1000 225.8000 46.2000 ;
	    RECT 215.0000 45.8000 242.5000 46.1000 ;
	    RECT 248.6000 45.8000 249.0000 46.2000 ;
	    RECT 82.2000 45.2000 82.5000 45.8000 ;
	    RECT 133.4000 45.2000 133.7000 45.8000 ;
	    RECT 143.8000 45.2000 144.1000 45.8000 ;
	    RECT 189.4000 45.2000 189.7000 45.8000 ;
	    RECT 192.6000 45.2000 192.9000 45.8000 ;
	    RECT 232.6000 45.2000 232.9000 45.8000 ;
	    RECT 242.2000 45.2000 242.5000 45.8000 ;
	    RECT 9.4000 45.1000 9.8000 45.2000 ;
	    RECT 15.0000 45.1000 15.4000 45.2000 ;
	    RECT 9.4000 44.8000 15.4000 45.1000 ;
	    RECT 31.8000 44.8000 32.2000 45.2000 ;
	    RECT 69.4000 45.1000 69.8000 45.2000 ;
	    RECT 75.8000 45.1000 76.2000 45.2000 ;
	    RECT 69.4000 44.8000 76.2000 45.1000 ;
	    RECT 82.2000 44.8000 82.6000 45.2000 ;
	    RECT 87.0000 45.1000 87.4000 45.2000 ;
	    RECT 95.8000 45.1000 96.2000 45.2000 ;
	    RECT 87.0000 44.8000 96.2000 45.1000 ;
	    RECT 105.4000 45.1000 105.8000 45.2000 ;
	    RECT 108.6000 45.1000 109.0000 45.2000 ;
	    RECT 105.4000 44.8000 109.0000 45.1000 ;
	    RECT 111.0000 44.8000 111.4000 45.2000 ;
	    RECT 125.4000 45.1000 125.8000 45.2000 ;
	    RECT 127.8000 45.1000 128.2000 45.2000 ;
	    RECT 125.4000 44.8000 128.2000 45.1000 ;
	    RECT 129.4000 45.1000 129.8000 45.2000 ;
	    RECT 130.2000 45.1000 130.6000 45.2000 ;
	    RECT 129.4000 44.8000 130.6000 45.1000 ;
	    RECT 133.4000 44.8000 133.8000 45.2000 ;
	    RECT 135.0000 44.8000 135.4000 45.2000 ;
	    RECT 143.8000 44.8000 144.2000 45.2000 ;
	    RECT 189.4000 44.8000 189.8000 45.2000 ;
	    RECT 192.6000 44.8000 193.0000 45.2000 ;
	    RECT 232.6000 44.8000 233.0000 45.2000 ;
	    RECT 235.8000 45.1000 236.2000 45.2000 ;
	    RECT 239.0000 45.1000 239.4000 45.2000 ;
	    RECT 235.8000 44.8000 239.4000 45.1000 ;
	    RECT 242.2000 45.1000 242.6000 45.2000 ;
	    RECT 250.2000 45.1000 250.6000 45.2000 ;
	    RECT 242.2000 44.8000 250.6000 45.1000 ;
	    RECT 252.6000 44.8000 253.0000 45.2000 ;
	    RECT 253.4000 45.1000 253.8000 45.2000 ;
	    RECT 255.8000 45.1000 256.2000 45.2000 ;
	    RECT 253.4000 44.8000 256.2000 45.1000 ;
	    RECT 31.8000 44.2000 32.1000 44.8000 ;
	    RECT 111.0000 44.2000 111.3000 44.8000 ;
	    RECT 31.8000 43.8000 32.2000 44.2000 ;
	    RECT 111.0000 43.8000 111.4000 44.2000 ;
	    RECT 121.4000 44.1000 121.8000 44.2000 ;
	    RECT 135.0000 44.1000 135.3000 44.8000 ;
	    RECT 252.6000 44.2000 252.9000 44.8000 ;
	    RECT 121.4000 43.8000 135.3000 44.1000 ;
	    RECT 153.4000 44.1000 153.8000 44.2000 ;
	    RECT 174.2000 44.1000 174.6000 44.2000 ;
	    RECT 153.4000 43.8000 174.6000 44.1000 ;
	    RECT 252.6000 43.8000 253.0000 44.2000 ;
	    RECT 63.8000 43.1000 64.2000 43.2000 ;
	    RECT 67.0000 43.1000 67.4000 43.2000 ;
	    RECT 83.0000 43.1000 83.4000 43.2000 ;
	    RECT 63.8000 42.8000 83.4000 43.1000 ;
	    RECT 105.4000 43.1000 105.8000 43.2000 ;
	    RECT 123.0000 43.1000 123.4000 43.2000 ;
	    RECT 124.6000 43.1000 125.0000 43.2000 ;
	    RECT 105.4000 42.8000 125.0000 43.1000 ;
	    RECT 250.2000 43.1000 250.6000 43.2000 ;
	    RECT 261.4000 43.1000 261.8000 43.2000 ;
	    RECT 250.2000 42.8000 261.8000 43.1000 ;
	    RECT 55.8000 42.1000 56.2000 42.2000 ;
	    RECT 157.4000 42.1000 157.8000 42.2000 ;
	    RECT 163.0000 42.1000 163.4000 42.2000 ;
	    RECT 175.8000 42.1000 176.2000 42.2000 ;
	    RECT 55.8000 41.8000 176.2000 42.1000 ;
	    RECT 259.0000 42.1000 259.4000 42.2000 ;
	    RECT 259.8000 42.1000 260.2000 42.2000 ;
	    RECT 259.0000 41.8000 260.2000 42.1000 ;
	    RECT 82.2000 40.8000 82.6000 41.2000 ;
	    RECT 82.2000 40.2000 82.5000 40.8000 ;
	    RECT 82.2000 39.8000 82.6000 40.2000 ;
	    RECT 255.8000 40.1000 256.2000 40.2000 ;
	    RECT 261.4000 40.1000 261.8000 40.2000 ;
	    RECT 255.8000 39.8000 261.8000 40.1000 ;
	    RECT 56.6000 39.1000 57.0000 39.2000 ;
	    RECT 77.4000 39.1000 77.8000 39.2000 ;
	    RECT 56.6000 38.8000 77.8000 39.1000 ;
	    RECT 104.6000 39.1000 105.0000 39.2000 ;
	    RECT 106.2000 39.1000 106.6000 39.2000 ;
	    RECT 115.0000 39.1000 115.4000 39.2000 ;
	    RECT 123.8000 39.1000 124.2000 39.2000 ;
	    RECT 104.6000 38.8000 124.2000 39.1000 ;
	    RECT 202.2000 39.1000 202.6000 39.2000 ;
	    RECT 217.4000 39.1000 217.8000 39.2000 ;
	    RECT 202.2000 38.8000 217.8000 39.1000 ;
	    RECT 231.8000 39.1000 232.2000 39.2000 ;
	    RECT 233.4000 39.1000 233.8000 39.2000 ;
	    RECT 231.8000 38.8000 233.8000 39.1000 ;
	    RECT 83.0000 38.1000 83.4000 38.2000 ;
	    RECT 86.2000 38.1000 86.6000 38.2000 ;
	    RECT 111.0000 38.1000 111.4000 38.2000 ;
	    RECT 83.0000 37.8000 111.4000 38.1000 ;
	    RECT 119.0000 38.1000 119.4000 38.2000 ;
	    RECT 119.8000 38.1000 120.2000 38.2000 ;
	    RECT 119.0000 37.8000 120.2000 38.1000 ;
	    RECT 254.2000 38.1000 254.6000 38.2000 ;
	    RECT 259.0000 38.1000 259.4000 38.2000 ;
	    RECT 254.2000 37.8000 259.4000 38.1000 ;
	    RECT 3.0000 37.1000 3.4000 37.2000 ;
	    RECT 27.8000 37.1000 28.2000 37.2000 ;
	    RECT 3.0000 36.8000 28.2000 37.1000 ;
	    RECT 78.2000 37.1000 78.6000 37.2000 ;
	    RECT 98.2000 37.1000 98.6000 37.2000 ;
	    RECT 145.4000 37.1000 145.8000 37.2000 ;
	    RECT 78.2000 36.8000 98.6000 37.1000 ;
	    RECT 139.0000 36.8000 145.8000 37.1000 ;
	    RECT 164.6000 37.1000 165.0000 37.2000 ;
	    RECT 197.4000 37.1000 197.8000 37.2000 ;
	    RECT 164.6000 36.8000 197.8000 37.1000 ;
	    RECT 233.4000 37.1000 233.8000 37.2000 ;
	    RECT 239.8000 37.1000 240.2000 37.2000 ;
	    RECT 233.4000 36.8000 240.2000 37.1000 ;
	    RECT 139.0000 36.2000 139.3000 36.8000 ;
	    RECT 19.8000 36.1000 20.2000 36.2000 ;
	    RECT 27.0000 36.1000 27.4000 36.2000 ;
	    RECT 19.8000 35.8000 27.4000 36.1000 ;
	    RECT 30.2000 36.1000 30.6000 36.2000 ;
	    RECT 37.4000 36.1000 37.8000 36.2000 ;
	    RECT 30.2000 35.8000 37.8000 36.1000 ;
	    RECT 49.4000 36.1000 49.8000 36.2000 ;
	    RECT 55.8000 36.1000 56.2000 36.2000 ;
	    RECT 49.4000 35.8000 56.2000 36.1000 ;
	    RECT 62.2000 36.1000 62.6000 36.2000 ;
	    RECT 66.2000 36.1000 66.6000 36.2000 ;
	    RECT 62.2000 35.8000 66.6000 36.1000 ;
	    RECT 85.4000 35.8000 85.8000 36.2000 ;
	    RECT 106.2000 36.1000 106.6000 36.2000 ;
	    RECT 120.6000 36.1000 121.0000 36.2000 ;
	    RECT 106.2000 35.8000 121.0000 36.1000 ;
	    RECT 123.0000 36.1000 123.4000 36.2000 ;
	    RECT 124.6000 36.1000 125.0000 36.2000 ;
	    RECT 129.4000 36.1000 129.8000 36.2000 ;
	    RECT 123.0000 35.8000 129.8000 36.1000 ;
	    RECT 139.0000 35.8000 139.4000 36.2000 ;
	    RECT 139.8000 35.8000 140.2000 36.2000 ;
	    RECT 140.6000 36.1000 141.0000 36.2000 ;
	    RECT 157.4000 36.1000 157.8000 36.2000 ;
	    RECT 173.4000 36.1000 173.8000 36.2000 ;
	    RECT 140.6000 35.8000 173.8000 36.1000 ;
	    RECT 181.4000 35.8000 181.8000 36.2000 ;
	    RECT 187.8000 36.1000 188.2000 36.2000 ;
	    RECT 189.4000 36.1000 189.8000 36.2000 ;
	    RECT 191.8000 36.1000 192.2000 36.2000 ;
	    RECT 187.8000 35.8000 192.2000 36.1000 ;
	    RECT 204.6000 36.1000 205.0000 36.2000 ;
	    RECT 206.2000 36.1000 206.6000 36.2000 ;
	    RECT 204.6000 35.8000 206.6000 36.1000 ;
	    RECT 211.8000 35.8000 212.2000 36.2000 ;
	    RECT 229.4000 36.1000 229.8000 36.2000 ;
	    RECT 246.2000 36.1000 246.6000 36.2000 ;
	    RECT 254.2000 36.1000 254.6000 36.2000 ;
	    RECT 258.2000 36.1000 258.6000 36.2000 ;
	    RECT 229.4000 35.8000 258.6000 36.1000 ;
	    RECT 261.4000 36.1000 261.8000 36.2000 ;
	    RECT 267.8000 36.1000 268.2000 36.2000 ;
	    RECT 261.4000 35.8000 268.2000 36.1000 ;
	    RECT 12.6000 35.1000 13.0000 35.2000 ;
	    RECT 15.0000 35.1000 15.4000 35.2000 ;
	    RECT 12.6000 34.8000 15.4000 35.1000 ;
	    RECT 15.8000 35.1000 16.2000 35.2000 ;
	    RECT 18.2000 35.1000 18.6000 35.2000 ;
	    RECT 15.8000 34.8000 18.6000 35.1000 ;
	    RECT 27.0000 35.1000 27.4000 35.2000 ;
	    RECT 32.6000 35.1000 33.0000 35.2000 ;
	    RECT 27.0000 34.8000 33.0000 35.1000 ;
	    RECT 45.4000 35.1000 45.8000 35.2000 ;
	    RECT 47.0000 35.1000 47.4000 35.2000 ;
	    RECT 45.4000 34.8000 47.4000 35.1000 ;
	    RECT 50.2000 35.1000 50.6000 35.2000 ;
	    RECT 63.8000 35.1000 64.2000 35.2000 ;
	    RECT 70.2000 35.1000 70.6000 35.2000 ;
	    RECT 76.6000 35.1000 77.0000 35.2000 ;
	    RECT 50.2000 34.8000 77.0000 35.1000 ;
	    RECT 82.2000 35.1000 82.6000 35.2000 ;
	    RECT 85.4000 35.1000 85.7000 35.8000 ;
	    RECT 82.2000 34.8000 85.7000 35.1000 ;
	    RECT 95.0000 35.1000 95.4000 35.2000 ;
	    RECT 99.0000 35.1000 99.4000 35.2000 ;
	    RECT 95.0000 34.8000 99.4000 35.1000 ;
	    RECT 101.4000 35.1000 101.8000 35.2000 ;
	    RECT 119.0000 35.1000 119.4000 35.2000 ;
	    RECT 122.2000 35.1000 122.6000 35.2000 ;
	    RECT 138.2000 35.1000 138.6000 35.2000 ;
	    RECT 139.8000 35.1000 140.1000 35.8000 ;
	    RECT 181.4000 35.2000 181.7000 35.8000 ;
	    RECT 101.4000 34.8000 119.4000 35.1000 ;
	    RECT 121.4000 34.8000 129.7000 35.1000 ;
	    RECT 138.2000 34.8000 140.1000 35.1000 ;
	    RECT 155.8000 35.1000 156.2000 35.2000 ;
	    RECT 159.0000 35.1000 159.4000 35.2000 ;
	    RECT 171.8000 35.1000 172.2000 35.2000 ;
	    RECT 155.8000 34.8000 164.1000 35.1000 ;
	    RECT 31.0000 34.2000 31.3000 34.8000 ;
	    RECT 129.4000 34.2000 129.7000 34.8000 ;
	    RECT 163.8000 34.2000 164.1000 34.8000 ;
	    RECT 167.0000 34.8000 172.2000 35.1000 ;
	    RECT 174.2000 35.1000 174.6000 35.2000 ;
	    RECT 177.4000 35.1000 177.8000 35.2000 ;
	    RECT 174.2000 34.8000 177.8000 35.1000 ;
	    RECT 179.8000 34.8000 180.2000 35.2000 ;
	    RECT 181.4000 34.8000 181.8000 35.2000 ;
	    RECT 203.8000 35.1000 204.2000 35.2000 ;
	    RECT 206.2000 35.1000 206.6000 35.2000 ;
	    RECT 191.0000 34.8000 206.6000 35.1000 ;
	    RECT 208.6000 35.1000 209.0000 35.2000 ;
	    RECT 211.8000 35.1000 212.1000 35.8000 ;
	    RECT 208.6000 34.8000 212.1000 35.1000 ;
	    RECT 224.6000 34.8000 225.0000 35.2000 ;
	    RECT 234.2000 35.1000 234.6000 35.2000 ;
	    RECT 246.2000 35.1000 246.6000 35.2000 ;
	    RECT 247.0000 35.1000 247.4000 35.2000 ;
	    RECT 262.2000 35.1000 262.6000 35.2000 ;
	    RECT 234.2000 34.8000 262.6000 35.1000 ;
	    RECT 167.0000 34.2000 167.3000 34.8000 ;
	    RECT 14.2000 34.1000 14.6000 34.2000 ;
	    RECT 15.0000 34.1000 15.4000 34.2000 ;
	    RECT 14.2000 33.8000 15.4000 34.1000 ;
	    RECT 16.6000 34.1000 17.0000 34.2000 ;
	    RECT 19.8000 34.1000 20.2000 34.2000 ;
	    RECT 16.6000 33.8000 20.2000 34.1000 ;
	    RECT 23.8000 34.1000 24.2000 34.2000 ;
	    RECT 24.6000 34.1000 25.0000 34.2000 ;
	    RECT 23.8000 33.8000 25.0000 34.1000 ;
	    RECT 31.0000 33.8000 31.4000 34.2000 ;
	    RECT 41.4000 34.1000 41.8000 34.2000 ;
	    RECT 44.6000 34.1000 45.0000 34.2000 ;
	    RECT 41.4000 33.8000 45.0000 34.1000 ;
	    RECT 99.0000 33.8000 99.4000 34.2000 ;
	    RECT 119.0000 34.1000 119.4000 34.2000 ;
	    RECT 121.4000 34.1000 121.8000 34.2000 ;
	    RECT 119.0000 33.8000 121.8000 34.1000 ;
	    RECT 123.8000 34.1000 124.2000 34.2000 ;
	    RECT 124.6000 34.1000 125.0000 34.2000 ;
	    RECT 123.8000 33.8000 125.0000 34.1000 ;
	    RECT 129.4000 33.8000 129.8000 34.2000 ;
	    RECT 134.2000 34.1000 134.6000 34.2000 ;
	    RECT 140.6000 34.1000 141.0000 34.2000 ;
	    RECT 151.8000 34.1000 152.2000 34.2000 ;
	    RECT 154.2000 34.1000 154.6000 34.2000 ;
	    RECT 134.2000 33.8000 154.6000 34.1000 ;
	    RECT 163.8000 33.8000 164.2000 34.2000 ;
	    RECT 167.0000 33.8000 167.4000 34.2000 ;
	    RECT 168.6000 34.1000 169.0000 34.2000 ;
	    RECT 179.8000 34.1000 180.1000 34.8000 ;
	    RECT 168.6000 33.8000 180.1000 34.1000 ;
	    RECT 188.6000 34.1000 189.0000 34.2000 ;
	    RECT 191.0000 34.1000 191.3000 34.8000 ;
	    RECT 224.6000 34.2000 224.9000 34.8000 ;
	    RECT 191.8000 34.1000 192.2000 34.2000 ;
	    RECT 188.6000 33.8000 192.2000 34.1000 ;
	    RECT 200.6000 34.1000 201.0000 34.2000 ;
	    RECT 220.6000 34.1000 221.0000 34.2000 ;
	    RECT 200.6000 33.8000 210.5000 34.1000 ;
	    RECT 99.0000 33.2000 99.3000 33.8000 ;
	    RECT 210.2000 33.2000 210.5000 33.8000 ;
	    RECT 219.0000 33.8000 221.0000 34.1000 ;
	    RECT 224.6000 33.8000 225.0000 34.2000 ;
	    RECT 231.8000 34.1000 232.2000 34.2000 ;
	    RECT 231.8000 33.8000 236.1000 34.1000 ;
	    RECT 219.0000 33.2000 219.3000 33.8000 ;
	    RECT 235.8000 33.2000 236.1000 33.8000 ;
	    RECT 242.2000 33.8000 242.6000 34.2000 ;
	    RECT 246.2000 34.1000 246.6000 34.2000 ;
	    RECT 255.8000 34.1000 256.2000 34.2000 ;
	    RECT 246.2000 33.8000 256.2000 34.1000 ;
	    RECT 260.6000 34.1000 261.0000 34.2000 ;
	    RECT 263.0000 34.1000 263.4000 34.2000 ;
	    RECT 260.6000 33.8000 263.4000 34.1000 ;
	    RECT 242.2000 33.2000 242.5000 33.8000 ;
	    RECT 18.2000 33.1000 18.6000 33.2000 ;
	    RECT 93.4000 33.1000 93.8000 33.2000 ;
	    RECT 97.4000 33.1000 97.8000 33.2000 ;
	    RECT 18.2000 32.8000 24.1000 33.1000 ;
	    RECT 93.4000 32.8000 97.8000 33.1000 ;
	    RECT 99.0000 32.8000 99.4000 33.2000 ;
	    RECT 103.8000 33.1000 104.2000 33.2000 ;
	    RECT 116.6000 33.1000 117.0000 33.2000 ;
	    RECT 103.8000 32.8000 117.0000 33.1000 ;
	    RECT 122.2000 33.1000 122.6000 33.2000 ;
	    RECT 136.6000 33.1000 137.0000 33.2000 ;
	    RECT 122.2000 32.8000 137.0000 33.1000 ;
	    RECT 139.0000 33.1000 139.4000 33.2000 ;
	    RECT 141.4000 33.1000 141.8000 33.2000 ;
	    RECT 142.2000 33.1000 142.6000 33.2000 ;
	    RECT 139.0000 32.8000 142.6000 33.1000 ;
	    RECT 176.6000 33.1000 177.0000 33.2000 ;
	    RECT 177.4000 33.1000 177.8000 33.2000 ;
	    RECT 176.6000 32.8000 177.8000 33.1000 ;
	    RECT 191.8000 33.1000 192.2000 33.2000 ;
	    RECT 193.4000 33.1000 193.8000 33.2000 ;
	    RECT 191.8000 32.8000 193.8000 33.1000 ;
	    RECT 210.2000 32.8000 210.6000 33.2000 ;
	    RECT 219.0000 32.8000 219.4000 33.2000 ;
	    RECT 223.0000 33.1000 223.4000 33.2000 ;
	    RECT 231.0000 33.1000 231.4000 33.2000 ;
	    RECT 223.0000 32.8000 231.4000 33.1000 ;
	    RECT 235.8000 32.8000 236.2000 33.2000 ;
	    RECT 242.2000 32.8000 242.6000 33.2000 ;
	    RECT 243.8000 33.1000 244.2000 33.2000 ;
	    RECT 244.6000 33.1000 245.0000 33.2000 ;
	    RECT 243.8000 32.8000 245.0000 33.1000 ;
	    RECT 23.8000 32.2000 24.1000 32.8000 ;
	    RECT 23.8000 31.8000 24.2000 32.2000 ;
	    RECT 72.6000 32.1000 73.0000 32.2000 ;
	    RECT 76.6000 32.1000 77.0000 32.2000 ;
	    RECT 95.0000 32.1000 95.4000 32.2000 ;
	    RECT 72.6000 31.8000 95.4000 32.1000 ;
	    RECT 99.0000 32.1000 99.4000 32.2000 ;
	    RECT 102.2000 32.1000 102.6000 32.2000 ;
	    RECT 99.0000 31.8000 102.6000 32.1000 ;
	    RECT 103.8000 32.1000 104.2000 32.2000 ;
	    RECT 110.2000 32.1000 110.6000 32.2000 ;
	    RECT 103.8000 31.8000 110.6000 32.1000 ;
	    RECT 127.8000 32.1000 128.2000 32.2000 ;
	    RECT 156.6000 32.1000 157.0000 32.2000 ;
	    RECT 127.8000 31.8000 157.0000 32.1000 ;
	    RECT 161.4000 32.1000 161.8000 32.2000 ;
	    RECT 170.2000 32.1000 170.6000 32.2000 ;
	    RECT 161.4000 31.8000 170.6000 32.1000 ;
	    RECT 205.4000 32.1000 205.8000 32.2000 ;
	    RECT 224.6000 32.1000 225.0000 32.2000 ;
	    RECT 205.4000 31.8000 225.0000 32.1000 ;
	    RECT 225.4000 32.1000 225.8000 32.2000 ;
	    RECT 242.2000 32.1000 242.6000 32.2000 ;
	    RECT 225.4000 31.8000 242.6000 32.1000 ;
	    RECT 259.8000 32.1000 260.2000 32.2000 ;
	    RECT 263.8000 32.1000 264.2000 32.2000 ;
	    RECT 265.4000 32.1000 265.8000 32.2000 ;
	    RECT 259.8000 31.8000 265.8000 32.1000 ;
	    RECT 91.0000 31.1000 91.4000 31.2000 ;
	    RECT 98.2000 31.1000 98.6000 31.2000 ;
	    RECT 105.4000 31.1000 105.8000 31.2000 ;
	    RECT 91.0000 30.8000 105.8000 31.1000 ;
	    RECT 125.4000 31.1000 125.8000 31.2000 ;
	    RECT 131.8000 31.1000 132.2000 31.2000 ;
	    RECT 135.8000 31.1000 136.2000 31.2000 ;
	    RECT 152.6000 31.1000 153.0000 31.2000 ;
	    RECT 125.4000 30.8000 153.0000 31.1000 ;
	    RECT 185.4000 31.1000 185.8000 31.2000 ;
	    RECT 186.2000 31.1000 186.6000 31.2000 ;
	    RECT 185.4000 30.8000 186.6000 31.1000 ;
	    RECT 215.8000 31.1000 216.2000 31.2000 ;
	    RECT 219.8000 31.1000 220.2000 31.2000 ;
	    RECT 215.8000 30.8000 220.2000 31.1000 ;
	    RECT 220.6000 31.1000 221.0000 31.2000 ;
	    RECT 236.6000 31.1000 237.0000 31.2000 ;
	    RECT 220.6000 30.8000 237.0000 31.1000 ;
	    RECT 237.4000 31.1000 237.8000 31.2000 ;
	    RECT 256.6000 31.1000 257.0000 31.2000 ;
	    RECT 237.4000 30.8000 257.0000 31.1000 ;
	    RECT 8.6000 30.1000 9.0000 30.2000 ;
	    RECT 20.6000 30.1000 21.0000 30.2000 ;
	    RECT 8.6000 29.8000 21.0000 30.1000 ;
	    RECT 130.2000 30.1000 130.6000 30.2000 ;
	    RECT 132.6000 30.1000 133.0000 30.2000 ;
	    RECT 145.4000 30.1000 145.8000 30.2000 ;
	    RECT 130.2000 29.8000 145.8000 30.1000 ;
	    RECT 163.0000 30.1000 163.4000 30.2000 ;
	    RECT 166.2000 30.1000 166.6000 30.2000 ;
	    RECT 175.0000 30.1000 175.4000 30.2000 ;
	    RECT 178.2000 30.1000 178.6000 30.2000 ;
	    RECT 163.0000 29.8000 178.6000 30.1000 ;
	    RECT 238.2000 29.8000 238.6000 30.2000 ;
	    RECT 240.6000 30.1000 241.0000 30.2000 ;
	    RECT 243.0000 30.1000 243.4000 30.2000 ;
	    RECT 240.6000 29.8000 243.4000 30.1000 ;
	    RECT 251.8000 30.1000 252.2000 30.2000 ;
	    RECT 259.0000 30.1000 259.4000 30.2000 ;
	    RECT 251.8000 29.8000 259.4000 30.1000 ;
	    RECT 238.2000 29.2000 238.5000 29.8000 ;
	    RECT 15.0000 28.8000 15.4000 29.2000 ;
	    RECT 20.6000 29.1000 21.0000 29.2000 ;
	    RECT 22.2000 29.1000 22.6000 29.2000 ;
	    RECT 20.6000 28.8000 22.6000 29.1000 ;
	    RECT 67.8000 29.1000 68.2000 29.2000 ;
	    RECT 72.6000 29.1000 73.0000 29.2000 ;
	    RECT 67.8000 28.8000 73.0000 29.1000 ;
	    RECT 83.8000 29.1000 84.2000 29.2000 ;
	    RECT 84.6000 29.1000 85.0000 29.2000 ;
	    RECT 83.8000 28.8000 85.0000 29.1000 ;
	    RECT 101.4000 29.1000 101.8000 29.2000 ;
	    RECT 117.4000 29.1000 117.8000 29.2000 ;
	    RECT 101.4000 28.8000 117.8000 29.1000 ;
	    RECT 121.4000 29.1000 121.8000 29.2000 ;
	    RECT 122.2000 29.1000 122.6000 29.2000 ;
	    RECT 121.4000 28.8000 122.6000 29.1000 ;
	    RECT 126.2000 29.1000 126.6000 29.2000 ;
	    RECT 129.4000 29.1000 129.8000 29.2000 ;
	    RECT 126.2000 28.8000 129.8000 29.1000 ;
	    RECT 131.0000 29.1000 131.4000 29.2000 ;
	    RECT 133.4000 29.1000 133.8000 29.2000 ;
	    RECT 131.0000 28.8000 133.8000 29.1000 ;
	    RECT 153.4000 29.1000 153.8000 29.2000 ;
	    RECT 204.6000 29.1000 205.0000 29.2000 ;
	    RECT 233.4000 29.1000 233.8000 29.2000 ;
	    RECT 153.4000 28.8000 168.1000 29.1000 ;
	    RECT 204.6000 28.8000 233.8000 29.1000 ;
	    RECT 238.2000 28.8000 238.6000 29.2000 ;
	    RECT 239.0000 29.1000 239.4000 29.2000 ;
	    RECT 244.6000 29.1000 245.0000 29.2000 ;
	    RECT 239.0000 28.8000 245.0000 29.1000 ;
	    RECT 254.2000 29.1000 254.6000 29.2000 ;
	    RECT 257.4000 29.1000 257.8000 29.2000 ;
	    RECT 254.2000 28.8000 257.8000 29.1000 ;
	    RECT 15.0000 28.1000 15.3000 28.8000 ;
	    RECT 167.8000 28.2000 168.1000 28.8000 ;
	    RECT 18.2000 28.1000 18.6000 28.2000 ;
	    RECT 15.0000 27.8000 18.6000 28.1000 ;
	    RECT 21.4000 28.1000 21.8000 28.2000 ;
	    RECT 22.2000 28.1000 22.6000 28.2000 ;
	    RECT 21.4000 27.8000 22.6000 28.1000 ;
	    RECT 66.2000 28.1000 66.6000 28.2000 ;
	    RECT 68.6000 28.1000 69.0000 28.2000 ;
	    RECT 92.6000 28.1000 93.0000 28.2000 ;
	    RECT 66.2000 27.8000 93.0000 28.1000 ;
	    RECT 97.4000 28.1000 97.8000 28.2000 ;
	    RECT 104.6000 28.1000 105.0000 28.2000 ;
	    RECT 107.8000 28.1000 108.2000 28.2000 ;
	    RECT 97.4000 27.8000 108.2000 28.1000 ;
	    RECT 108.6000 28.1000 109.0000 28.2000 ;
	    RECT 111.0000 28.1000 111.4000 28.2000 ;
	    RECT 108.6000 27.8000 111.4000 28.1000 ;
	    RECT 119.0000 28.1000 119.4000 28.2000 ;
	    RECT 123.0000 28.1000 123.4000 28.2000 ;
	    RECT 139.0000 28.1000 139.4000 28.2000 ;
	    RECT 119.0000 27.8000 139.4000 28.1000 ;
	    RECT 149.4000 27.8000 149.8000 28.2000 ;
	    RECT 151.0000 28.1000 151.4000 28.2000 ;
	    RECT 157.4000 28.1000 157.8000 28.2000 ;
	    RECT 165.4000 28.1000 165.8000 28.2000 ;
	    RECT 151.0000 27.8000 165.8000 28.1000 ;
	    RECT 167.8000 27.8000 168.2000 28.2000 ;
	    RECT 182.2000 28.1000 182.6000 28.2000 ;
	    RECT 194.2000 28.1000 194.6000 28.2000 ;
	    RECT 182.2000 27.8000 194.6000 28.1000 ;
	    RECT 207.8000 28.1000 208.2000 28.2000 ;
	    RECT 210.2000 28.1000 210.6000 28.2000 ;
	    RECT 207.8000 27.8000 210.6000 28.1000 ;
	    RECT 217.4000 27.8000 217.8000 28.2000 ;
	    RECT 229.4000 28.1000 229.8000 28.2000 ;
	    RECT 231.0000 28.1000 231.4000 28.2000 ;
	    RECT 228.6000 27.8000 231.4000 28.1000 ;
	    RECT 232.6000 28.1000 233.0000 28.2000 ;
	    RECT 237.4000 28.1000 237.8000 28.2000 ;
	    RECT 232.6000 27.8000 237.8000 28.1000 ;
	    RECT 248.6000 28.1000 249.0000 28.2000 ;
	    RECT 254.2000 28.1000 254.6000 28.2000 ;
	    RECT 248.6000 27.8000 254.6000 28.1000 ;
	    RECT 257.4000 28.1000 257.8000 28.2000 ;
	    RECT 266.2000 28.1000 266.6000 28.2000 ;
	    RECT 257.4000 27.8000 266.6000 28.1000 ;
	    RECT 3.8000 27.1000 4.2000 27.2000 ;
	    RECT 7.0000 27.1000 7.4000 27.2000 ;
	    RECT 3.8000 26.8000 7.4000 27.1000 ;
	    RECT 9.4000 27.1000 9.8000 27.2000 ;
	    RECT 16.6000 27.1000 17.0000 27.2000 ;
	    RECT 9.4000 26.8000 17.0000 27.1000 ;
	    RECT 25.4000 27.1000 25.8000 27.2000 ;
	    RECT 29.4000 27.1000 29.8000 27.2000 ;
	    RECT 25.4000 26.8000 29.8000 27.1000 ;
	    RECT 36.6000 27.1000 37.0000 27.2000 ;
	    RECT 43.8000 27.1000 44.2000 27.2000 ;
	    RECT 36.6000 26.8000 44.2000 27.1000 ;
	    RECT 60.6000 26.8000 61.0000 27.2000 ;
	    RECT 65.4000 27.1000 65.8000 27.2000 ;
	    RECT 99.8000 27.1000 100.2000 27.2000 ;
	    RECT 65.4000 26.8000 100.2000 27.1000 ;
	    RECT 105.4000 27.1000 105.8000 27.2000 ;
	    RECT 111.0000 27.1000 111.4000 27.2000 ;
	    RECT 105.4000 26.8000 111.4000 27.1000 ;
	    RECT 131.8000 27.1000 132.2000 27.2000 ;
	    RECT 135.0000 27.1000 135.4000 27.2000 ;
	    RECT 140.6000 27.1000 141.0000 27.2000 ;
	    RECT 131.8000 26.8000 141.0000 27.1000 ;
	    RECT 149.4000 27.1000 149.7000 27.8000 ;
	    RECT 152.6000 27.1000 153.0000 27.2000 ;
	    RECT 171.8000 27.1000 172.2000 27.2000 ;
	    RECT 190.2000 27.1000 190.6000 27.2000 ;
	    RECT 149.4000 26.8000 153.7000 27.1000 ;
	    RECT 171.8000 26.8000 190.6000 27.1000 ;
	    RECT 192.6000 27.1000 193.0000 27.2000 ;
	    RECT 201.4000 27.1000 201.8000 27.2000 ;
	    RECT 192.6000 26.8000 201.8000 27.1000 ;
	    RECT 208.6000 27.1000 209.0000 27.2000 ;
	    RECT 217.4000 27.1000 217.7000 27.8000 ;
	    RECT 208.6000 26.8000 217.7000 27.1000 ;
	    RECT 219.8000 27.1000 220.2000 27.2000 ;
	    RECT 227.0000 27.1000 227.4000 27.2000 ;
	    RECT 229.4000 27.1000 229.8000 27.2000 ;
	    RECT 219.8000 26.8000 229.8000 27.1000 ;
	    RECT 237.4000 26.8000 237.8000 27.2000 ;
	    RECT 243.0000 27.1000 243.4000 27.2000 ;
	    RECT 248.6000 27.1000 248.9000 27.8000 ;
	    RECT 243.0000 26.8000 248.9000 27.1000 ;
	    RECT 255.0000 27.1000 255.4000 27.2000 ;
	    RECT 255.0000 26.8000 261.7000 27.1000 ;
	    RECT 6.2000 26.1000 6.6000 26.2000 ;
	    RECT 11.0000 26.1000 11.4000 26.2000 ;
	    RECT 11.8000 26.1000 12.2000 26.2000 ;
	    RECT 6.2000 25.8000 12.2000 26.1000 ;
	    RECT 27.8000 26.1000 28.2000 26.2000 ;
	    RECT 31.0000 26.1000 31.4000 26.2000 ;
	    RECT 27.8000 25.8000 31.4000 26.1000 ;
	    RECT 43.8000 26.1000 44.2000 26.2000 ;
	    RECT 47.0000 26.1000 47.4000 26.2000 ;
	    RECT 51.8000 26.1000 52.2000 26.2000 ;
	    RECT 43.8000 25.8000 45.7000 26.1000 ;
	    RECT 47.0000 25.8000 52.2000 26.1000 ;
	    RECT 54.2000 26.1000 54.6000 26.2000 ;
	    RECT 60.6000 26.1000 60.9000 26.8000 ;
	    RECT 237.4000 26.2000 237.7000 26.8000 ;
	    RECT 261.4000 26.2000 261.7000 26.8000 ;
	    RECT 263.8000 26.8000 264.2000 27.2000 ;
	    RECT 263.8000 26.2000 264.1000 26.8000 ;
	    RECT 54.2000 25.8000 60.9000 26.1000 ;
	    RECT 70.2000 26.1000 70.6000 26.2000 ;
	    RECT 71.0000 26.1000 71.4000 26.2000 ;
	    RECT 95.0000 26.1000 95.4000 26.2000 ;
	    RECT 107.0000 26.1000 107.4000 26.2000 ;
	    RECT 125.4000 26.1000 125.8000 26.2000 ;
	    RECT 70.2000 25.8000 125.8000 26.1000 ;
	    RECT 127.8000 26.1000 128.2000 26.2000 ;
	    RECT 128.6000 26.1000 129.0000 26.2000 ;
	    RECT 127.8000 25.8000 129.0000 26.1000 ;
	    RECT 136.6000 26.1000 137.0000 26.2000 ;
	    RECT 151.8000 26.1000 152.2000 26.2000 ;
	    RECT 200.6000 26.1000 201.0000 26.2000 ;
	    RECT 221.4000 26.1000 221.8000 26.2000 ;
	    RECT 226.2000 26.1000 226.6000 26.2000 ;
	    RECT 227.8000 26.1000 228.2000 26.2000 ;
	    RECT 136.6000 25.8000 152.2000 26.1000 ;
	    RECT 153.4000 25.8000 156.9000 26.1000 ;
	    RECT 200.6000 25.8000 228.2000 26.1000 ;
	    RECT 237.4000 25.8000 237.8000 26.2000 ;
	    RECT 243.8000 26.1000 244.2000 26.2000 ;
	    RECT 246.2000 26.1000 246.6000 26.2000 ;
	    RECT 243.8000 25.8000 246.6000 26.1000 ;
	    RECT 248.6000 25.8000 252.1000 26.1000 ;
	    RECT 261.4000 25.8000 261.8000 26.2000 ;
	    RECT 263.8000 25.8000 264.2000 26.2000 ;
	    RECT 45.4000 25.2000 45.7000 25.8000 ;
	    RECT 153.4000 25.2000 153.7000 25.8000 ;
	    RECT 156.6000 25.2000 156.9000 25.8000 ;
	    RECT 248.6000 25.2000 248.9000 25.8000 ;
	    RECT 251.8000 25.2000 252.1000 25.8000 ;
	    RECT 17.4000 25.1000 17.8000 25.2000 ;
	    RECT 19.8000 25.1000 20.2000 25.2000 ;
	    RECT 17.4000 24.8000 20.2000 25.1000 ;
	    RECT 24.6000 25.1000 25.0000 25.2000 ;
	    RECT 29.4000 25.1000 29.8000 25.2000 ;
	    RECT 24.6000 24.8000 29.8000 25.1000 ;
	    RECT 45.4000 24.8000 45.8000 25.2000 ;
	    RECT 75.8000 25.1000 76.2000 25.2000 ;
	    RECT 71.8000 24.8000 76.2000 25.1000 ;
	    RECT 78.2000 25.1000 78.6000 25.2000 ;
	    RECT 86.2000 25.1000 86.6000 25.2000 ;
	    RECT 78.2000 24.8000 86.6000 25.1000 ;
	    RECT 89.4000 25.1000 89.8000 25.2000 ;
	    RECT 94.2000 25.1000 94.6000 25.2000 ;
	    RECT 101.4000 25.1000 101.8000 25.2000 ;
	    RECT 89.4000 24.8000 93.7000 25.1000 ;
	    RECT 94.2000 24.8000 101.8000 25.1000 ;
	    RECT 106.2000 25.1000 106.6000 25.2000 ;
	    RECT 110.2000 25.1000 110.6000 25.2000 ;
	    RECT 115.0000 25.1000 115.4000 25.2000 ;
	    RECT 106.2000 24.8000 110.6000 25.1000 ;
	    RECT 111.8000 24.8000 115.4000 25.1000 ;
	    RECT 118.2000 25.1000 118.6000 25.2000 ;
	    RECT 130.2000 25.1000 130.6000 25.2000 ;
	    RECT 118.2000 24.8000 130.6000 25.1000 ;
	    RECT 135.8000 25.1000 136.2000 25.2000 ;
	    RECT 136.6000 25.1000 137.0000 25.2000 ;
	    RECT 147.0000 25.1000 147.4000 25.2000 ;
	    RECT 135.8000 24.8000 137.0000 25.1000 ;
	    RECT 138.2000 24.8000 147.4000 25.1000 ;
	    RECT 153.4000 24.8000 153.8000 25.2000 ;
	    RECT 156.6000 24.8000 157.0000 25.2000 ;
	    RECT 167.0000 25.1000 167.4000 25.2000 ;
	    RECT 181.4000 25.1000 181.8000 25.2000 ;
	    RECT 167.0000 24.8000 181.8000 25.1000 ;
	    RECT 209.4000 25.1000 209.8000 25.2000 ;
	    RECT 211.8000 25.1000 212.2000 25.2000 ;
	    RECT 237.4000 25.1000 237.8000 25.2000 ;
	    RECT 238.2000 25.1000 238.6000 25.2000 ;
	    RECT 209.4000 24.8000 212.2000 25.1000 ;
	    RECT 236.6000 24.8000 238.6000 25.1000 ;
	    RECT 248.6000 24.8000 249.0000 25.2000 ;
	    RECT 251.8000 24.8000 252.2000 25.2000 ;
	    RECT 71.8000 24.2000 72.1000 24.8000 ;
	    RECT 93.4000 24.2000 93.7000 24.8000 ;
	    RECT 111.8000 24.2000 112.1000 24.8000 ;
	    RECT 138.2000 24.2000 138.5000 24.8000 ;
	    RECT 55.8000 24.1000 56.2000 24.2000 ;
	    RECT 66.2000 24.1000 66.6000 24.2000 ;
	    RECT 55.8000 23.8000 66.6000 24.1000 ;
	    RECT 71.8000 23.8000 72.2000 24.2000 ;
	    RECT 93.4000 23.8000 93.8000 24.2000 ;
	    RECT 111.8000 23.8000 112.2000 24.2000 ;
	    RECT 138.2000 23.8000 138.6000 24.2000 ;
	    RECT 179.0000 24.1000 179.4000 24.2000 ;
	    RECT 207.0000 24.1000 207.4000 24.2000 ;
	    RECT 179.0000 23.8000 207.4000 24.1000 ;
	    RECT 214.2000 24.1000 214.6000 24.2000 ;
	    RECT 216.6000 24.1000 217.0000 24.2000 ;
	    RECT 242.2000 24.1000 242.6000 24.2000 ;
	    RECT 243.0000 24.1000 243.4000 24.2000 ;
	    RECT 214.2000 23.8000 243.4000 24.1000 ;
	    RECT 243.8000 24.1000 244.2000 24.2000 ;
	    RECT 244.6000 24.1000 245.0000 24.2000 ;
	    RECT 243.8000 23.8000 245.0000 24.1000 ;
	    RECT 35.8000 23.1000 36.2000 23.2000 ;
	    RECT 39.0000 23.1000 39.4000 23.2000 ;
	    RECT 48.6000 23.1000 49.0000 23.2000 ;
	    RECT 63.8000 23.1000 64.2000 23.2000 ;
	    RECT 78.2000 23.1000 78.6000 23.2000 ;
	    RECT 35.8000 22.8000 78.6000 23.1000 ;
	    RECT 91.8000 23.1000 92.2000 23.2000 ;
	    RECT 98.2000 23.1000 98.6000 23.2000 ;
	    RECT 91.8000 22.8000 98.6000 23.1000 ;
	    RECT 211.0000 23.1000 211.4000 23.2000 ;
	    RECT 234.2000 23.1000 234.6000 23.2000 ;
	    RECT 211.0000 22.8000 234.6000 23.1000 ;
	    RECT 46.2000 22.1000 46.6000 22.2000 ;
	    RECT 51.0000 22.1000 51.4000 22.2000 ;
	    RECT 68.6000 22.1000 69.0000 22.2000 ;
	    RECT 46.2000 21.8000 69.0000 22.1000 ;
	    RECT 85.4000 22.1000 85.8000 22.2000 ;
	    RECT 97.4000 22.1000 97.8000 22.2000 ;
	    RECT 100.6000 22.1000 101.0000 22.2000 ;
	    RECT 85.4000 21.8000 101.0000 22.1000 ;
	    RECT 119.0000 22.1000 119.4000 22.2000 ;
	    RECT 143.0000 22.1000 143.4000 22.2000 ;
	    RECT 161.4000 22.1000 161.8000 22.2000 ;
	    RECT 119.0000 21.8000 161.8000 22.1000 ;
	    RECT 255.8000 22.1000 256.2000 22.2000 ;
	    RECT 257.4000 22.1000 257.8000 22.2000 ;
	    RECT 255.8000 21.8000 257.8000 22.1000 ;
	    RECT 89.4000 21.1000 89.8000 21.2000 ;
	    RECT 99.0000 21.1000 99.4000 21.2000 ;
	    RECT 89.4000 20.8000 99.4000 21.1000 ;
	    RECT 207.0000 19.1000 207.4000 19.2000 ;
	    RECT 224.6000 19.1000 225.0000 19.2000 ;
	    RECT 238.2000 19.1000 238.6000 19.2000 ;
	    RECT 247.8000 19.1000 248.2000 19.2000 ;
	    RECT 250.2000 19.1000 250.6000 19.2000 ;
	    RECT 207.0000 18.8000 250.6000 19.1000 ;
	    RECT 67.8000 17.8000 68.2000 18.2000 ;
	    RECT 251.0000 17.8000 251.4000 18.2000 ;
	    RECT 67.8000 17.2000 68.1000 17.8000 ;
	    RECT 53.4000 17.1000 53.8000 17.2000 ;
	    RECT 63.0000 17.1000 63.4000 17.2000 ;
	    RECT 53.4000 16.8000 63.4000 17.1000 ;
	    RECT 67.8000 16.8000 68.2000 17.2000 ;
	    RECT 69.4000 16.8000 69.8000 17.2000 ;
	    RECT 205.4000 17.1000 205.8000 17.2000 ;
	    RECT 207.0000 17.1000 207.4000 17.2000 ;
	    RECT 205.4000 16.8000 207.4000 17.1000 ;
	    RECT 209.4000 17.1000 209.8000 17.2000 ;
	    RECT 223.0000 17.1000 223.4000 17.2000 ;
	    RECT 209.4000 16.8000 223.4000 17.1000 ;
	    RECT 227.8000 17.1000 228.2000 17.2000 ;
	    RECT 231.0000 17.1000 231.4000 17.2000 ;
	    RECT 235.0000 17.1000 235.4000 17.2000 ;
	    RECT 227.8000 16.8000 235.4000 17.1000 ;
	    RECT 240.6000 17.1000 241.0000 17.2000 ;
	    RECT 251.0000 17.1000 251.3000 17.8000 ;
	    RECT 240.6000 16.8000 251.3000 17.1000 ;
	    RECT 39.8000 15.8000 40.2000 16.2000 ;
	    RECT 59.0000 16.1000 59.4000 16.2000 ;
	    RECT 65.4000 16.1000 65.8000 16.2000 ;
	    RECT 69.4000 16.1000 69.7000 16.8000 ;
	    RECT 59.0000 15.8000 64.1000 16.1000 ;
	    RECT 65.4000 15.8000 69.7000 16.1000 ;
	    RECT 71.8000 16.1000 72.2000 16.2000 ;
	    RECT 82.2000 16.1000 82.6000 16.2000 ;
	    RECT 71.8000 15.8000 82.6000 16.1000 ;
	    RECT 87.0000 16.1000 87.4000 16.2000 ;
	    RECT 91.0000 16.1000 91.4000 16.2000 ;
	    RECT 87.0000 15.8000 91.4000 16.1000 ;
	    RECT 110.2000 16.1000 110.6000 16.2000 ;
	    RECT 113.4000 16.1000 113.8000 16.2000 ;
	    RECT 110.2000 15.8000 113.8000 16.1000 ;
	    RECT 118.2000 15.8000 118.6000 16.2000 ;
	    RECT 131.0000 16.1000 131.4000 16.2000 ;
	    RECT 137.4000 16.1000 137.8000 16.2000 ;
	    RECT 131.0000 15.8000 137.8000 16.1000 ;
	    RECT 157.4000 15.8000 157.8000 16.2000 ;
	    RECT 169.4000 16.1000 169.8000 16.2000 ;
	    RECT 176.6000 16.1000 177.0000 16.2000 ;
	    RECT 169.4000 15.8000 177.0000 16.1000 ;
	    RECT 187.8000 16.1000 188.2000 16.2000 ;
	    RECT 198.2000 16.1000 198.6000 16.2000 ;
	    RECT 187.8000 15.8000 198.6000 16.1000 ;
	    RECT 200.6000 16.1000 201.0000 16.2000 ;
	    RECT 251.8000 16.1000 252.2000 16.2000 ;
	    RECT 263.8000 16.1000 264.2000 16.2000 ;
	    RECT 200.6000 15.8000 252.2000 16.1000 ;
	    RECT 252.6000 15.8000 264.2000 16.1000 ;
	    RECT 3.0000 15.1000 3.4000 15.2000 ;
	    RECT 9.4000 15.1000 9.8000 15.2000 ;
	    RECT 3.0000 14.8000 9.8000 15.1000 ;
	    RECT 15.8000 15.1000 16.2000 15.2000 ;
	    RECT 23.0000 15.1000 23.4000 15.2000 ;
	    RECT 15.8000 14.8000 23.4000 15.1000 ;
	    RECT 26.2000 14.8000 26.6000 15.2000 ;
	    RECT 31.0000 14.8000 31.4000 15.2000 ;
	    RECT 34.2000 15.1000 34.6000 15.2000 ;
	    RECT 39.8000 15.1000 40.1000 15.8000 ;
	    RECT 63.8000 15.2000 64.1000 15.8000 ;
	    RECT 34.2000 14.8000 40.1000 15.1000 ;
	    RECT 43.8000 15.1000 44.2000 15.2000 ;
	    RECT 47.0000 15.1000 47.4000 15.2000 ;
	    RECT 43.8000 14.8000 47.4000 15.1000 ;
	    RECT 63.8000 14.8000 64.2000 15.2000 ;
	    RECT 67.8000 15.1000 68.2000 15.2000 ;
	    RECT 70.2000 15.1000 70.6000 15.2000 ;
	    RECT 67.8000 14.8000 70.6000 15.1000 ;
	    RECT 71.8000 15.1000 72.2000 15.2000 ;
	    RECT 91.8000 15.1000 92.2000 15.2000 ;
	    RECT 92.6000 15.1000 93.0000 15.2000 ;
	    RECT 71.8000 14.8000 84.9000 15.1000 ;
	    RECT 91.8000 14.8000 93.0000 15.1000 ;
	    RECT 94.2000 15.1000 94.6000 15.2000 ;
	    RECT 95.0000 15.1000 95.4000 15.2000 ;
	    RECT 94.2000 14.8000 95.4000 15.1000 ;
	    RECT 111.8000 15.1000 112.2000 15.2000 ;
	    RECT 115.8000 15.1000 116.2000 15.2000 ;
	    RECT 111.8000 14.8000 116.2000 15.1000 ;
	    RECT 118.2000 15.1000 118.5000 15.8000 ;
	    RECT 157.4000 15.2000 157.7000 15.8000 ;
	    RECT 252.6000 15.2000 252.9000 15.8000 ;
	    RECT 122.2000 15.1000 122.6000 15.2000 ;
	    RECT 118.2000 14.8000 122.6000 15.1000 ;
	    RECT 123.0000 15.1000 123.4000 15.2000 ;
	    RECT 138.2000 15.1000 138.6000 15.2000 ;
	    RECT 123.0000 14.8000 138.6000 15.1000 ;
	    RECT 147.8000 15.1000 148.2000 15.2000 ;
	    RECT 155.0000 15.1000 155.4000 15.2000 ;
	    RECT 147.8000 14.8000 155.4000 15.1000 ;
	    RECT 157.4000 14.8000 157.8000 15.2000 ;
	    RECT 173.4000 15.1000 173.8000 15.2000 ;
	    RECT 183.0000 15.1000 183.4000 15.2000 ;
	    RECT 173.4000 14.8000 183.4000 15.1000 ;
	    RECT 188.6000 15.1000 189.0000 15.2000 ;
	    RECT 192.6000 15.1000 193.0000 15.2000 ;
	    RECT 188.6000 14.8000 193.0000 15.1000 ;
	    RECT 199.8000 15.1000 200.2000 15.2000 ;
	    RECT 206.2000 15.1000 206.6000 15.2000 ;
	    RECT 199.8000 14.8000 206.6000 15.1000 ;
	    RECT 207.8000 15.1000 208.2000 15.2000 ;
	    RECT 211.0000 15.1000 211.4000 15.2000 ;
	    RECT 207.8000 14.8000 211.4000 15.1000 ;
	    RECT 218.2000 15.1000 218.6000 15.2000 ;
	    RECT 223.0000 15.1000 223.4000 15.2000 ;
	    RECT 223.8000 15.1000 224.2000 15.2000 ;
	    RECT 218.2000 14.8000 220.1000 15.1000 ;
	    RECT 223.0000 14.8000 224.2000 15.1000 ;
	    RECT 233.4000 15.1000 233.8000 15.2000 ;
	    RECT 235.8000 15.1000 236.2000 15.2000 ;
	    RECT 233.4000 14.8000 236.2000 15.1000 ;
	    RECT 239.8000 15.1000 240.2000 15.2000 ;
	    RECT 246.2000 15.1000 246.6000 15.2000 ;
	    RECT 247.0000 15.1000 247.4000 15.2000 ;
	    RECT 239.8000 14.8000 247.4000 15.1000 ;
	    RECT 248.6000 14.8000 249.0000 15.2000 ;
	    RECT 252.6000 14.8000 253.0000 15.2000 ;
	    RECT 259.0000 14.8000 259.4000 15.2000 ;
	    RECT 26.2000 14.1000 26.5000 14.8000 ;
	    RECT 31.0000 14.1000 31.3000 14.8000 ;
	    RECT 84.6000 14.2000 84.9000 14.8000 ;
	    RECT 123.0000 14.2000 123.3000 14.8000 ;
	    RECT 219.8000 14.2000 220.1000 14.8000 ;
	    RECT 26.2000 13.8000 31.3000 14.1000 ;
	    RECT 50.2000 14.1000 50.6000 14.2000 ;
	    RECT 60.6000 14.1000 61.0000 14.2000 ;
	    RECT 50.2000 13.8000 61.0000 14.1000 ;
	    RECT 63.0000 14.1000 63.4000 14.2000 ;
	    RECT 65.4000 14.1000 65.8000 14.2000 ;
	    RECT 67.0000 14.1000 67.4000 14.2000 ;
	    RECT 63.0000 13.8000 67.4000 14.1000 ;
	    RECT 67.8000 13.8000 68.2000 14.2000 ;
	    RECT 68.6000 14.1000 69.0000 14.2000 ;
	    RECT 71.8000 14.1000 72.2000 14.2000 ;
	    RECT 78.2000 14.1000 78.6000 14.2000 ;
	    RECT 68.6000 13.8000 78.6000 14.1000 ;
	    RECT 84.6000 13.8000 85.0000 14.2000 ;
	    RECT 88.6000 14.1000 89.0000 14.2000 ;
	    RECT 89.4000 14.1000 89.8000 14.2000 ;
	    RECT 88.6000 13.8000 89.8000 14.1000 ;
	    RECT 99.8000 14.1000 100.2000 14.2000 ;
	    RECT 102.2000 14.1000 102.6000 14.2000 ;
	    RECT 111.0000 14.1000 111.4000 14.2000 ;
	    RECT 99.8000 13.8000 111.4000 14.1000 ;
	    RECT 115.8000 14.1000 116.2000 14.2000 ;
	    RECT 123.0000 14.1000 123.4000 14.2000 ;
	    RECT 115.8000 13.8000 123.4000 14.1000 ;
	    RECT 137.4000 14.1000 137.8000 14.2000 ;
	    RECT 147.0000 14.1000 147.4000 14.2000 ;
	    RECT 137.4000 13.8000 147.4000 14.1000 ;
	    RECT 179.8000 14.1000 180.2000 14.2000 ;
	    RECT 184.6000 14.1000 185.0000 14.2000 ;
	    RECT 179.8000 13.8000 185.0000 14.1000 ;
	    RECT 203.8000 14.1000 204.2000 14.2000 ;
	    RECT 205.4000 14.1000 205.8000 14.2000 ;
	    RECT 214.2000 14.1000 214.6000 14.2000 ;
	    RECT 203.8000 13.8000 214.6000 14.1000 ;
	    RECT 219.8000 13.8000 220.2000 14.2000 ;
	    RECT 227.0000 14.1000 227.4000 14.2000 ;
	    RECT 228.6000 14.1000 229.0000 14.2000 ;
	    RECT 241.4000 14.1000 241.8000 14.2000 ;
	    RECT 246.2000 14.1000 246.6000 14.2000 ;
	    RECT 248.6000 14.1000 248.9000 14.8000 ;
	    RECT 259.0000 14.2000 259.3000 14.8000 ;
	    RECT 227.0000 13.8000 248.9000 14.1000 ;
	    RECT 252.6000 13.8000 253.0000 14.2000 ;
	    RECT 256.6000 13.8000 257.0000 14.2000 ;
	    RECT 259.0000 13.8000 259.4000 14.2000 ;
	    RECT 67.8000 13.2000 68.1000 13.8000 ;
	    RECT 252.6000 13.2000 252.9000 13.8000 ;
	    RECT 256.6000 13.2000 256.9000 13.8000 ;
	    RECT 4.6000 12.8000 5.0000 13.2000 ;
	    RECT 49.4000 13.1000 49.8000 13.2000 ;
	    RECT 56.6000 13.1000 57.0000 13.2000 ;
	    RECT 49.4000 12.8000 57.0000 13.1000 ;
	    RECT 67.8000 13.1000 68.2000 13.2000 ;
	    RECT 80.6000 13.1000 81.0000 13.2000 ;
	    RECT 84.6000 13.1000 85.0000 13.2000 ;
	    RECT 67.8000 12.8000 85.0000 13.1000 ;
	    RECT 90.2000 13.1000 90.6000 13.2000 ;
	    RECT 92.6000 13.1000 93.0000 13.2000 ;
	    RECT 90.2000 12.8000 93.0000 13.1000 ;
	    RECT 94.2000 13.1000 94.6000 13.2000 ;
	    RECT 95.0000 13.1000 95.4000 13.2000 ;
	    RECT 94.2000 12.8000 95.4000 13.1000 ;
	    RECT 98.2000 13.1000 98.6000 13.2000 ;
	    RECT 100.6000 13.1000 101.0000 13.2000 ;
	    RECT 101.4000 13.1000 101.8000 13.2000 ;
	    RECT 98.2000 12.8000 101.8000 13.1000 ;
	    RECT 102.2000 13.1000 102.6000 13.2000 ;
	    RECT 105.4000 13.1000 105.8000 13.2000 ;
	    RECT 102.2000 12.8000 105.8000 13.1000 ;
	    RECT 113.4000 13.1000 113.8000 13.2000 ;
	    RECT 119.0000 13.1000 119.4000 13.2000 ;
	    RECT 113.4000 12.8000 119.4000 13.1000 ;
	    RECT 119.8000 13.1000 120.2000 13.2000 ;
	    RECT 123.0000 13.1000 123.4000 13.2000 ;
	    RECT 119.8000 12.8000 123.4000 13.1000 ;
	    RECT 124.6000 13.1000 125.0000 13.2000 ;
	    RECT 136.6000 13.1000 137.0000 13.2000 ;
	    RECT 124.6000 12.8000 137.0000 13.1000 ;
	    RECT 155.0000 13.1000 155.4000 13.2000 ;
	    RECT 162.2000 13.1000 162.6000 13.2000 ;
	    RECT 169.4000 13.1000 169.8000 13.2000 ;
	    RECT 155.0000 12.8000 169.8000 13.1000 ;
	    RECT 195.0000 12.8000 195.4000 13.2000 ;
	    RECT 207.0000 13.1000 207.4000 13.2000 ;
	    RECT 210.2000 13.1000 210.6000 13.2000 ;
	    RECT 216.6000 13.1000 217.0000 13.2000 ;
	    RECT 207.0000 12.8000 217.0000 13.1000 ;
	    RECT 224.6000 13.1000 225.0000 13.2000 ;
	    RECT 229.4000 13.1000 229.8000 13.2000 ;
	    RECT 237.4000 13.1000 237.8000 13.2000 ;
	    RECT 242.2000 13.1000 242.6000 13.2000 ;
	    RECT 248.6000 13.1000 249.0000 13.2000 ;
	    RECT 224.6000 12.8000 249.0000 13.1000 ;
	    RECT 252.6000 12.8000 253.0000 13.2000 ;
	    RECT 256.6000 12.8000 257.0000 13.2000 ;
	    RECT 1.4000 12.1000 1.8000 12.2000 ;
	    RECT 2.2000 12.1000 2.6000 12.2000 ;
	    RECT 4.6000 12.1000 4.9000 12.8000 ;
	    RECT 1.4000 11.8000 4.9000 12.1000 ;
	    RECT 39.8000 12.1000 40.2000 12.2000 ;
	    RECT 41.4000 12.1000 41.8000 12.2000 ;
	    RECT 47.0000 12.1000 47.4000 12.2000 ;
	    RECT 39.8000 11.8000 47.4000 12.1000 ;
	    RECT 50.2000 12.1000 50.6000 12.2000 ;
	    RECT 52.6000 12.1000 53.0000 12.2000 ;
	    RECT 50.2000 11.8000 53.0000 12.1000 ;
	    RECT 75.0000 12.1000 75.4000 12.2000 ;
	    RECT 88.6000 12.1000 89.0000 12.2000 ;
	    RECT 111.0000 12.1000 111.4000 12.2000 ;
	    RECT 117.4000 12.1000 117.8000 12.2000 ;
	    RECT 75.0000 11.8000 110.5000 12.1000 ;
	    RECT 111.0000 11.8000 117.8000 12.1000 ;
	    RECT 120.6000 12.1000 121.0000 12.2000 ;
	    RECT 123.8000 12.1000 124.2000 12.2000 ;
	    RECT 120.6000 11.8000 124.2000 12.1000 ;
	    RECT 124.6000 12.1000 125.0000 12.2000 ;
	    RECT 132.6000 12.1000 133.0000 12.2000 ;
	    RECT 124.6000 11.8000 133.0000 12.1000 ;
	    RECT 134.2000 12.1000 134.6000 12.2000 ;
	    RECT 141.4000 12.1000 141.8000 12.2000 ;
	    RECT 134.2000 11.8000 141.8000 12.1000 ;
	    RECT 195.0000 12.1000 195.3000 12.8000 ;
	    RECT 213.4000 12.1000 213.8000 12.2000 ;
	    RECT 195.0000 11.8000 213.8000 12.1000 ;
	    RECT 255.0000 12.1000 255.4000 12.2000 ;
	    RECT 267.8000 12.1000 268.2000 12.2000 ;
	    RECT 268.6000 12.1000 269.0000 12.2000 ;
	    RECT 255.0000 11.8000 269.0000 12.1000 ;
	    RECT 87.0000 11.1000 87.4000 11.2000 ;
	    RECT 98.2000 11.1000 98.6000 11.2000 ;
	    RECT 87.0000 10.8000 98.6000 11.1000 ;
	    RECT 104.6000 11.1000 105.0000 11.2000 ;
	    RECT 105.4000 11.1000 105.8000 11.2000 ;
	    RECT 104.6000 10.8000 105.8000 11.1000 ;
	    RECT 110.2000 11.1000 110.5000 11.8000 ;
	    RECT 143.8000 11.1000 144.2000 11.2000 ;
	    RECT 110.2000 10.8000 144.2000 11.1000 ;
	    RECT 215.8000 11.1000 216.2000 11.2000 ;
	    RECT 234.2000 11.1000 234.6000 11.2000 ;
	    RECT 255.0000 11.1000 255.4000 11.2000 ;
	    RECT 215.8000 10.8000 255.4000 11.1000 ;
	    RECT 263.0000 11.1000 263.4000 11.2000 ;
	    RECT 269.4000 11.1000 269.8000 11.2000 ;
	    RECT 263.0000 10.8000 269.8000 11.1000 ;
	    RECT 47.0000 10.1000 47.4000 10.2000 ;
	    RECT 58.2000 10.1000 58.6000 10.2000 ;
	    RECT 64.6000 10.1000 65.0000 10.2000 ;
	    RECT 47.0000 9.8000 65.0000 10.1000 ;
	    RECT 86.2000 10.1000 86.6000 10.2000 ;
	    RECT 89.4000 10.1000 89.8000 10.2000 ;
	    RECT 86.2000 9.8000 89.8000 10.1000 ;
	    RECT 110.2000 10.1000 110.6000 10.2000 ;
	    RECT 112.6000 10.1000 113.0000 10.2000 ;
	    RECT 110.2000 9.8000 113.0000 10.1000 ;
	    RECT 116.6000 10.1000 117.0000 10.2000 ;
	    RECT 124.6000 10.1000 125.0000 10.2000 ;
	    RECT 151.0000 10.1000 151.4000 10.2000 ;
	    RECT 153.4000 10.1000 153.8000 10.2000 ;
	    RECT 159.0000 10.1000 159.4000 10.2000 ;
	    RECT 164.6000 10.1000 165.0000 10.2000 ;
	    RECT 175.8000 10.1000 176.2000 10.2000 ;
	    RECT 116.6000 9.8000 140.1000 10.1000 ;
	    RECT 151.0000 9.8000 176.2000 10.1000 ;
	    RECT 181.4000 10.1000 181.8000 10.2000 ;
	    RECT 191.0000 10.1000 191.4000 10.2000 ;
	    RECT 205.4000 10.1000 205.8000 10.2000 ;
	    RECT 181.4000 9.8000 205.8000 10.1000 ;
	    RECT 221.4000 10.1000 221.8000 10.2000 ;
	    RECT 233.4000 10.1000 233.8000 10.2000 ;
	    RECT 241.4000 10.1000 241.8000 10.2000 ;
	    RECT 221.4000 9.8000 232.1000 10.1000 ;
	    RECT 233.4000 9.8000 241.8000 10.1000 ;
	    RECT 253.4000 10.1000 253.8000 10.2000 ;
	    RECT 257.4000 10.1000 257.8000 10.2000 ;
	    RECT 253.4000 9.8000 257.8000 10.1000 ;
	    RECT 139.8000 9.2000 140.1000 9.8000 ;
	    RECT 5.4000 9.1000 5.8000 9.2000 ;
	    RECT 8.6000 9.1000 9.0000 9.2000 ;
	    RECT 5.4000 8.8000 9.0000 9.1000 ;
	    RECT 12.6000 9.1000 13.0000 9.2000 ;
	    RECT 15.8000 9.1000 16.2000 9.2000 ;
	    RECT 26.2000 9.1000 26.6000 9.2000 ;
	    RECT 27.8000 9.1000 28.2000 9.2000 ;
	    RECT 43.8000 9.1000 44.2000 9.2000 ;
	    RECT 12.6000 8.8000 44.2000 9.1000 ;
	    RECT 55.8000 9.1000 56.2000 9.2000 ;
	    RECT 63.8000 9.1000 64.2000 9.2000 ;
	    RECT 55.8000 8.8000 64.2000 9.1000 ;
	    RECT 67.0000 9.1000 67.4000 9.2000 ;
	    RECT 73.4000 9.1000 73.8000 9.2000 ;
	    RECT 67.0000 8.8000 73.8000 9.1000 ;
	    RECT 74.2000 9.1000 74.6000 9.2000 ;
	    RECT 91.0000 9.1000 91.4000 9.2000 ;
	    RECT 94.2000 9.1000 94.6000 9.2000 ;
	    RECT 74.2000 8.8000 94.6000 9.1000 ;
	    RECT 105.4000 9.1000 105.8000 9.2000 ;
	    RECT 106.2000 9.1000 106.6000 9.2000 ;
	    RECT 111.0000 9.1000 111.4000 9.2000 ;
	    RECT 105.4000 8.8000 111.4000 9.1000 ;
	    RECT 115.8000 9.1000 116.2000 9.2000 ;
	    RECT 125.4000 9.1000 125.8000 9.2000 ;
	    RECT 130.2000 9.1000 130.6000 9.2000 ;
	    RECT 134.2000 9.1000 134.6000 9.2000 ;
	    RECT 115.8000 8.8000 134.6000 9.1000 ;
	    RECT 139.8000 9.1000 140.2000 9.2000 ;
	    RECT 154.2000 9.1000 154.6000 9.2000 ;
	    RECT 139.8000 8.8000 154.6000 9.1000 ;
	    RECT 170.2000 9.1000 170.6000 9.2000 ;
	    RECT 171.8000 9.1000 172.2000 9.2000 ;
	    RECT 170.2000 8.8000 172.2000 9.1000 ;
	    RECT 189.4000 9.1000 189.8000 9.2000 ;
	    RECT 218.2000 9.1000 218.6000 9.2000 ;
	    RECT 227.0000 9.1000 227.4000 9.2000 ;
	    RECT 189.4000 8.8000 227.4000 9.1000 ;
	    RECT 231.8000 9.1000 232.1000 9.8000 ;
	    RECT 241.4000 9.1000 241.8000 9.2000 ;
	    RECT 231.8000 8.8000 241.8000 9.1000 ;
	    RECT 257.4000 9.1000 257.8000 9.2000 ;
	    RECT 262.2000 9.1000 262.6000 9.2000 ;
	    RECT 257.4000 8.8000 262.6000 9.1000 ;
	    RECT 268.6000 8.8000 269.0000 9.2000 ;
	    RECT 268.6000 8.2000 268.9000 8.8000 ;
	    RECT 24.6000 8.1000 25.0000 8.2000 ;
	    RECT 34.2000 8.1000 34.6000 8.2000 ;
	    RECT 24.6000 7.8000 34.6000 8.1000 ;
	    RECT 40.6000 8.1000 41.0000 8.2000 ;
	    RECT 50.2000 8.1000 50.6000 8.2000 ;
	    RECT 40.6000 7.8000 50.6000 8.1000 ;
	    RECT 60.6000 8.1000 61.0000 8.2000 ;
	    RECT 75.0000 8.1000 75.4000 8.2000 ;
	    RECT 60.6000 7.8000 75.4000 8.1000 ;
	    RECT 79.8000 8.1000 80.2000 8.2000 ;
	    RECT 83.8000 8.1000 84.2000 8.2000 ;
	    RECT 79.8000 7.8000 84.2000 8.1000 ;
	    RECT 91.8000 7.8000 92.2000 8.2000 ;
	    RECT 98.2000 8.1000 98.6000 8.2000 ;
	    RECT 100.6000 8.1000 101.0000 8.2000 ;
	    RECT 98.2000 7.8000 101.0000 8.1000 ;
	    RECT 103.0000 8.1000 103.4000 8.2000 ;
	    RECT 103.8000 8.1000 104.2000 8.2000 ;
	    RECT 116.6000 8.1000 117.0000 8.2000 ;
	    RECT 103.0000 7.8000 117.0000 8.1000 ;
	    RECT 117.4000 8.1000 117.8000 8.2000 ;
	    RECT 121.4000 8.1000 121.8000 8.2000 ;
	    RECT 117.4000 7.8000 121.8000 8.1000 ;
	    RECT 122.2000 8.1000 122.6000 8.2000 ;
	    RECT 123.0000 8.1000 123.4000 8.2000 ;
	    RECT 122.2000 7.8000 123.4000 8.1000 ;
	    RECT 125.4000 7.8000 125.8000 8.2000 ;
	    RECT 131.0000 8.1000 131.4000 8.2000 ;
	    RECT 131.8000 8.1000 132.2000 8.2000 ;
	    RECT 131.0000 7.8000 132.2000 8.1000 ;
	    RECT 135.0000 8.1000 135.4000 8.2000 ;
	    RECT 136.6000 8.1000 137.0000 8.2000 ;
	    RECT 152.6000 8.1000 153.0000 8.2000 ;
	    RECT 135.0000 7.8000 153.0000 8.1000 ;
	    RECT 184.6000 8.1000 185.0000 8.2000 ;
	    RECT 194.2000 8.1000 194.6000 8.2000 ;
	    RECT 184.6000 7.8000 194.6000 8.1000 ;
	    RECT 198.2000 8.1000 198.6000 8.2000 ;
	    RECT 222.2000 8.1000 222.6000 8.2000 ;
	    RECT 198.2000 7.8000 222.6000 8.1000 ;
	    RECT 223.8000 8.1000 224.2000 8.2000 ;
	    RECT 229.4000 8.1000 229.8000 8.2000 ;
	    RECT 223.8000 7.8000 229.8000 8.1000 ;
	    RECT 251.0000 8.1000 251.4000 8.2000 ;
	    RECT 252.6000 8.1000 253.0000 8.2000 ;
	    RECT 251.0000 7.8000 253.0000 8.1000 ;
	    RECT 256.6000 8.1000 257.0000 8.2000 ;
	    RECT 259.0000 8.1000 259.4000 8.2000 ;
	    RECT 256.6000 7.8000 259.4000 8.1000 ;
	    RECT 263.8000 7.8000 264.2000 8.2000 ;
	    RECT 268.6000 7.8000 269.0000 8.2000 ;
	    RECT 38.2000 6.8000 38.6000 7.2000 ;
	    RECT 52.6000 7.1000 53.0000 7.2000 ;
	    RECT 69.4000 7.1000 69.8000 7.2000 ;
	    RECT 70.2000 7.1000 70.6000 7.2000 ;
	    RECT 52.6000 6.8000 70.6000 7.1000 ;
	    RECT 73.4000 7.1000 73.8000 7.2000 ;
	    RECT 77.4000 7.1000 77.8000 7.2000 ;
	    RECT 73.4000 6.8000 77.8000 7.1000 ;
	    RECT 78.2000 7.1000 78.6000 7.2000 ;
	    RECT 80.6000 7.1000 81.0000 7.2000 ;
	    RECT 78.2000 6.8000 81.0000 7.1000 ;
	    RECT 82.2000 7.1000 82.6000 7.2000 ;
	    RECT 85.4000 7.1000 85.8000 7.2000 ;
	    RECT 82.2000 6.8000 85.8000 7.1000 ;
	    RECT 89.4000 7.1000 89.8000 7.2000 ;
	    RECT 91.8000 7.1000 92.1000 7.8000 ;
	    RECT 89.4000 6.8000 92.1000 7.1000 ;
	    RECT 93.4000 7.1000 93.8000 7.2000 ;
	    RECT 96.6000 7.1000 97.0000 7.2000 ;
	    RECT 93.4000 6.8000 97.0000 7.1000 ;
	    RECT 98.2000 7.1000 98.6000 7.2000 ;
	    RECT 99.0000 7.1000 99.4000 7.2000 ;
	    RECT 98.2000 6.8000 99.4000 7.1000 ;
	    RECT 99.8000 7.1000 100.2000 7.2000 ;
	    RECT 102.2000 7.1000 102.6000 7.2000 ;
	    RECT 99.8000 6.8000 102.6000 7.1000 ;
	    RECT 103.8000 7.1000 104.2000 7.2000 ;
	    RECT 105.4000 7.1000 105.8000 7.2000 ;
	    RECT 103.8000 6.8000 105.8000 7.1000 ;
	    RECT 111.0000 7.1000 111.4000 7.2000 ;
	    RECT 125.4000 7.1000 125.7000 7.8000 ;
	    RECT 111.0000 6.8000 125.7000 7.1000 ;
	    RECT 131.0000 7.1000 131.4000 7.2000 ;
	    RECT 137.4000 7.1000 137.8000 7.2000 ;
	    RECT 131.0000 6.8000 137.8000 7.1000 ;
	    RECT 191.0000 6.8000 191.4000 7.2000 ;
	    RECT 198.2000 7.1000 198.6000 7.2000 ;
	    RECT 203.8000 7.1000 204.2000 7.2000 ;
	    RECT 213.4000 7.1000 213.8000 7.2000 ;
	    RECT 198.2000 6.8000 213.8000 7.1000 ;
	    RECT 227.8000 7.1000 228.2000 7.2000 ;
	    RECT 231.8000 7.1000 232.2000 7.2000 ;
	    RECT 245.4000 7.1000 245.8000 7.2000 ;
	    RECT 227.8000 6.8000 245.8000 7.1000 ;
	    RECT 250.2000 7.1000 250.6000 7.2000 ;
	    RECT 263.8000 7.1000 264.1000 7.8000 ;
	    RECT 250.2000 6.8000 264.1000 7.1000 ;
	    RECT 38.2000 6.2000 38.5000 6.8000 ;
	    RECT 3.8000 6.1000 4.2000 6.2000 ;
	    RECT 9.4000 6.1000 9.8000 6.2000 ;
	    RECT 14.2000 6.1000 14.6000 6.2000 ;
	    RECT 22.2000 6.1000 22.6000 6.2000 ;
	    RECT 38.2000 6.1000 38.6000 6.2000 ;
	    RECT 3.8000 5.8000 38.6000 6.1000 ;
	    RECT 39.0000 6.1000 39.4000 6.2000 ;
	    RECT 63.8000 6.1000 64.2000 6.2000 ;
	    RECT 70.2000 6.1000 70.6000 6.2000 ;
	    RECT 39.0000 5.8000 44.1000 6.1000 ;
	    RECT 63.8000 5.8000 70.6000 6.1000 ;
	    RECT 76.6000 6.1000 77.0000 6.2000 ;
	    RECT 81.4000 6.1000 81.8000 6.2000 ;
	    RECT 76.6000 5.8000 81.8000 6.1000 ;
	    RECT 86.2000 6.1000 86.6000 6.2000 ;
	    RECT 89.4000 6.1000 89.8000 6.2000 ;
	    RECT 94.2000 6.1000 94.6000 6.2000 ;
	    RECT 86.2000 5.8000 94.6000 6.1000 ;
	    RECT 101.4000 6.1000 101.8000 6.2000 ;
	    RECT 103.0000 6.1000 103.4000 6.2000 ;
	    RECT 117.4000 6.1000 117.8000 6.2000 ;
	    RECT 101.4000 5.8000 117.8000 6.1000 ;
	    RECT 118.2000 6.1000 118.6000 6.2000 ;
	    RECT 120.6000 6.1000 121.0000 6.2000 ;
	    RECT 170.2000 6.1000 170.6000 6.2000 ;
	    RECT 177.4000 6.1000 177.8000 6.2000 ;
	    RECT 118.2000 5.8000 170.6000 6.1000 ;
	    RECT 171.8000 5.8000 177.8000 6.1000 ;
	    RECT 191.0000 6.1000 191.3000 6.8000 ;
	    RECT 195.8000 6.1000 196.2000 6.2000 ;
	    RECT 191.0000 5.8000 196.2000 6.1000 ;
	    RECT 202.2000 6.1000 202.6000 6.2000 ;
	    RECT 215.8000 6.1000 216.2000 6.2000 ;
	    RECT 228.6000 6.1000 229.0000 6.2000 ;
	    RECT 202.2000 5.8000 207.3000 6.1000 ;
	    RECT 215.8000 5.8000 229.0000 6.1000 ;
	    RECT 233.4000 6.1000 233.8000 6.2000 ;
	    RECT 235.8000 6.1000 236.2000 6.2000 ;
	    RECT 233.4000 5.8000 236.2000 6.1000 ;
	    RECT 239.8000 5.8000 240.2000 6.2000 ;
	    RECT 242.2000 6.1000 242.6000 6.2000 ;
	    RECT 251.8000 6.1000 252.2000 6.2000 ;
	    RECT 242.2000 5.8000 252.2000 6.1000 ;
	    RECT 255.0000 6.1000 255.4000 6.2000 ;
	    RECT 255.8000 6.1000 256.2000 6.2000 ;
	    RECT 255.0000 5.8000 256.2000 6.1000 ;
	    RECT 43.8000 5.2000 44.1000 5.8000 ;
	    RECT 171.8000 5.2000 172.1000 5.8000 ;
	    RECT 207.0000 5.2000 207.3000 5.8000 ;
	    RECT 8.6000 5.1000 9.0000 5.2000 ;
	    RECT 15.0000 5.1000 15.4000 5.2000 ;
	    RECT 27.8000 5.1000 28.2000 5.2000 ;
	    RECT 8.6000 4.8000 15.4000 5.1000 ;
	    RECT 22.2000 4.8000 28.2000 5.1000 ;
	    RECT 43.8000 4.8000 44.2000 5.2000 ;
	    RECT 83.0000 5.1000 83.4000 5.2000 ;
	    RECT 87.0000 5.1000 87.4000 5.2000 ;
	    RECT 83.0000 4.8000 87.4000 5.1000 ;
	    RECT 95.8000 5.1000 96.2000 5.2000 ;
	    RECT 113.4000 5.1000 113.8000 5.2000 ;
	    RECT 95.8000 4.8000 113.8000 5.1000 ;
	    RECT 116.6000 5.1000 117.0000 5.2000 ;
	    RECT 122.2000 5.1000 122.6000 5.2000 ;
	    RECT 116.6000 4.8000 122.6000 5.1000 ;
	    RECT 126.2000 5.1000 126.6000 5.2000 ;
	    RECT 127.0000 5.1000 127.4000 5.2000 ;
	    RECT 126.2000 4.8000 127.4000 5.1000 ;
	    RECT 135.8000 5.1000 136.2000 5.2000 ;
	    RECT 138.2000 5.1000 138.6000 5.2000 ;
	    RECT 135.8000 4.8000 138.6000 5.1000 ;
	    RECT 142.2000 5.1000 142.6000 5.2000 ;
	    RECT 142.2000 4.8000 154.5000 5.1000 ;
	    RECT 171.8000 4.8000 172.2000 5.2000 ;
	    RECT 186.2000 5.1000 186.6000 5.2000 ;
	    RECT 197.4000 5.1000 197.8000 5.2000 ;
	    RECT 200.6000 5.1000 201.0000 5.2000 ;
	    RECT 186.2000 4.8000 201.0000 5.1000 ;
	    RECT 207.0000 4.8000 207.4000 5.2000 ;
	    RECT 239.8000 5.1000 240.1000 5.8000 ;
	    RECT 246.2000 5.1000 246.6000 5.2000 ;
	    RECT 239.8000 4.8000 246.6000 5.1000 ;
	    RECT 260.6000 5.1000 261.0000 5.2000 ;
	    RECT 261.4000 5.1000 261.8000 5.2000 ;
	    RECT 265.4000 5.1000 265.8000 5.2000 ;
	    RECT 260.6000 4.8000 265.8000 5.1000 ;
	    RECT 22.2000 4.2000 22.5000 4.8000 ;
	    RECT 154.2000 4.2000 154.5000 4.8000 ;
	    RECT 22.2000 3.8000 22.6000 4.2000 ;
	    RECT 154.2000 3.8000 154.6000 4.2000 ;
         LAYER metal4 ;
	    RECT 92.6000 174.8000 93.0000 175.2000 ;
	    RECT 219.0000 174.8000 219.4000 175.2000 ;
	    RECT 223.8000 175.1000 224.2000 175.2000 ;
	    RECT 223.0000 174.8000 224.2000 175.1000 ;
	    RECT 14.2000 171.8000 14.6000 172.2000 ;
	    RECT 14.2000 156.2000 14.5000 171.8000 ;
	    RECT 92.6000 166.2000 92.9000 174.8000 ;
	    RECT 199.8000 173.8000 200.2000 174.2000 ;
	    RECT 92.6000 165.8000 93.0000 166.2000 ;
	    RECT 199.8000 163.2000 200.1000 173.8000 ;
	    RECT 200.6000 172.8000 201.0000 173.2000 ;
	    RECT 200.6000 169.2000 200.9000 172.8000 ;
	    RECT 215.8000 171.8000 216.2000 172.2000 ;
	    RECT 215.8000 170.2000 216.1000 171.8000 ;
	    RECT 219.0000 171.2000 219.3000 174.8000 ;
	    RECT 223.0000 174.2000 223.3000 174.8000 ;
	    RECT 223.0000 173.8000 223.4000 174.2000 ;
	    RECT 219.0000 170.8000 219.4000 171.2000 ;
	    RECT 214.2000 170.1000 214.6000 170.2000 ;
	    RECT 215.0000 170.1000 215.4000 170.2000 ;
	    RECT 214.2000 169.8000 215.4000 170.1000 ;
	    RECT 215.8000 169.8000 216.2000 170.2000 ;
	    RECT 221.4000 170.1000 221.8000 170.2000 ;
	    RECT 222.2000 170.1000 222.6000 170.2000 ;
	    RECT 221.4000 169.8000 222.6000 170.1000 ;
	    RECT 200.6000 168.8000 201.0000 169.2000 ;
	    RECT 244.6000 168.8000 245.0000 169.2000 ;
	    RECT 257.4000 168.8000 257.8000 169.2000 ;
	    RECT 199.8000 162.8000 200.2000 163.2000 ;
	    RECT 190.2000 161.8000 190.6000 162.2000 ;
	    RECT 29.4000 156.8000 29.8000 157.2000 ;
	    RECT 3.8000 155.8000 4.2000 156.2000 ;
	    RECT 14.2000 155.8000 14.6000 156.2000 ;
	    RECT 3.8000 146.2000 4.1000 155.8000 ;
	    RECT 29.4000 148.2000 29.7000 156.8000 ;
	    RECT 50.2000 154.8000 50.6000 155.2000 ;
	    RECT 29.4000 147.8000 29.8000 148.2000 ;
	    RECT 3.8000 145.8000 4.2000 146.2000 ;
	    RECT 39.0000 139.8000 39.4000 140.2000 ;
	    RECT 38.2000 138.8000 38.6000 139.2000 ;
	    RECT 19.0000 135.8000 19.4000 136.2000 ;
	    RECT 27.0000 135.8000 27.4000 136.2000 ;
	    RECT 19.0000 126.2000 19.3000 135.8000 ;
	    RECT 19.0000 125.8000 19.4000 126.2000 ;
	    RECT 27.0000 124.2000 27.3000 135.8000 ;
	    RECT 27.0000 123.8000 27.4000 124.2000 ;
	    RECT 17.4000 113.8000 17.8000 114.2000 ;
	    RECT 31.0000 113.8000 31.4000 114.2000 ;
	    RECT 10.2000 106.1000 10.6000 106.2000 ;
	    RECT 9.4000 105.8000 10.6000 106.1000 ;
	    RECT 8.6000 77.8000 9.0000 78.2000 ;
	    RECT 8.6000 77.2000 8.9000 77.8000 ;
	    RECT 8.6000 76.8000 9.0000 77.2000 ;
	    RECT 5.4000 75.8000 5.8000 76.2000 ;
	    RECT 5.4000 75.2000 5.7000 75.8000 ;
	    RECT 9.4000 75.2000 9.7000 105.8000 ;
	    RECT 14.2000 104.1000 14.6000 104.2000 ;
	    RECT 13.4000 103.8000 14.6000 104.1000 ;
	    RECT 11.8000 77.1000 12.2000 77.2000 ;
	    RECT 12.6000 77.1000 13.0000 77.2000 ;
	    RECT 11.8000 76.8000 13.0000 77.1000 ;
	    RECT 5.4000 74.8000 5.8000 75.2000 ;
	    RECT 9.4000 74.8000 9.8000 75.2000 ;
	    RECT 13.4000 72.2000 13.7000 103.8000 ;
	    RECT 17.4000 72.2000 17.7000 113.8000 ;
	    RECT 27.0000 113.1000 27.4000 113.2000 ;
	    RECT 26.2000 112.8000 27.4000 113.1000 ;
	    RECT 25.4000 94.8000 25.8000 95.2000 ;
	    RECT 22.2000 93.8000 22.6000 94.2000 ;
	    RECT 18.2000 77.8000 18.6000 78.2000 ;
	    RECT 13.4000 71.8000 13.8000 72.2000 ;
	    RECT 17.4000 71.8000 17.8000 72.2000 ;
	    RECT 18.2000 68.2000 18.5000 77.8000 ;
	    RECT 22.2000 71.2000 22.5000 93.8000 ;
	    RECT 23.0000 76.1000 23.4000 76.2000 ;
	    RECT 23.8000 76.1000 24.2000 76.2000 ;
	    RECT 23.0000 75.8000 24.2000 76.1000 ;
	    RECT 24.6000 74.8000 25.0000 75.2000 ;
	    RECT 24.6000 74.2000 24.9000 74.8000 ;
	    RECT 24.6000 73.8000 25.0000 74.2000 ;
	    RECT 23.0000 71.8000 23.4000 72.2000 ;
	    RECT 22.2000 70.8000 22.6000 71.2000 ;
	    RECT 23.0000 68.2000 23.3000 71.8000 ;
	    RECT 25.4000 69.2000 25.7000 94.8000 ;
	    RECT 26.2000 73.2000 26.5000 112.8000 ;
	    RECT 30.2000 88.8000 30.6000 89.2000 ;
	    RECT 27.0000 87.8000 27.4000 88.2000 ;
	    RECT 27.0000 75.2000 27.3000 87.8000 ;
	    RECT 30.2000 78.2000 30.5000 88.8000 ;
	    RECT 30.2000 77.8000 30.6000 78.2000 ;
	    RECT 27.0000 74.8000 27.4000 75.2000 ;
	    RECT 27.8000 75.1000 28.2000 75.2000 ;
	    RECT 28.6000 75.1000 29.0000 75.2000 ;
	    RECT 27.8000 74.8000 29.0000 75.1000 ;
	    RECT 26.2000 72.8000 26.6000 73.2000 ;
	    RECT 31.0000 71.2000 31.3000 113.8000 ;
	    RECT 31.0000 70.8000 31.4000 71.2000 ;
	    RECT 25.4000 68.8000 25.8000 69.2000 ;
	    RECT 18.2000 67.8000 18.6000 68.2000 ;
	    RECT 23.0000 67.8000 23.4000 68.2000 ;
	    RECT 8.6000 66.8000 9.0000 67.2000 ;
	    RECT 22.2000 66.8000 22.6000 67.2000 ;
	    RECT 8.6000 64.2000 8.9000 66.8000 ;
	    RECT 20.6000 65.8000 21.0000 66.2000 ;
	    RECT 8.6000 63.8000 9.0000 64.2000 ;
	    RECT 20.6000 56.2000 20.9000 65.8000 ;
	    RECT 20.6000 55.8000 21.0000 56.2000 ;
	    RECT 15.8000 35.1000 16.2000 35.2000 ;
	    RECT 15.0000 34.8000 16.2000 35.1000 ;
	    RECT 15.0000 34.2000 15.3000 34.8000 ;
	    RECT 15.0000 33.8000 15.4000 34.2000 ;
	    RECT 20.6000 30.2000 20.9000 55.8000 ;
	    RECT 20.6000 29.8000 21.0000 30.2000 ;
	    RECT 22.2000 28.2000 22.5000 66.8000 ;
	    RECT 31.8000 64.8000 32.2000 65.2000 ;
	    RECT 31.8000 45.2000 32.1000 64.8000 ;
	    RECT 32.6000 53.8000 33.0000 54.2000 ;
	    RECT 36.6000 54.1000 37.0000 54.2000 ;
	    RECT 37.4000 54.1000 37.8000 54.2000 ;
	    RECT 36.6000 53.8000 37.8000 54.1000 ;
	    RECT 31.8000 44.8000 32.2000 45.2000 ;
	    RECT 32.6000 35.2000 32.9000 53.8000 ;
	    RECT 32.6000 34.8000 33.0000 35.2000 ;
	    RECT 22.2000 27.8000 22.6000 28.2000 ;
	    RECT 38.2000 7.2000 38.5000 138.8000 ;
	    RECT 39.0000 132.2000 39.3000 139.8000 ;
	    RECT 50.2000 139.2000 50.5000 154.8000 ;
	    RECT 135.0000 153.8000 135.4000 154.2000 ;
	    RECT 179.8000 153.8000 180.2000 154.2000 ;
	    RECT 50.2000 138.8000 50.6000 139.2000 ;
	    RECT 117.4000 134.8000 117.8000 135.2000 ;
	    RECT 117.4000 133.2000 117.7000 134.8000 ;
	    RECT 117.4000 132.8000 117.8000 133.2000 ;
	    RECT 39.0000 131.8000 39.4000 132.2000 ;
	    RECT 88.6000 130.8000 89.0000 131.2000 ;
	    RECT 75.0000 114.8000 75.4000 115.2000 ;
	    RECT 63.0000 111.1000 63.4000 111.2000 ;
	    RECT 63.0000 110.8000 64.1000 111.1000 ;
	    RECT 50.2000 95.8000 50.6000 96.2000 ;
	    RECT 50.2000 95.2000 50.5000 95.8000 ;
	    RECT 49.4000 94.8000 49.8000 95.2000 ;
	    RECT 50.2000 94.8000 50.6000 95.2000 ;
	    RECT 49.4000 84.2000 49.7000 94.8000 ;
	    RECT 55.8000 92.8000 56.2000 93.2000 ;
	    RECT 60.6000 93.1000 61.0000 93.2000 ;
	    RECT 59.8000 92.8000 61.0000 93.1000 ;
	    RECT 49.4000 83.8000 49.8000 84.2000 ;
	    RECT 55.8000 79.2000 56.1000 92.8000 ;
	    RECT 55.8000 78.8000 56.2000 79.2000 ;
	    RECT 49.4000 74.8000 49.8000 75.2000 ;
	    RECT 49.4000 59.2000 49.7000 74.8000 ;
	    RECT 59.8000 73.2000 60.1000 92.8000 ;
	    RECT 59.8000 72.8000 60.2000 73.2000 ;
	    RECT 49.4000 58.8000 49.8000 59.2000 ;
	    RECT 63.8000 49.2000 64.1000 110.8000 ;
	    RECT 75.0000 95.2000 75.3000 114.8000 ;
	    RECT 88.6000 95.2000 88.9000 130.8000 ;
	    RECT 113.4000 127.8000 113.8000 128.2000 ;
	    RECT 126.2000 127.8000 126.6000 128.2000 ;
	    RECT 113.4000 125.2000 113.7000 127.8000 ;
	    RECT 126.2000 127.2000 126.5000 127.8000 ;
	    RECT 126.2000 126.8000 126.6000 127.2000 ;
	    RECT 113.4000 124.8000 113.8000 125.2000 ;
	    RECT 121.4000 123.8000 121.8000 124.2000 ;
	    RECT 97.4000 122.8000 97.8000 123.2000 ;
	    RECT 95.0000 119.8000 95.4000 120.2000 ;
	    RECT 90.2000 106.8000 90.6000 107.2000 ;
	    RECT 75.0000 94.8000 75.4000 95.2000 ;
	    RECT 88.6000 94.8000 89.0000 95.2000 ;
	    RECT 65.4000 82.8000 65.8000 83.2000 ;
	    RECT 65.4000 65.2000 65.7000 82.8000 ;
	    RECT 70.2000 74.1000 70.6000 74.2000 ;
	    RECT 71.0000 74.1000 71.4000 74.2000 ;
	    RECT 70.2000 73.8000 71.4000 74.1000 ;
	    RECT 88.6000 72.2000 88.9000 94.8000 ;
	    RECT 90.2000 87.2000 90.5000 106.8000 ;
	    RECT 95.0000 95.2000 95.3000 119.8000 ;
	    RECT 95.0000 94.8000 95.4000 95.2000 ;
	    RECT 90.2000 86.8000 90.6000 87.2000 ;
	    RECT 95.0000 74.2000 95.3000 94.8000 ;
	    RECT 95.0000 73.8000 95.4000 74.2000 ;
	    RECT 79.0000 71.8000 79.4000 72.2000 ;
	    RECT 88.6000 71.8000 89.0000 72.2000 ;
	    RECT 79.0000 66.2000 79.3000 71.8000 ;
	    RECT 97.4000 66.2000 97.7000 122.8000 ;
	    RECT 121.4000 121.2000 121.7000 123.8000 ;
	    RECT 121.4000 120.8000 121.8000 121.2000 ;
	    RECT 100.6000 111.8000 101.0000 112.2000 ;
	    RECT 100.6000 105.2000 100.9000 111.8000 ;
	    RECT 121.4000 105.2000 121.7000 120.8000 ;
	    RECT 133.4000 114.8000 133.8000 115.2000 ;
	    RECT 133.4000 113.2000 133.7000 114.8000 ;
	    RECT 133.4000 112.8000 133.8000 113.2000 ;
	    RECT 100.6000 104.8000 101.0000 105.2000 ;
	    RECT 121.4000 104.8000 121.8000 105.2000 ;
	    RECT 98.2000 98.8000 98.6000 99.2000 ;
	    RECT 98.2000 80.2000 98.5000 98.8000 ;
	    RECT 103.8000 96.8000 104.2000 97.2000 ;
	    RECT 98.2000 79.8000 98.6000 80.2000 ;
	    RECT 101.4000 74.1000 101.8000 74.2000 ;
	    RECT 102.2000 74.1000 102.6000 74.2000 ;
	    RECT 101.4000 73.8000 102.6000 74.1000 ;
	    RECT 103.8000 73.2000 104.1000 96.8000 ;
	    RECT 103.8000 72.8000 104.2000 73.2000 ;
	    RECT 104.6000 72.8000 105.0000 73.2000 ;
	    RECT 79.0000 65.8000 79.4000 66.2000 ;
	    RECT 97.4000 65.8000 97.8000 66.2000 ;
	    RECT 65.4000 64.8000 65.8000 65.2000 ;
	    RECT 71.0000 64.1000 71.4000 64.2000 ;
	    RECT 71.0000 63.8000 72.1000 64.1000 ;
	    RECT 69.4000 50.8000 69.8000 51.2000 ;
	    RECT 63.8000 48.8000 64.2000 49.2000 ;
	    RECT 67.8000 16.8000 68.2000 17.2000 ;
	    RECT 67.0000 14.8000 67.4000 15.2000 ;
	    RECT 67.0000 14.2000 67.3000 14.8000 ;
	    RECT 67.8000 14.2000 68.1000 16.8000 ;
	    RECT 67.0000 13.8000 67.4000 14.2000 ;
	    RECT 67.8000 13.8000 68.2000 14.2000 ;
	    RECT 38.2000 6.8000 38.6000 7.2000 ;
	    RECT 69.4000 7.1000 69.7000 50.8000 ;
	    RECT 71.8000 50.2000 72.1000 63.8000 ;
	    RECT 104.6000 58.2000 104.9000 72.8000 ;
	    RECT 135.0000 68.2000 135.3000 153.8000 ;
	    RECT 179.8000 153.2000 180.1000 153.8000 ;
	    RECT 179.8000 152.8000 180.2000 153.2000 ;
	    RECT 188.6000 147.1000 189.0000 147.2000 ;
	    RECT 189.4000 147.1000 189.8000 147.2000 ;
	    RECT 188.6000 146.8000 189.8000 147.1000 ;
	    RECT 141.4000 145.8000 141.8000 146.2000 ;
	    RECT 142.2000 146.1000 142.6000 146.2000 ;
	    RECT 142.2000 145.8000 143.3000 146.1000 ;
	    RECT 140.6000 123.8000 141.0000 124.2000 ;
	    RECT 135.8000 117.8000 136.2000 118.2000 ;
	    RECT 135.8000 114.1000 136.1000 117.8000 ;
	    RECT 136.6000 114.1000 137.0000 114.2000 ;
	    RECT 135.8000 113.8000 137.0000 114.1000 ;
	    RECT 138.2000 109.8000 138.6000 110.2000 ;
	    RECT 138.2000 94.2000 138.5000 109.8000 ;
	    RECT 140.6000 96.2000 140.9000 123.8000 ;
	    RECT 141.4000 105.2000 141.7000 145.8000 ;
	    RECT 141.4000 104.8000 141.8000 105.2000 ;
	    RECT 140.6000 95.8000 141.0000 96.2000 ;
	    RECT 138.2000 93.8000 138.6000 94.2000 ;
	    RECT 143.0000 93.2000 143.3000 145.8000 ;
	    RECT 190.2000 144.2000 190.5000 161.8000 ;
	    RECT 199.8000 151.2000 200.1000 162.8000 ;
	    RECT 199.8000 150.8000 200.2000 151.2000 ;
	    RECT 190.2000 143.8000 190.6000 144.2000 ;
	    RECT 200.6000 142.2000 200.9000 168.8000 ;
	    RECT 232.6000 166.8000 233.0000 167.2000 ;
	    RECT 215.8000 147.8000 216.2000 148.2000 ;
	    RECT 212.6000 147.1000 213.0000 147.2000 ;
	    RECT 213.4000 147.1000 213.8000 147.2000 ;
	    RECT 212.6000 146.8000 213.8000 147.1000 ;
	    RECT 200.6000 141.8000 201.0000 142.2000 ;
	    RECT 175.8000 140.1000 176.2000 140.2000 ;
	    RECT 175.8000 139.8000 176.9000 140.1000 ;
	    RECT 176.6000 134.2000 176.9000 139.8000 ;
	    RECT 200.6000 138.8000 201.0000 139.2000 ;
	    RECT 177.4000 136.8000 177.8000 137.2000 ;
	    RECT 176.6000 133.8000 177.0000 134.2000 ;
	    RECT 174.2000 127.8000 174.6000 128.2000 ;
	    RECT 145.4000 127.1000 145.8000 127.2000 ;
	    RECT 146.2000 127.1000 146.6000 127.2000 ;
	    RECT 145.4000 126.8000 146.6000 127.1000 ;
	    RECT 174.2000 107.2000 174.5000 127.8000 ;
	    RECT 174.2000 106.8000 174.6000 107.2000 ;
	    RECT 177.4000 107.1000 177.7000 136.8000 ;
	    RECT 180.6000 133.8000 181.0000 134.2000 ;
	    RECT 180.6000 115.1000 180.9000 133.8000 ;
	    RECT 186.2000 116.8000 186.6000 117.2000 ;
	    RECT 194.2000 116.8000 194.6000 117.2000 ;
	    RECT 181.4000 115.1000 181.8000 115.2000 ;
	    RECT 180.6000 114.8000 181.8000 115.1000 ;
	    RECT 178.2000 107.1000 178.6000 107.2000 ;
	    RECT 177.4000 106.8000 178.6000 107.1000 ;
	    RECT 182.2000 106.8000 182.6000 107.2000 ;
	    RECT 170.2000 105.8000 170.6000 106.2000 ;
	    RECT 168.6000 95.8000 169.0000 96.2000 ;
	    RECT 143.0000 92.8000 143.4000 93.2000 ;
	    RECT 168.6000 92.2000 168.9000 95.8000 ;
	    RECT 168.6000 91.8000 169.0000 92.2000 ;
	    RECT 159.0000 88.8000 159.4000 89.2000 ;
	    RECT 140.6000 81.8000 141.0000 82.2000 ;
	    RECT 135.0000 67.8000 135.4000 68.2000 ;
	    RECT 111.0000 62.8000 111.4000 63.2000 ;
	    RECT 104.6000 57.8000 105.0000 58.2000 ;
	    RECT 82.2000 52.8000 82.6000 53.2000 ;
	    RECT 71.8000 49.8000 72.2000 50.2000 ;
	    RECT 82.2000 41.2000 82.5000 52.8000 ;
	    RECT 111.0000 44.2000 111.3000 62.8000 ;
	    RECT 132.6000 56.8000 133.0000 57.2000 ;
	    RECT 130.2000 54.8000 130.6000 55.2000 ;
	    RECT 124.6000 52.8000 125.0000 53.2000 ;
	    RECT 121.4000 48.8000 121.8000 49.2000 ;
	    RECT 111.0000 43.8000 111.4000 44.2000 ;
	    RECT 82.2000 40.8000 82.6000 41.2000 ;
	    RECT 106.2000 38.8000 106.6000 39.2000 ;
	    RECT 99.0000 33.8000 99.4000 34.2000 ;
	    RECT 99.0000 21.2000 99.3000 33.8000 ;
	    RECT 99.0000 20.8000 99.4000 21.2000 ;
	    RECT 71.0000 15.1000 71.4000 15.2000 ;
	    RECT 71.8000 15.1000 72.2000 15.2000 ;
	    RECT 71.0000 14.8000 72.2000 15.1000 ;
	    RECT 91.8000 15.1000 92.2000 15.2000 ;
	    RECT 92.6000 15.1000 93.0000 15.2000 ;
	    RECT 91.8000 14.8000 93.0000 15.1000 ;
	    RECT 88.6000 14.1000 89.0000 14.2000 ;
	    RECT 89.4000 14.1000 89.8000 14.2000 ;
	    RECT 88.6000 13.8000 89.8000 14.1000 ;
	    RECT 102.2000 13.8000 102.6000 14.2000 ;
	    RECT 102.2000 13.2000 102.5000 13.8000 ;
	    RECT 95.0000 12.8000 95.4000 13.2000 ;
	    RECT 100.6000 13.1000 101.0000 13.2000 ;
	    RECT 101.4000 13.1000 101.8000 13.2000 ;
	    RECT 100.6000 12.8000 101.8000 13.1000 ;
	    RECT 102.2000 12.8000 102.6000 13.2000 ;
	    RECT 95.0000 12.2000 95.3000 12.8000 ;
	    RECT 95.0000 11.8000 95.4000 12.2000 ;
	    RECT 105.4000 11.1000 105.8000 11.2000 ;
	    RECT 104.6000 10.8000 105.8000 11.1000 ;
	    RECT 104.6000 9.2000 104.9000 10.8000 ;
	    RECT 106.2000 9.2000 106.5000 38.8000 ;
	    RECT 111.0000 38.2000 111.3000 43.8000 ;
	    RECT 111.0000 37.8000 111.4000 38.2000 ;
	    RECT 119.8000 38.1000 120.2000 38.2000 ;
	    RECT 119.0000 37.8000 120.2000 38.1000 ;
	    RECT 119.0000 28.2000 119.3000 37.8000 ;
	    RECT 121.4000 29.2000 121.7000 48.8000 ;
	    RECT 123.0000 35.8000 123.4000 36.2000 ;
	    RECT 121.4000 28.8000 121.8000 29.2000 ;
	    RECT 119.0000 27.8000 119.4000 28.2000 ;
	    RECT 110.2000 25.1000 110.6000 25.2000 ;
	    RECT 111.0000 25.1000 111.4000 25.2000 ;
	    RECT 110.2000 24.8000 111.4000 25.1000 ;
	    RECT 113.4000 15.8000 113.8000 16.2000 ;
	    RECT 113.4000 14.2000 113.7000 15.8000 ;
	    RECT 123.0000 15.2000 123.3000 35.8000 ;
	    RECT 123.8000 34.1000 124.2000 34.2000 ;
	    RECT 124.6000 34.1000 124.9000 52.8000 ;
	    RECT 129.4000 45.1000 129.8000 45.2000 ;
	    RECT 130.2000 45.1000 130.5000 54.8000 ;
	    RECT 132.6000 54.2000 132.9000 56.8000 ;
	    RECT 135.0000 54.2000 135.3000 67.8000 ;
	    RECT 132.6000 53.8000 133.0000 54.2000 ;
	    RECT 135.0000 53.8000 135.4000 54.2000 ;
	    RECT 129.4000 44.8000 130.5000 45.1000 ;
	    RECT 129.4000 36.2000 129.7000 44.8000 ;
	    RECT 140.6000 36.2000 140.9000 81.8000 ;
	    RECT 159.0000 76.2000 159.3000 88.8000 ;
	    RECT 170.2000 87.2000 170.5000 105.8000 ;
	    RECT 170.2000 86.8000 170.6000 87.2000 ;
	    RECT 178.2000 84.2000 178.5000 106.8000 ;
	    RECT 182.2000 98.2000 182.5000 106.8000 ;
	    RECT 182.2000 97.8000 182.6000 98.2000 ;
	    RECT 179.8000 92.8000 180.2000 93.2000 ;
	    RECT 178.2000 83.8000 178.6000 84.2000 ;
	    RECT 159.0000 75.8000 159.4000 76.2000 ;
	    RECT 179.8000 73.2000 180.1000 92.8000 ;
	    RECT 179.8000 72.8000 180.2000 73.2000 ;
	    RECT 142.2000 61.8000 142.6000 62.2000 ;
	    RECT 129.4000 35.8000 129.8000 36.2000 ;
	    RECT 140.6000 35.8000 141.0000 36.2000 ;
	    RECT 123.8000 33.8000 124.9000 34.1000 ;
	    RECT 142.2000 33.2000 142.5000 61.8000 ;
	    RECT 181.4000 59.8000 181.8000 60.2000 ;
	    RECT 176.6000 52.8000 177.0000 53.2000 ;
	    RECT 157.4000 41.8000 157.8000 42.2000 ;
	    RECT 142.2000 32.8000 142.6000 33.2000 ;
	    RECT 127.8000 31.8000 128.2000 32.2000 ;
	    RECT 127.8000 26.2000 128.1000 31.8000 ;
	    RECT 127.8000 25.8000 128.2000 26.2000 ;
	    RECT 135.8000 25.1000 136.2000 25.2000 ;
	    RECT 136.6000 25.1000 137.0000 25.2000 ;
	    RECT 135.8000 24.8000 137.0000 25.1000 ;
	    RECT 157.4000 15.2000 157.7000 41.8000 ;
	    RECT 176.6000 33.2000 176.9000 52.8000 ;
	    RECT 181.4000 35.2000 181.7000 59.8000 ;
	    RECT 181.4000 34.8000 181.8000 35.2000 ;
	    RECT 176.6000 32.8000 177.0000 33.2000 ;
	    RECT 185.4000 31.1000 185.8000 31.2000 ;
	    RECT 186.2000 31.1000 186.5000 116.8000 ;
	    RECT 189.4000 110.8000 189.8000 111.2000 ;
	    RECT 189.4000 100.2000 189.7000 110.8000 ;
	    RECT 189.4000 99.8000 189.8000 100.2000 ;
	    RECT 187.8000 89.1000 188.2000 89.2000 ;
	    RECT 188.6000 89.1000 189.0000 89.2000 ;
	    RECT 187.8000 88.8000 189.0000 89.1000 ;
	    RECT 188.6000 74.1000 189.0000 74.2000 ;
	    RECT 189.4000 74.1000 189.7000 99.8000 ;
	    RECT 190.2000 91.8000 190.6000 92.2000 ;
	    RECT 190.2000 89.1000 190.5000 91.8000 ;
	    RECT 191.0000 89.1000 191.4000 89.2000 ;
	    RECT 190.2000 88.8000 191.4000 89.1000 ;
	    RECT 194.2000 76.2000 194.5000 116.8000 ;
	    RECT 200.6000 114.2000 200.9000 138.8000 ;
	    RECT 207.0000 132.8000 207.4000 133.2000 ;
	    RECT 205.4000 131.8000 205.8000 132.2000 ;
	    RECT 205.4000 126.2000 205.7000 131.8000 ;
	    RECT 205.4000 125.8000 205.8000 126.2000 ;
	    RECT 207.0000 114.2000 207.3000 132.8000 ;
	    RECT 195.8000 113.8000 196.2000 114.2000 ;
	    RECT 200.6000 113.8000 201.0000 114.2000 ;
	    RECT 207.0000 113.8000 207.4000 114.2000 ;
	    RECT 195.8000 88.2000 196.1000 113.8000 ;
	    RECT 200.6000 110.2000 200.9000 113.8000 ;
	    RECT 208.6000 112.8000 209.0000 113.2000 ;
	    RECT 200.6000 109.8000 201.0000 110.2000 ;
	    RECT 201.4000 109.8000 201.8000 110.2000 ;
	    RECT 200.6000 108.8000 201.0000 109.2000 ;
	    RECT 200.6000 93.2000 200.9000 108.8000 ;
	    RECT 201.4000 108.2000 201.7000 109.8000 ;
	    RECT 201.4000 107.8000 201.8000 108.2000 ;
	    RECT 200.6000 92.8000 201.0000 93.2000 ;
	    RECT 195.8000 87.8000 196.2000 88.2000 ;
	    RECT 195.8000 85.8000 196.2000 86.2000 ;
	    RECT 194.2000 75.8000 194.6000 76.2000 ;
	    RECT 195.8000 75.2000 196.1000 85.8000 ;
	    RECT 195.8000 74.8000 196.2000 75.2000 ;
	    RECT 188.6000 73.8000 189.7000 74.1000 ;
	    RECT 200.6000 68.2000 200.9000 92.8000 ;
	    RECT 206.2000 87.1000 206.6000 87.2000 ;
	    RECT 207.0000 87.1000 207.4000 87.2000 ;
	    RECT 206.2000 86.8000 207.4000 87.1000 ;
	    RECT 207.8000 85.1000 208.2000 85.2000 ;
	    RECT 208.6000 85.1000 208.9000 112.8000 ;
	    RECT 215.8000 94.2000 216.1000 147.8000 ;
	    RECT 231.8000 145.8000 232.2000 146.2000 ;
	    RECT 224.6000 144.8000 225.0000 145.2000 ;
	    RECT 224.6000 139.2000 224.9000 144.8000 ;
	    RECT 224.6000 138.8000 225.0000 139.2000 ;
	    RECT 225.4000 134.8000 225.8000 135.2000 ;
	    RECT 225.4000 133.2000 225.7000 134.8000 ;
	    RECT 230.2000 133.8000 230.6000 134.2000 ;
	    RECT 225.4000 132.8000 225.8000 133.2000 ;
	    RECT 230.2000 131.2000 230.5000 133.8000 ;
	    RECT 231.8000 131.2000 232.1000 145.8000 ;
	    RECT 230.2000 130.8000 230.6000 131.2000 ;
	    RECT 231.8000 130.8000 232.2000 131.2000 ;
	    RECT 217.4000 127.8000 217.8000 128.2000 ;
	    RECT 217.4000 123.2000 217.7000 127.8000 ;
	    RECT 223.8000 126.8000 224.2000 127.2000 ;
	    RECT 221.4000 123.8000 221.8000 124.2000 ;
	    RECT 223.0000 124.1000 223.4000 124.2000 ;
	    RECT 222.2000 123.8000 223.4000 124.1000 ;
	    RECT 217.4000 122.8000 217.8000 123.2000 ;
	    RECT 219.8000 105.8000 220.2000 106.2000 ;
	    RECT 215.8000 93.8000 216.2000 94.2000 ;
	    RECT 207.8000 84.8000 208.9000 85.1000 ;
	    RECT 209.4000 90.8000 209.8000 91.2000 ;
	    RECT 205.4000 83.8000 205.8000 84.2000 ;
	    RECT 205.4000 71.2000 205.7000 83.8000 ;
	    RECT 209.4000 74.2000 209.7000 90.8000 ;
	    RECT 215.0000 87.8000 215.4000 88.2000 ;
	    RECT 207.0000 74.1000 207.4000 74.2000 ;
	    RECT 207.8000 74.1000 208.2000 74.2000 ;
	    RECT 207.0000 73.8000 208.2000 74.1000 ;
	    RECT 209.4000 73.8000 209.8000 74.2000 ;
	    RECT 205.4000 70.8000 205.8000 71.2000 ;
	    RECT 204.6000 68.8000 205.0000 69.2000 ;
	    RECT 200.6000 67.8000 201.0000 68.2000 ;
	    RECT 204.6000 55.2000 204.9000 68.8000 ;
	    RECT 205.4000 67.2000 205.7000 70.8000 ;
	    RECT 215.0000 67.2000 215.3000 87.8000 ;
	    RECT 219.8000 85.2000 220.1000 105.8000 ;
	    RECT 219.8000 84.8000 220.2000 85.2000 ;
	    RECT 221.4000 72.2000 221.7000 123.8000 ;
	    RECT 222.2000 107.2000 222.5000 123.8000 ;
	    RECT 222.2000 106.8000 222.6000 107.2000 ;
	    RECT 223.8000 104.2000 224.1000 126.8000 ;
	    RECT 230.2000 120.2000 230.5000 130.8000 ;
	    RECT 230.2000 119.8000 230.6000 120.2000 ;
	    RECT 230.2000 114.1000 230.6000 114.2000 ;
	    RECT 231.0000 114.1000 231.4000 114.2000 ;
	    RECT 230.2000 113.8000 231.4000 114.1000 ;
	    RECT 230.2000 106.8000 230.6000 107.2000 ;
	    RECT 223.8000 103.8000 224.2000 104.2000 ;
	    RECT 223.8000 88.8000 224.2000 89.2000 ;
	    RECT 223.8000 86.2000 224.1000 88.8000 ;
	    RECT 225.4000 86.8000 225.8000 87.2000 ;
	    RECT 225.4000 86.2000 225.7000 86.8000 ;
	    RECT 222.2000 86.1000 222.6000 86.2000 ;
	    RECT 223.0000 86.1000 223.4000 86.2000 ;
	    RECT 222.2000 85.8000 223.4000 86.1000 ;
	    RECT 223.8000 85.8000 224.2000 86.2000 ;
	    RECT 225.4000 85.8000 225.8000 86.2000 ;
	    RECT 229.4000 76.8000 229.8000 77.2000 ;
	    RECT 228.6000 75.8000 229.0000 76.2000 ;
	    RECT 227.8000 72.8000 228.2000 73.2000 ;
	    RECT 221.4000 71.8000 221.8000 72.2000 ;
	    RECT 227.0000 70.8000 227.4000 71.2000 ;
	    RECT 205.4000 66.8000 205.8000 67.2000 ;
	    RECT 215.0000 66.8000 215.4000 67.2000 ;
	    RECT 204.6000 54.8000 205.0000 55.2000 ;
	    RECT 227.0000 51.2000 227.3000 70.8000 ;
	    RECT 227.0000 50.8000 227.4000 51.2000 ;
	    RECT 227.8000 50.2000 228.1000 72.8000 ;
	    RECT 228.6000 65.2000 228.9000 75.8000 ;
	    RECT 229.4000 65.2000 229.7000 76.8000 ;
	    RECT 230.2000 72.2000 230.5000 106.8000 ;
	    RECT 231.8000 106.2000 232.1000 130.8000 ;
	    RECT 232.6000 122.2000 232.9000 166.8000 ;
	    RECT 244.6000 166.2000 244.9000 168.8000 ;
	    RECT 244.6000 165.8000 245.0000 166.2000 ;
	    RECT 246.2000 166.1000 246.6000 166.2000 ;
	    RECT 247.0000 166.1000 247.4000 166.2000 ;
	    RECT 246.2000 165.8000 247.4000 166.1000 ;
	    RECT 236.6000 165.1000 237.0000 165.2000 ;
	    RECT 237.4000 165.1000 237.8000 165.2000 ;
	    RECT 236.6000 164.8000 237.8000 165.1000 ;
	    RECT 238.2000 164.8000 238.6000 165.2000 ;
	    RECT 239.8000 165.1000 240.2000 165.2000 ;
	    RECT 240.6000 165.1000 241.0000 165.2000 ;
	    RECT 239.8000 164.8000 241.0000 165.1000 ;
	    RECT 233.4000 158.8000 233.8000 159.2000 ;
	    RECT 232.6000 121.8000 233.0000 122.2000 ;
	    RECT 231.8000 105.8000 232.2000 106.2000 ;
	    RECT 233.4000 87.2000 233.7000 158.8000 ;
	    RECT 238.2000 151.2000 238.5000 164.8000 ;
	    RECT 241.4000 152.8000 241.8000 153.2000 ;
	    RECT 251.0000 152.8000 251.4000 153.2000 ;
	    RECT 254.2000 152.8000 254.6000 153.2000 ;
	    RECT 238.2000 150.8000 238.6000 151.2000 ;
	    RECT 241.4000 136.2000 241.7000 152.8000 ;
	    RECT 242.2000 147.1000 242.6000 147.2000 ;
	    RECT 242.2000 146.8000 243.3000 147.1000 ;
	    RECT 241.4000 135.8000 241.8000 136.2000 ;
	    RECT 242.2000 134.8000 242.6000 135.2000 ;
	    RECT 240.6000 125.8000 241.0000 126.2000 ;
	    RECT 235.0000 124.1000 235.4000 124.2000 ;
	    RECT 235.0000 123.8000 236.1000 124.1000 ;
	    RECT 235.8000 100.2000 236.1000 123.8000 ;
	    RECT 240.6000 117.2000 240.9000 125.8000 ;
	    RECT 239.0000 116.8000 239.4000 117.2000 ;
	    RECT 240.6000 116.8000 241.0000 117.2000 ;
	    RECT 235.8000 99.8000 236.2000 100.2000 ;
	    RECT 239.0000 97.2000 239.3000 116.8000 ;
	    RECT 239.0000 96.8000 239.4000 97.2000 ;
	    RECT 235.0000 95.8000 235.4000 96.2000 ;
	    RECT 233.4000 86.8000 233.8000 87.2000 ;
	    RECT 230.2000 71.8000 230.6000 72.2000 ;
	    RECT 228.6000 64.8000 229.0000 65.2000 ;
	    RECT 229.4000 64.8000 229.8000 65.2000 ;
	    RECT 233.4000 55.2000 233.7000 86.8000 ;
	    RECT 235.0000 84.2000 235.3000 95.8000 ;
	    RECT 240.6000 95.2000 240.9000 116.8000 ;
	    RECT 242.2000 116.2000 242.5000 134.8000 ;
	    RECT 243.0000 130.2000 243.3000 146.8000 ;
	    RECT 251.0000 146.2000 251.3000 152.8000 ;
	    RECT 254.2000 152.2000 254.5000 152.8000 ;
	    RECT 254.2000 151.8000 254.6000 152.2000 ;
	    RECT 251.0000 145.8000 251.4000 146.2000 ;
	    RECT 243.0000 129.8000 243.4000 130.2000 ;
	    RECT 243.0000 119.2000 243.3000 129.8000 ;
	    RECT 243.0000 118.8000 243.4000 119.2000 ;
	    RECT 242.2000 115.8000 242.6000 116.2000 ;
	    RECT 250.2000 114.1000 250.6000 114.2000 ;
	    RECT 251.0000 114.1000 251.4000 114.2000 ;
	    RECT 250.2000 113.8000 251.4000 114.1000 ;
	    RECT 243.8000 109.8000 244.2000 110.2000 ;
	    RECT 243.8000 102.2000 244.1000 109.8000 ;
	    RECT 243.8000 101.8000 244.2000 102.2000 ;
	    RECT 247.8000 101.8000 248.2000 102.2000 ;
	    RECT 240.6000 94.8000 241.0000 95.2000 ;
	    RECT 237.4000 92.1000 237.8000 92.2000 ;
	    RECT 238.2000 92.1000 238.6000 92.2000 ;
	    RECT 237.4000 91.8000 238.6000 92.1000 ;
	    RECT 235.0000 83.8000 235.4000 84.2000 ;
	    RECT 243.8000 73.8000 244.2000 74.2000 ;
	    RECT 243.8000 72.2000 244.1000 73.8000 ;
	    RECT 243.8000 71.8000 244.2000 72.2000 ;
	    RECT 238.2000 66.8000 238.6000 67.2000 ;
	    RECT 238.2000 66.2000 238.5000 66.8000 ;
	    RECT 247.8000 66.2000 248.1000 101.8000 ;
	    RECT 253.4000 94.8000 253.8000 95.2000 ;
	    RECT 251.8000 88.8000 252.2000 89.2000 ;
	    RECT 252.6000 88.8000 253.0000 89.2000 ;
	    RECT 238.2000 65.8000 238.6000 66.2000 ;
	    RECT 247.8000 65.8000 248.2000 66.2000 ;
	    RECT 233.4000 54.8000 233.8000 55.2000 ;
	    RECT 227.8000 49.8000 228.2000 50.2000 ;
	    RECT 233.4000 39.2000 233.7000 54.8000 ;
	    RECT 233.4000 38.8000 233.8000 39.2000 ;
	    RECT 224.6000 34.8000 225.0000 35.2000 ;
	    RECT 185.4000 30.8000 186.5000 31.1000 ;
	    RECT 220.6000 33.8000 221.0000 34.2000 ;
	    RECT 220.6000 31.2000 220.9000 33.8000 ;
	    RECT 224.6000 32.2000 224.9000 34.8000 ;
	    RECT 224.6000 31.8000 225.0000 32.2000 ;
	    RECT 220.6000 30.8000 221.0000 31.2000 ;
	    RECT 207.0000 16.8000 207.4000 17.2000 ;
	    RECT 122.2000 14.8000 122.6000 15.2000 ;
	    RECT 123.0000 14.8000 123.4000 15.2000 ;
	    RECT 124.6000 14.8000 125.0000 15.2000 ;
	    RECT 157.4000 14.8000 157.8000 15.2000 ;
	    RECT 113.4000 13.8000 113.8000 14.2000 ;
	    RECT 119.8000 13.8000 120.2000 14.2000 ;
	    RECT 119.8000 13.2000 120.1000 13.8000 ;
	    RECT 117.4000 12.8000 117.8000 13.2000 ;
	    RECT 119.8000 12.8000 120.2000 13.2000 ;
	    RECT 73.4000 8.8000 73.8000 9.2000 ;
	    RECT 104.6000 8.8000 105.0000 9.2000 ;
	    RECT 106.2000 8.8000 106.6000 9.2000 ;
	    RECT 73.4000 7.2000 73.7000 8.8000 ;
	    RECT 117.4000 8.2000 117.7000 12.8000 ;
	    RECT 122.2000 8.2000 122.5000 14.8000 ;
	    RECT 124.6000 12.2000 124.9000 14.8000 ;
	    RECT 207.0000 13.2000 207.3000 16.8000 ;
	    RECT 233.4000 15.2000 233.7000 38.8000 ;
	    RECT 246.2000 34.8000 246.6000 35.2000 ;
	    RECT 242.2000 32.8000 242.6000 33.2000 ;
	    RECT 243.8000 32.8000 244.2000 33.2000 ;
	    RECT 237.4000 30.8000 237.8000 31.2000 ;
	    RECT 237.4000 27.2000 237.7000 30.8000 ;
	    RECT 238.2000 28.8000 238.6000 29.2000 ;
	    RECT 237.4000 26.8000 237.8000 27.2000 ;
	    RECT 238.2000 19.2000 238.5000 28.8000 ;
	    RECT 242.2000 24.2000 242.5000 32.8000 ;
	    RECT 243.8000 24.2000 244.1000 32.8000 ;
	    RECT 242.2000 23.8000 242.6000 24.2000 ;
	    RECT 243.8000 23.8000 244.2000 24.2000 ;
	    RECT 238.2000 18.8000 238.6000 19.2000 ;
	    RECT 246.2000 15.2000 246.5000 34.8000 ;
	    RECT 251.8000 30.2000 252.1000 88.8000 ;
	    RECT 252.6000 87.2000 252.9000 88.8000 ;
	    RECT 252.6000 86.8000 253.0000 87.2000 ;
	    RECT 253.4000 48.2000 253.7000 94.8000 ;
	    RECT 254.2000 93.2000 254.5000 151.8000 ;
	    RECT 257.4000 113.2000 257.7000 168.8000 ;
	    RECT 266.2000 160.8000 266.6000 161.2000 ;
	    RECT 258.2000 141.8000 258.6000 142.2000 ;
	    RECT 258.2000 138.2000 258.5000 141.8000 ;
	    RECT 258.2000 137.8000 258.6000 138.2000 ;
	    RECT 266.2000 135.2000 266.5000 160.8000 ;
	    RECT 266.2000 134.8000 266.6000 135.2000 ;
	    RECT 257.4000 112.8000 257.8000 113.2000 ;
	    RECT 266.2000 98.2000 266.5000 134.8000 ;
	    RECT 266.2000 97.8000 266.6000 98.2000 ;
	    RECT 254.2000 92.8000 254.6000 93.2000 ;
	    RECT 253.4000 47.8000 253.8000 48.2000 ;
	    RECT 252.6000 43.8000 253.0000 44.2000 ;
	    RECT 251.8000 29.8000 252.2000 30.2000 ;
	    RECT 233.4000 14.8000 233.8000 15.2000 ;
	    RECT 246.2000 14.8000 246.6000 15.2000 ;
	    RECT 252.6000 14.2000 252.9000 43.8000 ;
	    RECT 254.2000 36.2000 254.5000 92.8000 ;
	    RECT 259.0000 89.8000 259.4000 90.2000 ;
	    RECT 255.0000 86.8000 255.4000 87.2000 ;
	    RECT 255.0000 51.2000 255.3000 86.8000 ;
	    RECT 257.4000 84.8000 257.8000 85.2000 ;
	    RECT 256.6000 76.8000 257.0000 77.2000 ;
	    RECT 255.0000 50.8000 255.4000 51.2000 ;
	    RECT 254.2000 35.8000 254.6000 36.2000 ;
	    RECT 252.6000 13.8000 253.0000 14.2000 ;
	    RECT 256.6000 13.2000 256.9000 76.8000 ;
	    RECT 257.4000 22.2000 257.7000 84.8000 ;
	    RECT 259.0000 75.2000 259.3000 89.8000 ;
	    RECT 259.0000 74.8000 259.4000 75.2000 ;
	    RECT 263.8000 73.1000 264.2000 73.2000 ;
	    RECT 263.0000 72.8000 264.2000 73.1000 ;
	    RECT 259.8000 41.8000 260.2000 42.2000 ;
	    RECT 259.0000 37.8000 259.4000 38.2000 ;
	    RECT 257.4000 21.8000 257.8000 22.2000 ;
	    RECT 259.0000 14.2000 259.3000 37.8000 ;
	    RECT 259.8000 32.2000 260.1000 41.8000 ;
	    RECT 259.8000 31.8000 260.2000 32.2000 ;
	    RECT 259.0000 13.8000 259.4000 14.2000 ;
	    RECT 207.0000 12.8000 207.4000 13.2000 ;
	    RECT 256.6000 12.8000 257.0000 13.2000 ;
	    RECT 123.8000 11.8000 124.2000 12.2000 ;
	    RECT 124.6000 11.8000 125.0000 12.2000 ;
	    RECT 133.4000 12.1000 133.8000 12.2000 ;
	    RECT 134.2000 12.1000 134.6000 12.2000 ;
	    RECT 133.4000 11.8000 134.6000 12.1000 ;
	    RECT 123.8000 8.2000 124.1000 11.8000 ;
	    RECT 263.0000 11.2000 263.3000 72.8000 ;
	    RECT 266.2000 66.2000 266.5000 97.8000 ;
	    RECT 268.6000 71.8000 269.0000 72.2000 ;
	    RECT 266.2000 65.8000 266.6000 66.2000 ;
	    RECT 263.8000 48.8000 264.2000 49.2000 ;
	    RECT 263.8000 26.2000 264.1000 48.8000 ;
	    RECT 263.8000 25.8000 264.2000 26.2000 ;
	    RECT 263.0000 10.8000 263.4000 11.2000 ;
	    RECT 126.2000 8.8000 126.6000 9.2000 ;
	    RECT 117.4000 7.8000 117.8000 8.2000 ;
	    RECT 122.2000 7.8000 122.6000 8.2000 ;
	    RECT 123.8000 7.8000 124.2000 8.2000 ;
	    RECT 70.2000 7.1000 70.6000 7.2000 ;
	    RECT 69.4000 6.8000 70.6000 7.1000 ;
	    RECT 73.4000 6.8000 73.8000 7.2000 ;
	    RECT 80.6000 7.1000 81.0000 7.2000 ;
	    RECT 81.4000 7.1000 81.8000 7.2000 ;
	    RECT 80.6000 6.8000 81.8000 7.1000 ;
	    RECT 88.6000 7.1000 89.0000 7.2000 ;
	    RECT 89.4000 7.1000 89.8000 7.2000 ;
	    RECT 88.6000 6.8000 89.8000 7.1000 ;
	    RECT 99.0000 7.1000 99.4000 7.2000 ;
	    RECT 99.8000 7.1000 100.2000 7.2000 ;
	    RECT 99.0000 6.8000 100.2000 7.1000 ;
	    RECT 103.0000 7.1000 103.4000 7.2000 ;
	    RECT 103.8000 7.1000 104.2000 7.2000 ;
	    RECT 103.0000 6.8000 104.2000 7.1000 ;
	    RECT 126.2000 5.2000 126.5000 8.8000 ;
	    RECT 268.6000 8.2000 268.9000 71.8000 ;
	    RECT 131.0000 8.1000 131.4000 8.2000 ;
	    RECT 131.8000 8.1000 132.2000 8.2000 ;
	    RECT 131.0000 7.8000 132.2000 8.1000 ;
	    RECT 268.6000 7.8000 269.0000 8.2000 ;
	    RECT 126.2000 4.8000 126.6000 5.2000 ;
         LAYER metal5 ;
	    RECT 214.2000 170.1000 214.6000 170.2000 ;
	    RECT 221.4000 170.1000 221.8000 170.2000 ;
	    RECT 214.2000 169.8000 221.8000 170.1000 ;
	    RECT 244.6000 166.1000 245.0000 166.2000 ;
	    RECT 247.0000 166.1000 247.4000 166.2000 ;
	    RECT 244.6000 165.8000 247.4000 166.1000 ;
	    RECT 236.6000 165.1000 237.0000 165.2000 ;
	    RECT 239.8000 165.1000 240.2000 165.2000 ;
	    RECT 236.6000 164.8000 240.2000 165.1000 ;
	    RECT 179.8000 153.1000 180.2000 153.2000 ;
	    RECT 254.2000 153.1000 254.6000 153.2000 ;
	    RECT 179.8000 152.8000 254.6000 153.1000 ;
	    RECT 189.4000 147.1000 189.8000 147.2000 ;
	    RECT 212.6000 147.1000 213.0000 147.2000 ;
	    RECT 189.4000 146.8000 213.0000 147.1000 ;
	    RECT 126.2000 127.1000 126.6000 127.2000 ;
	    RECT 145.4000 127.1000 145.8000 127.2000 ;
	    RECT 126.2000 126.8000 145.8000 127.1000 ;
	    RECT 231.0000 114.1000 231.4000 114.2000 ;
	    RECT 251.0000 114.1000 251.4000 114.2000 ;
	    RECT 231.0000 113.8000 251.4000 114.1000 ;
	    RECT 190.2000 92.1000 190.6000 92.2000 ;
	    RECT 237.4000 92.1000 237.8000 92.2000 ;
	    RECT 190.2000 91.8000 237.8000 92.1000 ;
	    RECT 187.8000 89.1000 188.2000 89.2000 ;
	    RECT 223.8000 89.1000 224.2000 89.2000 ;
	    RECT 187.8000 88.8000 224.2000 89.1000 ;
	    RECT 207.0000 87.1000 207.4000 87.2000 ;
	    RECT 252.6000 87.1000 253.0000 87.2000 ;
	    RECT 207.0000 86.8000 253.0000 87.1000 ;
	    RECT 223.0000 86.1000 223.4000 86.2000 ;
	    RECT 225.4000 86.1000 225.8000 86.2000 ;
	    RECT 223.0000 85.8000 225.8000 86.1000 ;
	    RECT 8.6000 77.1000 9.0000 77.2000 ;
	    RECT 11.8000 77.1000 12.2000 77.2000 ;
	    RECT 8.6000 76.8000 12.2000 77.1000 ;
	    RECT 5.4000 76.1000 5.8000 76.2000 ;
	    RECT 23.0000 76.1000 23.4000 76.2000 ;
	    RECT 5.4000 75.8000 23.4000 76.1000 ;
	    RECT 24.6000 75.1000 25.0000 75.2000 ;
	    RECT 27.8000 75.1000 28.2000 75.2000 ;
	    RECT 24.6000 74.8000 28.2000 75.1000 ;
	    RECT 71.0000 74.1000 71.4000 74.2000 ;
	    RECT 101.4000 74.1000 101.8000 74.2000 ;
	    RECT 71.0000 73.8000 101.8000 74.1000 ;
	    RECT 207.8000 74.1000 208.2000 74.2000 ;
	    RECT 243.8000 74.1000 244.2000 74.2000 ;
	    RECT 207.8000 73.8000 244.2000 74.1000 ;
	    RECT 205.4000 67.1000 205.8000 67.2000 ;
	    RECT 238.2000 67.1000 238.6000 67.2000 ;
	    RECT 205.4000 66.8000 238.6000 67.1000 ;
	    RECT 37.4000 54.1000 37.8000 54.2000 ;
	    RECT 135.0000 54.1000 135.4000 54.2000 ;
	    RECT 37.4000 53.8000 135.4000 54.1000 ;
	    RECT 111.0000 25.1000 111.4000 25.2000 ;
	    RECT 135.8000 25.1000 136.2000 25.2000 ;
	    RECT 111.0000 24.8000 136.2000 25.1000 ;
	    RECT 67.0000 15.1000 67.4000 15.2000 ;
	    RECT 71.0000 15.1000 71.4000 15.2000 ;
	    RECT 67.0000 14.8000 71.4000 15.1000 ;
	    RECT 92.6000 15.1000 93.0000 15.2000 ;
	    RECT 124.6000 15.1000 125.0000 15.2000 ;
	    RECT 92.6000 14.8000 125.0000 15.1000 ;
	    RECT 88.6000 14.1000 89.0000 14.2000 ;
	    RECT 102.2000 14.1000 102.6000 14.2000 ;
	    RECT 88.6000 13.8000 102.6000 14.1000 ;
	    RECT 113.4000 14.1000 113.8000 14.2000 ;
	    RECT 119.8000 14.1000 120.2000 14.2000 ;
	    RECT 113.4000 13.8000 120.2000 14.1000 ;
	    RECT 101.4000 13.1000 101.8000 13.2000 ;
	    RECT 117.4000 13.1000 117.8000 13.2000 ;
	    RECT 101.4000 12.8000 117.8000 13.1000 ;
	    RECT 95.0000 12.1000 95.4000 12.2000 ;
	    RECT 133.4000 12.1000 133.8000 12.2000 ;
	    RECT 95.0000 11.8000 133.8000 12.1000 ;
	    RECT 104.6000 9.1000 105.0000 9.2000 ;
	    RECT 126.2000 9.1000 126.6000 9.2000 ;
	    RECT 104.6000 8.8000 126.6000 9.1000 ;
	    RECT 123.8000 8.1000 124.2000 8.2000 ;
	    RECT 131.8000 8.1000 132.2000 8.2000 ;
	    RECT 123.8000 7.8000 132.2000 8.1000 ;
	    RECT 81.4000 7.1000 81.8000 7.2000 ;
	    RECT 88.6000 7.1000 89.0000 7.2000 ;
	    RECT 81.4000 6.8000 89.0000 7.1000 ;
	    RECT 99.8000 7.1000 100.2000 7.2000 ;
	    RECT 103.0000 7.1000 103.4000 7.2000 ;
	    RECT 99.8000 6.8000 103.4000 7.1000 ;
   END
END area_sys
