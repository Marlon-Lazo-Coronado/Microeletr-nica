* NGSPICE file created from area_sys.ext - technology: scmos

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 Q CLK D gnd vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

.subckt area_sys vdd gnd clk reset block0[0] block0[1] block0[2] block0[3] block0[4]
+ block0[5] block0[6] block0[7] block1[0] block1[1] block1[2] block1[3] block1[4]
+ block1[5] block1[6] block1[7] block2[0] block2[1] block2[2] block2[3] block2[4]
+ block2[5] block2[6] block2[7] block3[0] block3[1] block3[2] block3[3] block3[4]
+ block3[5] block3[6] block3[7] block4[0] block4[1] block4[2] block4[3] block4[4]
+ block4[5] block4[6] block4[7] block5[0] block5[1] block5[2] block5[3] block5[4]
+ block5[5] block5[6] block5[7] block6[0] block6[1] block6[2] block6[3] block6[4]
+ block6[5] block6[6] block6[7] block7[0] block7[1] block7[2] block7[3] block7[4]
+ block7[5] block7[6] block7[7] block8[0] block8[1] block8[2] block8[3] block8[4]
+ block8[5] block8[6] block8[7] block9[0] block9[1] block9[2] block9[3] block9[4]
+ block9[5] block9[6] block9[7] block10[0] block10[1] block10[2] block10[3] block10[4]
+ block10[5] block10[6] block10[7] block11[0] block11[1] block11[2] block11[3] block11[4]
+ block11[5] block11[6] block11[7] start target[0] target[1] target[2] target[3] target[4]
+ target[5] target[6] target[7] target[8] target[9] target[10] target[11] target[12]
+ target[13] target[14] target[15] nonce0[0] nonce0[1] nonce0[2] nonce0[3] nonce0[4]
+ nonce0[5] nonce0[6] nonce0[7] nonce1[0] nonce1[1] nonce1[2] nonce1[3] nonce1[4]
+ nonce1[5] nonce1[6] nonce1[7] nonce2[0] nonce2[1] nonce2[2] nonce2[3] nonce2[4]
+ nonce2[5] nonce2[6] nonce2[7] nonce3[0] nonce3[1] nonce3[2] nonce3[3] nonce3[4]
+ nonce3[5] nonce3[6] nonce3[7] finish
XNOR2X1_62 gnd OR2X2_6/A gnd NOR2X1_62/Y vdd NOR2X1
XINVX2_11 OR2X2_23/B gnd INVX2_11/Y vdd INVX2
XFILL_12_2_1 gnd vdd FILL
XFILL_14_0_0 gnd vdd FILL
XNOR2X1_26 NOR2X1_26/A NOR2X1_25/Y gnd NOR2X1_26/Y vdd NOR2X1
XOAI21X1_154 INVX4_5/Y INVX1_212/Y INVX4_4/Y gnd INVX1_215/A vdd OAI21X1
XNOR2X1_187 INVX4_3/Y NOR2X1_182/B gnd NOR2X1_187/Y vdd NOR2X1
XOAI21X1_118 INVX1_180/Y OAI21X1_117/Y OAI21X1_116/Y gnd OAI21X1_118/Y vdd OAI21X1
XNOR2X1_151 BUFX4_47/Y NOR2X1_117/B gnd OAI22X1_8/D vdd NOR2X1
XXNOR2X1_25 OR2X2_22/A OR2X2_23/B gnd AOI21X1_82/A vdd XNOR2X1
XNOR2X1_115 BUFX4_18/Y NAND2X1_80/Y gnd NOR2X1_115/Y vdd NOR2X1
XAOI21X1_94 AOI21X1_94/A AOI21X1_94/B INVX8_3/Y gnd AOI21X1_94/Y vdd AOI21X1
XAOI21X1_58 AOI21X1_58/A AOI21X1_58/B AOI21X1_58/C gnd AOI21X1_59/A vdd AOI21X1
XFILL_1_1_0 gnd vdd FILL
XOR2X2_11 OR2X2_11/A XOR2X1_7/B gnd OR2X2_11/Y vdd OR2X2
XFILL_9_1 gnd vdd FILL
XDFFPOSX1_2 INVX1_39/A CLKBUF1_9/Y DFFPOSX1_2/D gnd vdd DFFPOSX1
XNAND2X1_124 INVX2_14/Y INVX2_15/Y gnd NOR2X1_180/A vdd NAND2X1
XAOI21X1_22 INVX1_31/Y AOI22X1_1/B OR2X2_1/A gnd AOI21X1_22/Y vdd AOI21X1
XDFFPOSX1_88 NAND3X1_5/A CLKBUF1_6/Y NOR2X1_72/Y gnd vdd DFFPOSX1
XOAI21X1_70 NAND2X1_56/B INVX1_108/Y NOR2X1_70/Y gnd OAI21X1_70/Y vdd OAI21X1
XNAND2X1_85 NOR2X1_120/Y INVX2_12/Y gnd NOR2X1_155/B vdd NAND2X1
XBUFX2_25 INVX1_16/A gnd nonce2[7] vdd BUFX2
XBUFX2_3 BUFX2_3/A gnd nonce0[1] vdd BUFX2
XDFFPOSX1_118 AND2X2_28/A CLKBUF1_4/Y AND2X2_27/Y gnd vdd DFFPOSX1
XNAND2X1_49 INVX1_86/A INVX1_96/Y gnd AOI21X1_48/B vdd NAND2X1
XFILL_6_3_1 gnd vdd FILL
XDFFPOSX1_52 INVX1_103/A CLKBUF1_5/Y AOI21X1_9/Y gnd vdd DFFPOSX1
XOAI21X1_34 NOR2X1_48/B OAI21X1_33/Y OAI21X1_34/C gnd AOI21X1_40/C vdd OAI21X1
XFILL_8_1_0 gnd vdd FILL
XDFFPOSX1_16 BUFX2_7/A CLKBUF1_11/Y AOI21X1_22/Y gnd vdd DFFPOSX1
XNAND2X1_13 gnd INVX1_47/Y gnd NAND3X1_20/B vdd NAND2X1
XNAND2X1_2 BUFX4_44/Y INVX1_18/A gnd AOI22X1_1/B vdd NAND2X1
XINVX1_192 INVX1_192/A gnd MUX2X1_4/S vdd INVX1
XOAI22X1_1 INVX1_54/Y gnd INVX1_55/Y gnd gnd OAI22X1_1/Y vdd OAI22X1
XNAND3X1_18 INVX1_37/Y OR2X2_2/A INVX1_38/Y gnd NAND3X1_18/Y vdd NAND3X1
XINVX1_74 target[13] gnd INVX1_74/Y vdd INVX1
XAOI21X1_108 INVX1_215/Y AOI21X1_107/Y AOI21X1_106/Y gnd AOI21X1_108/Y vdd AOI21X1
XINVX1_156 INVX1_156/A gnd INVX1_156/Y vdd INVX1
XINVX1_38 INVX1_38/A gnd INVX1_38/Y vdd INVX1
XNOR2X1_99 INVX1_110/A NOR2X1_99/B gnd NOR2X1_99/Y vdd NOR2X1
XINVX1_120 INVX1_120/A gnd INVX1_120/Y vdd INVX1
XAND2X2_24 OR2X2_23/A OR2X2_23/B gnd AND2X2_24/Y vdd AND2X2
XBUFX4_45 reset gnd BUFX4_45/Y vdd BUFX4
XNOR2X1_63 target[13] INVX1_72/Y gnd OR2X2_7/B vdd NOR2X1
XINVX2_12 INVX2_12/A gnd INVX2_12/Y vdd INVX2
XNOR2X1_27 INVX1_34/A NAND2X1_6/Y gnd AND2X2_3/A vdd NOR2X1
XFILL_14_0_1 gnd vdd FILL
XOAI21X1_155 INVX4_5/Y INVX1_215/A AOI21X1_105/Y gnd NOR2X1_203/B vdd OAI21X1
XNOR2X1_188 AND2X2_34/B block9[0] gnd XOR2X1_16/A vdd NOR2X1
XOAI21X1_119 INVX1_181/Y NOR2X1_160/Y NOR2X1_152/Y gnd OAI21X1_119/Y vdd OAI21X1
XNOR2X1_152 BUFX4_48/Y NOR2X1_118/B gnd NOR2X1_152/Y vdd NOR2X1
XXNOR2X1_26 XNOR2X1_26/A INVX4_5/A gnd XNOR2X1_26/Y vdd XNOR2X1
XFILL_13_3_0 gnd vdd FILL
XNOR2X1_116 OR2X2_23/A INVX1_149/Y gnd NOR2X1_116/Y vdd NOR2X1
XFILL_1_1_1 gnd vdd FILL
XAOI21X1_59 AOI21X1_59/A AOI21X1_59/B AOI21X1_59/C gnd AOI21X1_59/Y vdd AOI21X1
XAOI21X1_95 AOI21X1_95/A AOI21X1_95/B INVX8_3/Y gnd AOI21X1_95/Y vdd AOI21X1
XOR2X2_12 BUFX4_9/Y OR2X2_12/B gnd OR2X2_12/Y vdd OR2X2
XFILL_9_2 gnd vdd FILL
XAOI21X1_23 INVX1_32/Y AOI22X1_1/B OR2X2_1/A gnd AOI21X1_23/Y vdd AOI21X1
XNAND2X1_125 XOR2X1_12/A NOR2X1_176/Y gnd AOI21X1_90/B vdd NAND2X1
XDFFPOSX1_3 NAND2X1_1/A CLKBUF1_12/Y NOR2X1_24/Y gnd vdd DFFPOSX1
XOAI21X1_71 INVX1_120/Y INVX1_40/A BUFX2_34/A gnd AOI21X1_56/C vdd OAI21X1
XDFFPOSX1_89 NAND3X1_6/A CLKBUF1_6/Y NOR2X1_73/Y gnd vdd DFFPOSX1
XNAND2X1_86 AND2X2_15/B NAND2X1_83/B gnd OR2X2_19/A vdd NAND2X1
XBUFX2_26 INVX1_1/A gnd nonce3[0] vdd BUFX2
XNAND2X1_50 NOR2X1_68/A OR2X2_17/B gnd NAND2X1_50/Y vdd NAND2X1
XDFFPOSX1_119 AND2X2_29/B CLKBUF1_9/Y NAND2X1_120/Y gnd vdd DFFPOSX1
XDFFPOSX1_53 OAI22X1_6/B CLKBUF1_5/Y AOI21X1_10/Y gnd vdd DFFPOSX1
XFILL_8_1_1 gnd vdd FILL
XOAI21X1_35 AOI21X1_34/Y AOI21X1_40/C AND2X2_4/Y gnd OAI21X1_35/Y vdd OAI21X1
XBUFX2_4 BUFX2_4/A gnd nonce0[2] vdd BUFX2
XDFFPOSX1_17 BUFX2_8/A CLKBUF1_12/Y AOI21X1_23/Y gnd vdd DFFPOSX1
XNAND2X1_14 gnd INVX2_3/Y gnd NAND2X1_14/Y vdd NAND2X1
XINVX1_193 INVX1_86/A gnd INVX1_193/Y vdd INVX1
XINVX1_75 target[12] gnd INVX1_75/Y vdd INVX1
XNAND3X1_19 NAND3X1_19/A NAND3X1_19/B AOI22X1_5/Y gnd NOR2X1_34/A vdd NAND3X1
XNAND2X1_3 start NAND2X1_1/A gnd INVX1_34/A vdd NAND2X1
XOAI22X1_2 INVX1_50/Y gnd INVX1_51/Y gnd gnd OAI22X1_2/Y vdd OAI22X1
XAOI21X1_109 INVX2_18/Y INVX2_21/Y OAI21X1_156/Y gnd AOI21X1_109/Y vdd AOI21X1
XINVX1_157 INVX1_187/A gnd INVX1_157/Y vdd INVX1
XINVX1_39 INVX1_39/A gnd INVX1_39/Y vdd INVX1
XBUFX4_46 reset gnd INVX8_4/A vdd BUFX4
XINVX1_121 INVX1_121/A gnd INVX1_121/Y vdd INVX1
XAND2X2_25 INVX8_2/A OR2X2_22/B gnd AND2X2_25/Y vdd AND2X2
XBUFX4_10 BUFX4_9/A gnd OR2X2_10/A vdd BUFX4
XNOR2X1_64 NOR2X1_64/A NOR2X1_64/B gnd NOR2X1_64/Y vdd NOR2X1
XNOR2X1_28 AND2X2_3/A NOR2X1_28/B gnd NOR2X1_28/Y vdd NOR2X1
XOAI21X1_156 INVX2_18/Y INVX2_21/Y INVX4_5/A gnd OAI21X1_156/Y vdd OAI21X1
XINVX2_13 OR2X2_22/B gnd OR2X2_20/B vdd INVX2
XNOR2X1_189 INVX4_3/Y NOR2X1_189/B gnd NOR2X1_189/Y vdd NOR2X1
XNOR2X1_153 BUFX4_49/Y NOR2X1_153/B gnd AOI21X1_74/A vdd NOR2X1
XOAI21X1_120 OAI21X1_118/Y NOR2X1_152/Y OAI21X1_119/Y gnd OAI22X1_8/C vdd OAI21X1
XNOR2X1_117 BUFX4_19/Y NOR2X1_117/B gnd INVX1_151/A vdd NOR2X1
XFILL_13_3_1 gnd vdd FILL
XFILL_15_1_0 gnd vdd FILL
XXOR2X1_1 gnd target[7] gnd XOR2X1_1/Y vdd XOR2X1
XAOI21X1_96 AOI21X1_96/A AOI21X1_96/B INVX8_3/Y gnd AOI21X1_96/Y vdd AOI21X1
XAOI21X1_60 AOI21X1_60/A XNOR2X1_14/Y NOR2X1_103/Y gnd AOI21X1_60/Y vdd AOI21X1
XNAND2X1_126 XOR2X1_12/A NOR2X1_177/Y gnd AOI21X1_91/B vdd NAND2X1
XOAI21X1_72 NOR2X1_99/Y OAI21X1_72/B OAI21X1_72/C gnd NAND2X1_68/A vdd OAI21X1
XFILL_2_2_0 gnd vdd FILL
XDFFPOSX1_90 NAND3X1_7/A CLKBUF1_1/Y NOR2X1_74/Y gnd vdd DFFPOSX1
XOR2X2_13 BUFX4_9/Y OR2X2_13/B gnd OR2X2_13/Y vdd OR2X2
XNAND2X1_87 block3[0] BUFX4_34/Y gnd INVX1_154/A vdd NAND2X1
XAOI21X1_24 INVX1_33/Y AOI22X1_1/B OR2X2_1/A gnd AOI21X1_24/Y vdd AOI21X1
XBUFX2_27 INVX1_2/A gnd nonce3[1] vdd BUFX2
XDFFPOSX1_4 NOR2X1_1/A CLKBUF1_12/Y NOR2X1_26/Y gnd vdd DFFPOSX1
XDFFPOSX1_120 AND2X2_27/B CLKBUF1_4/Y NAND2X1_119/Y gnd vdd DFFPOSX1
XNAND2X1_51 NAND2X1_50/Y BUFX4_11/Y gnd NOR2X1_70/B vdd NAND2X1
XDFFPOSX1_54 OR2X2_15/B CLKBUF1_1/Y AOI21X1_11/Y gnd vdd DFFPOSX1
XBUFX2_5 BUFX2_5/A gnd nonce0[3] vdd BUFX2
XOAI21X1_36 INVX1_48/Y target[9] OAI22X1_2/Y gnd OAI21X1_36/Y vdd OAI21X1
XDFFPOSX1_18 BUFX2_9/A CLKBUF1_11/Y AOI21X1_24/Y gnd vdd DFFPOSX1
XNAND2X1_15 gnd INVX1_50/Y gnd NAND3X1_22/A vdd NAND2X1
XFILL_9_2_0 gnd vdd FILL
XFILL_13_1 gnd vdd FILL
XINVX1_194 OR2X2_1/B gnd INVX1_194/Y vdd INVX1
XOAI22X1_3 INVX1_82/Y gnd INVX1_83/Y gnd gnd OAI22X1_3/Y vdd OAI22X1
XINVX1_76 gnd gnd INVX1_76/Y vdd INVX1
XNAND3X1_20 NAND3X1_20/A NAND3X1_20/B OR2X2_4/A gnd NOR2X1_34/B vdd NAND3X1
XNAND2X1_4 NAND2X1_4/A INVX1_34/A gnd NAND2X1_4/Y vdd NAND2X1
XINVX1_40 INVX1_40/A gnd INVX1_40/Y vdd INVX1
XINVX1_158 INVX1_158/A gnd INVX1_158/Y vdd INVX1
XAOI21X1_110 AND2X2_34/B AOI21X1_110/B OAI22X1_9/Y gnd AOI21X1_111/B vdd AOI21X1
XINVX1_122 INVX1_122/A gnd INVX1_122/Y vdd INVX1
XBUFX4_47 INVX8_2/Y gnd BUFX4_47/Y vdd BUFX4
XBUFX4_11 BUFX4_9/A gnd BUFX4_11/Y vdd BUFX4
XAND2X2_26 OR2X2_20/A OR2X2_20/B gnd NOR3X1_5/A vdd AND2X2
XNOR2X1_65 NOR2X1_65/A NOR2X1_65/B gnd NOR2X1_65/Y vdd NOR2X1
XINVX2_14 OR2X2_23/B gnd INVX2_14/Y vdd INVX2
XNOR2X1_29 NOR2X1_25/Y OR2X2_2/Y gnd NOR2X1_29/Y vdd NOR2X1
XOAI21X1_157 AOI21X1_109/Y AND2X2_34/Y NOR2X1_197/Y gnd OAI21X1_157/Y vdd OAI21X1
XNOR2X1_190 XOR2X1_11/A block8[0] gnd XOR2X1_17/A vdd NOR2X1
XNOR2X1_154 BUFX4_49/Y NAND2X1_84/Y gnd INVX1_172/A vdd NOR2X1
XOAI21X1_121 AND2X2_19/B BUFX4_31/Y OAI22X1_8/D gnd OAI22X1_8/B vdd OAI21X1
XFILL_15_1_1 gnd vdd FILL
XAOI21X1_97 AOI21X1_97/A AOI21X1_97/B INVX8_3/Y gnd AOI21X1_97/Y vdd AOI21X1
XNOR2X1_118 BUFX4_20/Y NOR2X1_118/B gnd INVX1_152/A vdd NOR2X1
XXOR2X1_2 target[6] gnd gnd XOR2X1_2/Y vdd XOR2X1
XAOI21X1_61 AOI21X1_61/A NAND3X1_33/C NOR2X1_105/Y gnd OAI21X1_77/C vdd AOI21X1
XNAND2X1_127 OR2X2_23/B INVX2_15/Y gnd NOR2X1_192/A vdd NAND2X1
XFILL_2_2_1 gnd vdd FILL
XFILL_4_0_0 gnd vdd FILL
XNAND2X1_88 AND2X2_15/B NAND2X1_93/B gnd NOR2X1_156/B vdd NAND2X1
XOR2X2_14 BUFX4_9/Y OR2X2_14/B gnd OR2X2_14/Y vdd OR2X2
XAOI21X1_25 NAND2X1_8/B OR2X2_2/A AOI21X1_25/C gnd DFFPOSX1_7/D vdd AOI21X1
XBUFX2_28 INVX1_3/A gnd nonce3[2] vdd BUFX2
XDFFPOSX1_5 NAND2X1_6/A CLKBUF1_11/Y NOR2X1_28/Y gnd vdd DFFPOSX1
XINVX2_1 INVX2_1/A gnd INVX2_1/Y vdd INVX2
XOAI21X1_73 INVX1_132/Y INVX1_134/A OAI22X1_5/Y gnd OAI21X1_74/B vdd OAI21X1
XNAND2X1_52 NOR3X1_1/C NOR2X1_70/Y gnd NOR2X1_71/B vdd NAND2X1
XDFFPOSX1_91 NAND3X1_8/A CLKBUF1_1/Y NOR2X1_76/Y gnd vdd DFFPOSX1
XDFFPOSX1_55 INVX1_106/A CLKBUF1_1/Y AOI21X1_12/Y gnd vdd DFFPOSX1
XBUFX2_6 BUFX2_6/A gnd nonce0[4] vdd BUFX2
XOAI21X1_37 NOR2X1_35/B OAI21X1_36/Y AOI21X1_36/Y gnd OAI21X1_37/Y vdd OAI21X1
XDFFPOSX1_121 AOI21X1_66/B CLKBUF1_3/Y AND2X2_30/Y gnd vdd DFFPOSX1
XDFFPOSX1_19 INVX1_17/A CLKBUF1_11/Y AOI22X1_3/Y gnd vdd DFFPOSX1
XNAND2X1_16 gnd INVX1_51/Y gnd NAND3X1_22/B vdd NAND2X1
XFILL_9_2_1 gnd vdd FILL
XFILL_13_2 gnd vdd FILL
XINVX1_77 gnd gnd INVX1_77/Y vdd INVX1
XOAI22X1_4 INVX1_78/Y gnd INVX1_79/Y gnd gnd OAI22X1_4/Y vdd OAI22X1
XNAND2X1_5 NOR2X1_1/A INVX1_34/Y gnd INVX1_35/A vdd NAND2X1
XINVX1_195 INVX1_195/A gnd INVX1_195/Y vdd INVX1
XINVX1_159 block0[0] gnd INVX1_159/Y vdd INVX1
XINVX1_41 gnd gnd INVX1_41/Y vdd INVX1
XNAND3X1_21 OR2X2_3/Y NAND2X1_14/Y XNOR2X1_1/Y gnd NOR2X1_35/B vdd NAND3X1
XAOI21X1_111 OAI21X1_157/Y AOI21X1_111/B INVX2_17/Y gnd AOI21X1_111/Y vdd AOI21X1
XINVX1_123 INVX1_118/A gnd INVX1_123/Y vdd INVX1
XBUFX4_48 INVX8_2/Y gnd BUFX4_48/Y vdd BUFX4
XAND2X2_27 BUFX2_34/A AND2X2_27/B gnd AND2X2_27/Y vdd AND2X2
XBUFX4_12 BUFX4_9/A gnd OR2X2_11/A vdd BUFX4
XNOR2X1_66 NOR2X1_66/A NOR2X1_66/B gnd NOR2X1_66/Y vdd NOR2X1
XINVX2_15 OR2X2_22/A gnd INVX2_15/Y vdd INVX2
XNOR2X1_30 NOR2X1_30/A NOR2X1_30/B gnd NOR2X1_30/Y vdd NOR2X1
XOAI21X1_158 INVX1_211/Y INVX4_5/A OAI21X1_158/C gnd AOI21X1_110/B vdd OAI21X1
XNOR2X1_191 XOR2X1_12/A block7[0] gnd NOR2X1_191/Y vdd NOR2X1
XNOR2X1_155 BUFX4_49/Y NOR2X1_155/B gnd NOR2X1_155/Y vdd NOR2X1
XOAI21X1_122 OAI22X1_8/Y NOR2X1_150/Y AOI21X1_75/Y gnd AOI21X1_77/B vdd OAI21X1
XAOI21X1_98 AOI21X1_98/A AOI21X1_98/B INVX8_3/Y gnd AOI21X1_98/Y vdd AOI21X1
XNOR2X1_119 INVX2_11/Y INVX2_10/Y gnd NAND2X1_83/B vdd NOR2X1
XXOR2X1_3 target[2] gnd gnd XOR2X1_3/Y vdd XOR2X1
XAOI21X1_62 INVX2_8/Y INVX1_121/A NAND3X1_31/B gnd AOI21X1_62/Y vdd AOI21X1
XFILL_16_2_0 gnd vdd FILL
XBUFX2_29 INVX1_4/A gnd nonce3[3] vdd BUFX2
XFILL_4_0_1 gnd vdd FILL
XOR2X2_15 INVX2_9/Y OR2X2_15/B gnd OR2X2_15/Y vdd OR2X2
XAOI21X1_26 NAND2X1_8/B OR2X2_2/A NAND2X1_8/A gnd NOR2X1_30/B vdd AOI21X1
XNAND2X1_128 XOR2X1_13/A NOR2X1_178/Y gnd AOI21X1_92/B vdd NAND2X1
XDFFPOSX1_6 AND2X2_3/B CLKBUF1_9/Y NOR2X1_29/Y gnd vdd DFFPOSX1
XOAI21X1_74 NAND2X1_70/Y OAI21X1_74/B AOI21X1_60/Y gnd OAI21X1_74/Y vdd OAI21X1
XDFFPOSX1_92 NAND3X1_9/A CLKBUF1_1/Y NOR2X1_77/Y gnd vdd DFFPOSX1
XNAND2X1_89 BUFX4_50/Y AND2X2_15/Y gnd INVX1_155/A vdd NAND2X1
XBUFX2_7 BUFX2_7/A gnd nonce0[5] vdd BUFX2
XINVX2_2 target[15] gnd INVX2_2/Y vdd INVX2
XNAND2X1_53 NAND2X1_53/A NOR2X1_70/Y gnd NOR2X1_72/B vdd NAND2X1
XDFFPOSX1_122 INVX1_202/A CLKBUF1_2/Y NOR3X1_6/Y gnd vdd DFFPOSX1
XNAND2X1_17 NOR2X1_36/Y AND2X2_5/Y gnd AOI21X1_34/C vdd NAND2X1
XDFFPOSX1_56 INVX1_107/A CLKBUF1_8/Y AOI21X1_13/Y gnd vdd DFFPOSX1
XOAI21X1_38 INVX2_2/Y gnd BUFX4_44/Y gnd NOR2X1_47/A vdd OAI21X1
XFILL_3_3_0 gnd vdd FILL
XDFFPOSX1_20 BUFX2_11/A CLKBUF1_11/Y NOR2X1_17/Y gnd vdd DFFPOSX1
XOAI22X1_5 INVX1_134/Y OAI22X1_5/B OAI22X1_5/C INVX1_99/A gnd OAI22X1_5/Y vdd OAI22X1
XINVX1_78 target[9] gnd INVX1_78/Y vdd INVX1
XNAND2X1_6 NAND2X1_6/A NOR2X1_1/A gnd NAND2X1_6/Y vdd NAND2X1
XINVX1_160 INVX1_160/A gnd INVX1_160/Y vdd INVX1
XINVX1_196 OR2X2_23/A gnd INVX1_196/Y vdd INVX1
XINVX1_42 gnd gnd INVX1_42/Y vdd INVX1
XNAND3X1_22 NAND3X1_22/A NAND3X1_22/B AOI22X1_7/Y gnd NOR2X1_35/A vdd NAND3X1
XAOI21X1_112 gnd OAI21X1_161/Y AOI21X1_112/C gnd AND2X2_36/A vdd AOI21X1
XBUFX4_49 INVX8_2/Y gnd BUFX4_49/Y vdd BUFX4
XINVX1_124 INVX1_124/A gnd INVX1_124/Y vdd INVX1
XAND2X2_28 AND2X2_28/A AND2X2_28/B gnd AND2X2_28/Y vdd AND2X2
XBUFX4_13 BUFX4_16/A gnd BUFX4_13/Y vdd BUFX4
XNOR2X1_67 gnd INVX1_95/Y gnd NOR2X1_67/Y vdd NOR2X1
XINVX2_16 gnd gnd MUX2X1_7/A vdd INVX2
XNOR2X1_31 NOR2X1_31/A NOR2X1_31/B gnd NOR2X1_31/Y vdd NOR2X1
XOAI21X1_159 AND2X2_35/Y NOR2X1_205/Y gnd gnd OAI21X1_159/Y vdd OAI21X1
XFILL_11_0_0 gnd vdd FILL
XNOR2X1_192 NOR2X1_192/A NAND3X1_41/Y gnd NOR2X1_192/Y vdd NOR2X1
XNOR2X1_156 BUFX4_50/Y NOR2X1_156/B gnd INVX1_177/A vdd NOR2X1
XOAI21X1_123 AND2X2_20/Y NOR2X1_165/Y NOR2X1_162/Y gnd OAI21X1_124/C vdd OAI21X1
XFILL_4_1 gnd vdd FILL
XAOI21X1_99 AOI21X1_99/A AOI21X1_99/B INVX8_3/Y gnd AOI21X1_99/Y vdd AOI21X1
XNOR2X1_120 OR2X2_22/B INVX1_150/Y gnd NOR2X1_120/Y vdd NOR2X1
XAOI21X1_63 AND2X2_11/B OAI21X1_77/Y AOI21X1_63/C gnd OAI21X1_83/C vdd AOI21X1
XXOR2X1_4 gnd target[7] gnd XOR2X1_4/Y vdd XOR2X1
XFILL_16_2_1 gnd vdd FILL
XOR2X2_16 OR2X2_16/A OR2X2_16/B gnd OR2X2_16/Y vdd OR2X2
XAOI21X1_27 INVX1_36/Y OR2X2_2/A NAND2X1_9/A gnd NOR2X1_31/B vdd AOI21X1
XDFFPOSX1_7 NAND2X1_8/B CLKBUF1_9/Y DFFPOSX1_7/D gnd vdd DFFPOSX1
XNAND2X1_129 block11[0] NOR2X1_179/Y gnd AOI21X1_93/B vdd NAND2X1
XBUFX2_30 INVX1_5/A gnd nonce3[4] vdd BUFX2
XOAI21X1_75 AOI21X1_59/Y OAI21X1_74/Y AND2X2_11/Y gnd OAI21X1_75/Y vdd OAI21X1
XNAND2X1_90 block1[0] BUFX4_34/Y gnd INVX1_156/A vdd NAND2X1
XDFFPOSX1_93 NAND3X1_10/A CLKBUF1_5/Y NOR2X1_78/Y gnd vdd DFFPOSX1
XBUFX2_8 BUFX2_8/A gnd nonce0[6] vdd BUFX2
XINVX2_3 target[10] gnd INVX2_3/Y vdd INVX2
XNAND2X1_54 OAI22X1_5/B NOR3X1_1/Y gnd INVX1_100/A vdd NAND2X1
XDFFPOSX1_123 INVX1_201/A CLKBUF1_7/Y AOI21X1_101/Y gnd vdd DFFPOSX1
XDFFPOSX1_57 INVX1_124/A CLKBUF1_5/Y AOI21X1_14/Y gnd vdd DFFPOSX1
XOAI21X1_39 NOR2X1_34/A OR2X2_4/Y NOR2X1_47/Y gnd AOI21X1_38/C vdd OAI21X1
XNOR2X1_1 NOR2X1_1/A NOR2X1_1/B gnd NOR2X1_1/Y vdd NOR2X1
XDFFPOSX1_21 INVX1_20/A CLKBUF1_6/Y NOR2X1_18/Y gnd vdd DFFPOSX1
XNAND2X1_18 target[3] gnd gnd INVX1_65/A vdd NAND2X1
XFILL_3_3_1 gnd vdd FILL
XFILL_5_1_0 gnd vdd FILL
XNAND2X1_7 AND2X2_3/B AND2X2_3/A gnd NAND2X1_7/Y vdd NAND2X1
XINVX1_197 OR2X2_22/B gnd INVX1_197/Y vdd INVX1
XOAI22X1_6 OAI22X1_6/A OAI22X1_6/B INVX1_131/Y INVX1_103/A gnd OAI22X1_6/Y vdd OAI22X1
XINVX1_79 target[8] gnd INVX1_79/Y vdd INVX1
XNAND3X1_23 NAND3X1_23/A NAND3X1_23/B NAND3X1_23/C gnd NOR2X1_51/A vdd NAND3X1
XINVX1_161 INVX1_161/A gnd INVX1_161/Y vdd INVX1
XINVX1_43 target[14] gnd INVX1_43/Y vdd INVX1
XAND2X2_29 BUFX2_34/A AND2X2_29/B gnd AND2X2_29/Y vdd AND2X2
XBUFX4_50 INVX8_2/Y gnd BUFX4_50/Y vdd BUFX4
XINVX1_125 INVX1_107/A gnd INVX1_125/Y vdd INVX1
XNOR2X1_68 NOR2X1_68/A OR2X2_17/B gnd OR2X2_9/A vdd NOR2X1
XBUFX4_14 BUFX4_16/A gnd BUFX4_14/Y vdd BUFX4
XINVX2_17 INVX2_17/A gnd INVX2_17/Y vdd INVX2
XNOR2X1_32 NOR2X1_32/A INVX1_18/Y gnd NOR2X1_33/B vdd NOR2X1
XOAI21X1_160 AOI22X1_23/D gnd OAI21X1_159/Y gnd NAND2X1_149/B vdd OAI21X1
XNOR2X1_193 INVX1_40/A INVX1_205/Y gnd INVX2_17/A vdd NOR2X1
XFILL_11_0_1 gnd vdd FILL
XNOR2X1_157 INVX1_200/A INVX4_1/A gnd NOR2X1_157/Y vdd NOR2X1
XOAI21X1_124 BUFX4_47/Y NAND2X1_78/Y OAI21X1_124/C gnd AOI21X1_77/C vdd OAI21X1
XFILL_10_3_0 gnd vdd FILL
XNOR2X1_121 INVX8_2/A NOR2X1_159/B gnd NOR2X1_121/Y vdd NOR2X1
XAOI21X1_64 AOI21X1_64/A AOI21X1_64/B AOI21X1_64/C gnd OAI21X1_82/B vdd AOI21X1
XFILL_4_2 gnd vdd FILL
XXOR2X1_5 target[6] gnd gnd XOR2X1_5/Y vdd XOR2X1
XOR2X2_17 INVX8_4/A OR2X2_17/B gnd OR2X2_17/Y vdd OR2X2
XAOI21X1_28 OAI21X1_27/Y NAND3X1_18/Y BUFX4_4/Y gnd AOI21X1_28/Y vdd AOI21X1
XDFFPOSX1_8 NAND2X1_8/A CLKBUF1_12/Y NOR2X1_30/Y gnd vdd DFFPOSX1
XNAND2X1_130 XOR2X1_10/Y NOR2X1_180/Y gnd AOI21X1_94/B vdd NAND2X1
XOAI21X1_76 INVX1_128/Y OR2X2_13/B OAI22X1_6/Y gnd OAI21X1_76/Y vdd OAI21X1
XDFFPOSX1_94 NAND3X1_11/A CLKBUF1_5/Y NOR2X1_79/Y gnd vdd DFFPOSX1
XNAND2X1_91 BUFX4_50/Y AND2X2_16/Y gnd INVX1_158/A vdd NAND2X1
XBUFX2_31 INVX1_6/A gnd nonce3[5] vdd BUFX2
XBUFX2_9 BUFX2_9/A gnd nonce0[7] vdd BUFX2
XINVX2_4 target[15] gnd INVX2_4/Y vdd INVX2
XOAI21X1_40 INVX1_56/A INVX1_65/Y XNOR2X1_4/Y gnd NOR2X1_49/B vdd OAI21X1
XNAND2X1_55 OAI22X1_6/B NOR3X1_2/Y gnd INVX1_104/A vdd NAND2X1
XDFFPOSX1_124 INVX1_200/A CLKBUF1_7/Y AOI21X1_100/Y gnd vdd DFFPOSX1
XDFFPOSX1_58 INVX1_122/A CLKBUF1_8/Y AOI21X1_15/Y gnd vdd DFFPOSX1
XFILL_17_3_0 gnd vdd FILL
XNAND2X1_19 target[1] INVX1_57/Y gnd OAI21X1_32/C vdd NAND2X1
XFILL_5_1_1 gnd vdd FILL
XDFFPOSX1_22 INVX1_21/A CLKBUF1_11/Y NOR2X1_19/Y gnd vdd DFFPOSX1
XNOR2X1_2 start BUFX4_1/Y gnd OR2X2_1/A vdd NOR2X1
XINVX1_198 INVX1_198/A gnd INVX1_198/Y vdd INVX1
XINVX1_80 gnd gnd INVX1_80/Y vdd INVX1
XNAND2X1_8 NAND2X1_8/A NAND2X1_8/B gnd INVX1_36/A vdd NAND2X1
XOAI22X1_7 OAI22X1_7/A OAI22X1_7/B OAI22X1_7/C OAI22X1_7/D gnd OAI22X1_7/Y vdd OAI22X1
XNAND3X1_24 NAND3X1_24/A NAND2X1_33/Y OR2X2_7/A gnd NOR2X1_51/B vdd NAND3X1
XINVX1_162 INVX1_162/A gnd INVX1_162/Y vdd INVX1
XINVX1_44 gnd gnd INVX1_44/Y vdd INVX1
XAND2X2_30 INVX1_39/A AND2X2_30/B gnd AND2X2_30/Y vdd AND2X2
XINVX1_126 INVX1_117/A gnd INVX1_126/Y vdd INVX1
XNOR2X1_69 INVX1_120/A INVX1_97/Y gnd BUFX4_9/A vdd NOR2X1
XBUFX4_15 BUFX4_16/A gnd BUFX4_15/Y vdd BUFX4
XNOR2X1_33 NOR2X1_33/A NOR2X1_33/B gnd NOR2X1_33/Y vdd NOR2X1
XINVX2_18 INVX2_18/A gnd INVX2_18/Y vdd INVX2
XOAI21X1_161 INVX4_4/Y XOR2X1_11/A NAND2X1_150/Y gnd OAI21X1_161/Y vdd OAI21X1
XOR2X2_1 OR2X2_1/A OR2X2_1/B gnd OR2X2_1/Y vdd OR2X2
XNOR2X1_194 INVX4_5/A INVX2_17/Y gnd INVX1_206/A vdd NOR2X1
XNOR2X1_158 NOR2X1_158/A INVX4_1/A gnd NOR2X1_158/Y vdd NOR2X1
XOAI21X1_125 AND2X2_21/B BUFX4_30/Y NOR2X1_166/Y gnd NOR2X1_167/B vdd OAI21X1
XNOR2X1_122 NOR3X1_4/A NAND2X1_84/Y gnd AOI21X1_67/A vdd NOR2X1
XXOR2X1_6 target[2] gnd gnd XOR2X1_6/Y vdd XOR2X1
XFILL_10_3_1 gnd vdd FILL
XFILL_12_1_0 gnd vdd FILL
XAOI21X1_65 NOR2X1_109/Y AOI21X1_65/B OAI21X1_74/Y gnd OAI21X1_83/A vdd AOI21X1
XNAND2X1_131 OR2X2_23/A INVX1_197/Y gnd INVX1_198/A vdd NAND2X1
XDFFPOSX1_9 NAND2X1_9/A CLKBUF1_9/Y NOR2X1_31/Y gnd vdd DFFPOSX1
XBUFX2_32 INVX1_7/A gnd nonce3[6] vdd BUFX2
XNAND2X1_92 block0[0] INVX4_1/A gnd NAND3X1_35/A vdd NAND2X1
XOAI21X1_77 NOR2X1_96/B OAI21X1_76/Y OAI21X1_77/C gnd OAI21X1_77/Y vdd OAI21X1
XDFFPOSX1_95 NAND3X1_12/A CLKBUF1_5/Y NOR2X1_81/Y gnd vdd DFFPOSX1
XAOI21X1_29 INVX2_1/Y INVX1_39/Y OAI21X1_29/Y gnd AOI21X1_30/B vdd AOI21X1
XOR2X2_18 BUFX4_32/Y block8[0] gnd OR2X2_18/Y vdd OR2X2
XINVX2_5 target[10] gnd OR2X2_6/A vdd INVX2
XDFFPOSX1_125 INVX1_178/A CLKBUF1_2/Y AOI21X1_99/Y gnd vdd DFFPOSX1
XDFFPOSX1_59 INVX1_121/A CLKBUF1_5/Y AOI21X1_16/Y gnd vdd DFFPOSX1
XNAND2X1_56 NOR2X1_70/Y NAND2X1_56/B gnd NOR2X1_83/B vdd NAND2X1
XOAI21X1_41 NAND2X1_24/Y NAND2X1_27/Y OR2X2_8/A gnd AND2X2_6/A vdd OAI21X1
XFILL_17_3_1 gnd vdd FILL
XDFFPOSX1_23 BUFX2_14/A CLKBUF1_4/Y NOR2X1_20/Y gnd vdd DFFPOSX1
XNAND2X1_20 NAND2X1_20/A AOI21X1_32/Y gnd NAND2X1_20/Y vdd NAND2X1
XNOR2X1_3 INVX1_2/Y NOR2X1_3/B gnd NOR2X1_3/Y vdd NOR2X1
XINVX1_199 INVX1_199/A gnd INVX1_199/Y vdd INVX1
XFILL_6_2_0 gnd vdd FILL
XINVX1_81 gnd gnd INVX1_81/Y vdd INVX1
XNAND2X1_9 NAND2X1_9/A INVX1_36/Y gnd INVX1_38/A vdd NAND2X1
XOAI22X1_8 OAI22X1_8/A OAI22X1_8/B OAI22X1_8/C OAI22X1_8/D gnd OAI22X1_8/Y vdd OAI22X1
XNAND3X1_25 OR2X2_6/Y NAND3X1_25/B XNOR2X1_7/Y gnd NOR2X1_52/B vdd NAND3X1
XOAI22X1_10 INVX1_217/A INVX1_216/Y AND2X2_37/Y NOR2X1_206/Y gnd NOR3X1_7/C vdd OAI22X1
XINVX1_163 block7[0] gnd INVX1_163/Y vdd INVX1
XINVX1_45 gnd gnd INVX1_45/Y vdd INVX1
XINVX1_127 OR2X2_14/B gnd INVX1_127/Y vdd INVX1
XAND2X2_31 AND2X2_31/A INVX1_202/Y gnd NOR3X1_6/C vdd AND2X2
XBUFX4_16 BUFX4_16/A gnd BUFX4_16/Y vdd BUFX4
XNOR2X1_70 OR2X2_9/Y NOR2X1_70/B gnd NOR2X1_70/Y vdd NOR2X1
XINVX2_19 gnd gnd INVX2_19/Y vdd INVX2
XOR2X2_2 OR2X2_2/A OR2X2_2/B gnd OR2X2_2/Y vdd OR2X2
XNOR2X1_34 NOR2X1_34/A NOR2X1_34/B gnd AND2X2_4/B vdd NOR2X1
XNOR2X1_195 gnd INVX4_4/Y gnd INVX1_207/A vdd NOR2X1
XOAI21X1_162 INVX4_5/A XOR2X1_11/A INVX2_17/A gnd AOI21X1_112/C vdd OAI21X1
XNOR2X1_159 BUFX4_49/Y NOR2X1_159/B gnd AOI21X1_74/C vdd NOR2X1
XOAI21X1_126 AOI21X1_77/Y NOR2X1_167/Y INVX1_171/Y gnd AOI21X1_79/B vdd OAI21X1
XXOR2X1_7 XOR2X1_7/A XOR2X1_7/B gnd XOR2X1_7/Y vdd XOR2X1
XNOR2X1_123 BUFX4_18/Y NOR2X1_155/B gnd INVX1_153/A vdd NOR2X1
XFILL_12_1_1 gnd vdd FILL
XAOI21X1_66 AND2X2_27/B AOI21X1_66/B AOI21X1_66/C gnd AOI21X1_66/Y vdd AOI21X1
XNAND2X1_132 XOR2X1_11/Y NOR2X1_181/Y gnd AOI21X1_95/B vdd NAND2X1
XBUFX2_33 INVX1_8/A gnd nonce3[7] vdd BUFX2
XINVX2_6 INVX2_6/A gnd INVX2_6/Y vdd INVX2
XOR2X2_19 OR2X2_19/A BUFX4_50/Y gnd OR2X2_19/Y vdd OR2X2
XAOI21X1_30 BUFX4_13/Y AOI21X1_30/B AOI21X1_30/C gnd DFFPOSX1_2/D vdd AOI21X1
XOAI21X1_78 INVX2_8/Y INVX1_121/A BUFX4_45/Y gnd NOR2X1_108/A vdd OAI21X1
XNAND2X1_93 NOR2X1_120/Y NAND2X1_93/B gnd NOR2X1_153/B vdd NAND2X1
XFILL_1_0_0 gnd vdd FILL
XNAND2X1_57 OR2X2_9/B OR2X2_9/A gnd NAND2X1_57/Y vdd NAND2X1
XOAI21X1_42 NOR2X1_49/B OAI21X1_42/B AOI21X1_33/Y gnd OAI21X1_42/Y vdd OAI21X1
XDFFPOSX1_96 NAND3X1_13/A CLKBUF1_8/Y NOR2X1_82/Y gnd vdd DFFPOSX1
XDFFPOSX1_60 NAND2X1_1/B CLKBUF1_9/Y NOR2X1_33/Y gnd vdd DFFPOSX1
XNAND2X1_21 gnd INVX1_59/Y gnd NAND2X1_21/Y vdd NAND2X1
XDFFPOSX1_126 NOR2X1_158/A CLKBUF1_2/Y AOI21X1_98/Y gnd vdd DFFPOSX1
XFILL_8_1 gnd vdd FILL
XDFFPOSX1_24 INVX1_23/A CLKBUF1_10/Y NOR2X1_21/Y gnd vdd DFFPOSX1
XNOR2X1_4 INVX1_3/Y BUFX4_39/Y gnd NOR2X1_4/Y vdd NOR2X1
XOAI22X1_9 OAI22X1_9/A MUX2X1_5/B INVX1_214/Y OAI22X1_9/D gnd OAI22X1_9/Y vdd OAI22X1
XFILL_6_2_1 gnd vdd FILL
XFILL_8_0_0 gnd vdd FILL
XINVX1_200 INVX1_200/A gnd INVX1_200/Y vdd INVX1
XINVX1_82 target[5] gnd INVX1_82/Y vdd INVX1
XINVX1_164 INVX1_164/A gnd INVX1_164/Y vdd INVX1
XNAND3X1_26 NAND3X1_26/A NAND3X1_26/B NAND3X1_26/C gnd NOR2X1_52/A vdd NAND3X1
XINVX1_46 target[13] gnd INVX1_46/Y vdd INVX1
XOAI22X1_11 INVX1_217/Y INVX1_216/A INVX1_218/Y OR2X2_5/B gnd NOR3X1_7/A vdd OAI22X1
XINVX1_10 BUFX2_19/A gnd INVX1_10/Y vdd INVX1
XINVX1_128 OAI22X1_6/B gnd INVX1_128/Y vdd INVX1
XAND2X2_32 AND2X2_32/A INVX2_17/A gnd AND2X2_32/Y vdd AND2X2
XBUFX4_17 BUFX4_18/A gnd NOR3X1_4/A vdd BUFX4
XNOR2X1_71 NOR2X1_71/A NOR2X1_71/B gnd NOR2X1_71/Y vdd NOR2X1
XINVX2_20 INVX2_20/A gnd MUX2X1_7/B vdd INVX2
XNOR2X1_35 NOR2X1_35/A NOR2X1_35/B gnd AND2X2_4/A vdd NOR2X1
XNOR2X1_196 INVX1_207/Y INVX1_206/Y gnd MUX2X1_5/S vdd NOR2X1
XOAI21X1_163 INVX2_19/Y INVX4_4/Y INVX2_17/A gnd XNOR2X1_26/A vdd OAI21X1
XOR2X2_3 INVX2_3/Y gnd gnd OR2X2_3/Y vdd OR2X2
XNOR2X1_160 NOR2X1_160/A BUFX4_30/Y gnd NOR2X1_160/Y vdd NOR2X1
XOAI21X1_127 AND2X2_22/Y NOR2X1_171/Y AOI21X1_78/C gnd OAI21X1_127/Y vdd OAI21X1
XNOR2X1_124 OR2X2_22/B OR2X2_23/A gnd AND2X2_15/B vdd NOR2X1
XXOR2X1_8 XOR2X1_8/A XOR2X1_8/B gnd XOR2X1_8/Y vdd XOR2X1
XAOI21X1_67 AOI21X1_67/A XNOR2X1_21/Y NOR2X1_133/Y gnd AOI21X1_67/Y vdd AOI21X1
XBUFX2_34 BUFX2_34/A gnd BUFX2_34/Y vdd BUFX2
XAOI21X1_31 INVX1_40/Y BUFX4_27/Y AOI21X1_31/C gnd DFFPOSX1_1/D vdd AOI21X1
XNAND2X1_133 XOR2X1_12/Y NOR2X1_182/Y gnd AOI21X1_96/B vdd NAND2X1
XOR2X2_20 OR2X2_20/A OR2X2_20/B gnd OR2X2_20/Y vdd OR2X2
XFILL_13_2_0 gnd vdd FILL
XFILL_1_0_1 gnd vdd FILL
XINVX2_7 INVX2_7/A gnd INVX2_7/Y vdd INVX2
XDFFPOSX1_97 NAND3X1_14/A CLKBUF1_5/Y AOI21X1_53/Y gnd vdd DFFPOSX1
XOAI21X1_79 NOR2X1_95/A OR2X2_16/Y OAI21X1_79/C gnd AOI21X1_63/C vdd OAI21X1
XNAND2X1_94 block6[0] BUFX4_32/Y gnd INVX1_162/A vdd NAND2X1
XNOR2X1_5 INVX1_4/Y NOR2X1_5/B gnd NOR2X1_5/Y vdd NOR2X1
XNAND2X1_58 INVX2_8/A INVX1_121/Y gnd NAND2X1_58/Y vdd NAND2X1
XNAND2X1_22 XNOR2X1_2/Y XNOR2X1_3/Y gnd NOR2X1_48/B vdd NAND2X1
XDFFPOSX1_127 XNOR2X1_22/B CLKBUF1_7/Y AOI21X1_97/Y gnd vdd DFFPOSX1
XDFFPOSX1_61 INVX1_216/A CLKBUF1_8/Y AOI22X1_10/Y gnd vdd DFFPOSX1
XOAI21X1_43 AOI21X1_40/Y NAND2X1_24/Y OAI21X1_43/C gnd OAI21X1_43/Y vdd OAI21X1
XFILL_0_3_0 gnd vdd FILL
XAOI21X1_1 AOI21X1_1/A OAI21X1_1/Y BUFX4_4/Y gnd AOI21X1_1/Y vdd AOI21X1
XDFFPOSX1_25 INVX1_24/A CLKBUF1_10/Y NOR2X1_22/Y gnd vdd DFFPOSX1
XFILL_8_0_1 gnd vdd FILL
XINVX1_83 target[4] gnd INVX1_83/Y vdd INVX1
XNAND3X1_27 INVX2_6/A INVX1_98/A XOR2X1_9/B gnd NOR3X1_1/C vdd NAND3X1
XINVX1_201 INVX1_201/A gnd INVX1_201/Y vdd INVX1
XINVX1_165 block9[0] gnd INVX1_165/Y vdd INVX1
XINVX1_47 target[12] gnd INVX1_47/Y vdd INVX1
XFILL_7_3_0 gnd vdd FILL
XINVX1_129 INVX1_103/A gnd INVX1_129/Y vdd INVX1
XINVX1_11 INVX1_11/A gnd INVX1_11/Y vdd INVX1
XAND2X2_33 AND2X2_33/A AND2X2_33/B gnd INVX1_214/A vdd AND2X2
XBUFX4_18 BUFX4_18/A gnd BUFX4_18/Y vdd BUFX4
XNOR2X1_72 NOR3X1_1/Y NOR2X1_72/B gnd NOR2X1_72/Y vdd NOR2X1
XINVX2_21 gnd gnd INVX2_21/Y vdd INVX2
XNOR2X1_36 XOR2X1_1/Y XOR2X1_2/Y gnd NOR2X1_36/Y vdd NOR2X1
XNAND3X1_1 NOR2X1_1/Y AND2X2_2/Y AND2X2_1/Y gnd BUFX4_24/A vdd NAND3X1
XNOR2X1_197 gnd INVX2_19/Y gnd NOR2X1_197/Y vdd NOR2X1
XOR2X2_4 OR2X2_4/A OR2X2_4/B gnd OR2X2_4/Y vdd OR2X2
XOAI21X1_164 INVX1_219/Y OR2X2_8/B BUFX4_44/Y gnd NOR3X1_7/B vdd OAI21X1
XOAI21X1_128 BUFX4_48/Y INVX1_184/Y OAI21X1_127/Y gnd AOI21X1_79/C vdd OAI21X1
XNOR2X1_161 BUFX4_47/Y NAND2X1_97/Y gnd AOI21X1_75/C vdd NOR2X1
XNOR2X1_125 BUFX4_19/Y OR2X2_19/A gnd INVX1_160/A vdd NOR2X1
XXOR2X1_9 XOR2X1_9/A XOR2X1_9/B gnd XOR2X1_9/Y vdd XOR2X1
XAOI21X1_68 AOI21X1_68/A OR2X2_18/Y INVX1_152/Y gnd AOI21X1_69/C vdd AOI21X1
XAOI21X1_32 INVX1_56/Y INVX1_65/A XOR2X1_3/Y gnd AOI21X1_32/Y vdd AOI21X1
XOR2X2_21 OR2X2_21/A OR2X2_21/B gnd MUX2X1_4/B vdd OR2X2
XNAND2X1_134 XOR2X1_13/Y NOR2X1_183/Y gnd AOI21X1_97/B vdd NAND2X1
XFILL_13_2_1 gnd vdd FILL
XFILL_15_0_0 gnd vdd FILL
XOAI21X1_80 NOR2X1_98/Y INVX1_145/Y XNOR2X1_16/Y gnd OAI21X1_82/A vdd OAI21X1
XDFFPOSX1_98 NAND3X1_15/A CLKBUF1_5/Y NOR2X1_83/Y gnd vdd DFFPOSX1
XINVX2_8 INVX2_8/A gnd INVX2_8/Y vdd INVX2
XNAND2X1_95 block8[0] BUFX4_32/Y gnd AOI21X1_68/A vdd NAND2X1
XBUFX2_35 gnd gnd BUFX2_35/Y vdd BUFX2
XNOR2X1_6 INVX1_5/Y NOR2X1_6/B gnd NOR2X1_6/Y vdd NOR2X1
XDFFPOSX1_128 XNOR2X1_23/B CLKBUF1_7/Y AOI21X1_96/Y gnd vdd DFFPOSX1
XNAND2X1_59 INVX1_118/A INVX1_122/Y gnd NAND3X1_31/B vdd NAND2X1
XOAI21X1_44 OR2X2_8/A INVX1_66/Y OAI21X1_43/Y gnd OAI21X1_44/Y vdd OAI21X1
XDFFPOSX1_62 OR2X2_5/B CLKBUF1_8/Y AND2X2_6/Y gnd vdd DFFPOSX1
XDFFPOSX1_26 BUFX2_17/A CLKBUF1_2/Y NOR2X1_23/Y gnd vdd DFFPOSX1
XFILL_2_1_0 gnd vdd FILL
XAOI21X1_2 AOI21X1_2/A OAI21X1_2/Y BUFX4_4/Y gnd AOI21X1_2/Y vdd AOI21X1
XNAND2X1_23 INVX1_216/A INVX1_64/Y gnd AOI22X1_10/A vdd NAND2X1
XFILL_0_3_1 gnd vdd FILL
XNAND3X1_28 OAI22X1_5/B XOR2X1_8/B NOR3X1_1/Y gnd NOR3X1_2/C vdd NAND3X1
XINVX1_84 INVX1_84/A gnd INVX1_84/Y vdd INVX1
XINVX1_202 INVX1_202/A gnd INVX1_202/Y vdd INVX1
XFILL_12_1 gnd vdd FILL
XINVX1_166 block11[0] gnd INVX1_166/Y vdd INVX1
XINVX1_12 INVX1_12/A gnd INVX1_12/Y vdd INVX1
XINVX1_48 gnd gnd INVX1_48/Y vdd INVX1
XAND2X2_34 INVX4_5/Y AND2X2_34/B gnd AND2X2_34/Y vdd AND2X2
XINVX1_130 OR2X2_13/B gnd OAI22X1_6/A vdd INVX1
XFILL_7_3_1 gnd vdd FILL
XFILL_9_1_0 gnd vdd FILL
XNOR2X1_73 NOR2X1_73/A NOR2X1_73/B gnd NOR2X1_73/Y vdd NOR2X1
XBUFX4_19 BUFX4_18/A gnd BUFX4_19/Y vdd BUFX4
XNOR2X1_37 target[3] gnd gnd INVX1_56/A vdd NOR2X1
XNAND3X1_2 NAND3X1_2/A BUFX4_27/Y BUFX4_13/Y gnd AOI21X1_2/A vdd NAND3X1
XNOR2X1_198 INVX4_5/A NOR2X1_198/B gnd MUX2X1_7/S vdd NOR2X1
XOR2X2_5 OR2X2_8/A OR2X2_5/B gnd OR2X2_5/Y vdd OR2X2
XOAI21X1_129 INVX1_202/A BUFX4_36/Y AND2X2_16/Y gnd OAI21X1_130/A vdd OAI21X1
XNOR2X1_162 BUFX4_47/Y NAND2X1_80/Y gnd NOR2X1_162/Y vdd NOR2X1
XNOR2X1_126 AND2X2_14/A AND2X2_14/B gnd NOR2X1_126/Y vdd NOR2X1
XAOI21X1_69 INVX1_152/Y AOI21X1_69/B AOI21X1_69/C gnd AOI21X1_70/B vdd AOI21X1
XAOI21X1_33 NAND2X1_21/Y NOR2X1_41/Y NOR2X1_40/Y gnd AOI21X1_33/Y vdd AOI21X1
XNAND2X1_135 INVX4_2/Y NOR2X1_184/Y gnd INVX1_199/A vdd NAND2X1
XOR2X2_22 OR2X2_22/A OR2X2_22/B gnd OR2X2_22/Y vdd OR2X2
XFILL_15_0_1 gnd vdd FILL
XOAI21X1_81 OAI21X1_83/B NAND2X1_75/Y INVX8_4/A gnd AND2X2_13/A vdd OAI21X1
XINVX2_9 INVX2_9/A gnd INVX2_9/Y vdd INVX2
XDFFPOSX1_99 NAND3X1_16/A CLKBUF1_5/Y AOI21X1_55/Y gnd vdd DFFPOSX1
XBUFX2_36 gnd gnd BUFX2_36/Y vdd BUFX2
XNAND2X1_96 NAND2X1_93/B NOR2X1_116/Y gnd NAND2X1_96/Y vdd NAND2X1
XOAI21X1_45 NOR2X1_55/Y NOR2X1_56/Y NAND2X1_39/Y gnd NAND2X1_40/A vdd OAI21X1
XDFFPOSX1_129 OAI21X1_142/C CLKBUF1_7/Y AOI21X1_95/Y gnd vdd DFFPOSX1
XNAND2X1_60 INVX1_124/A INVX1_126/Y gnd NAND3X1_32/A vdd NAND2X1
XDFFPOSX1_63 INVX1_66/A CLKBUF1_8/Y OAI21X1_44/Y gnd vdd DFFPOSX1
XFILL_14_3_0 gnd vdd FILL
XAOI21X1_3 AOI21X1_3/A OAI21X1_3/Y BUFX4_2/Y gnd AOI21X1_3/Y vdd AOI21X1
XNAND2X1_24 AND2X2_4/B AND2X2_4/A gnd NAND2X1_24/Y vdd NAND2X1
XNOR2X1_7 INVX1_6/Y BUFX4_39/Y gnd NOR2X1_7/Y vdd NOR2X1
XDFFPOSX1_27 INVX1_9/A CLKBUF1_12/Y AOI22X1_2/Y gnd vdd DFFPOSX1
XFILL_2_1_1 gnd vdd FILL
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XINVX1_85 gnd gnd INVX1_85/Y vdd INVX1
XINVX1_203 block2[0] gnd INVX1_203/Y vdd INVX1
XNAND3X1_29 OAI22X1_6/B OR2X2_15/B NOR3X1_2/Y gnd NOR3X1_3/C vdd NAND3X1
XFILL_12_2 gnd vdd FILL
XINVX1_49 gnd gnd INVX1_49/Y vdd INVX1
XINVX1_167 INVX1_167/A gnd INVX1_167/Y vdd INVX1
XAND2X2_35 INVX1_204/A gnd gnd AND2X2_35/Y vdd AND2X2
XINVX1_131 OR2X2_12/B gnd INVX1_131/Y vdd INVX1
XFILL_9_1_1 gnd vdd FILL
XINVX1_13 INVX1_13/A gnd INVX1_13/Y vdd INVX1
XNOR2X1_74 INVX1_101/Y NOR2X1_74/B gnd NOR2X1_74/Y vdd NOR2X1
XBUFX4_20 BUFX4_18/A gnd BUFX4_20/Y vdd BUFX4
XNOR2X1_38 target[1] INVX1_57/Y gnd NOR2X1_38/Y vdd NOR2X1
XNAND3X1_3 NAND3X1_3/A BUFX4_28/Y BUFX4_15/Y gnd AOI21X1_3/A vdd NAND3X1
XOR2X2_6 OR2X2_6/A gnd gnd OR2X2_6/Y vdd OR2X2
XNOR2X1_199 gnd INVX4_5/Y gnd INVX1_208/A vdd NOR2X1
XOAI21X1_130 OAI21X1_130/A AND2X2_23/Y BUFX4_20/Y gnd OAI21X1_130/Y vdd OAI21X1
XNOR2X1_163 NOR2X1_163/A BUFX4_31/Y gnd NOR2X1_163/Y vdd NOR2X1
XNOR2X1_127 NOR2X1_126/Y AND2X2_14/Y gnd BUFX4_35/A vdd NOR2X1
XNAND2X1_136 XOR2X1_15/Y NOR2X1_186/Y gnd AOI21X1_99/B vdd NAND2X1
XAOI21X1_70 INVX1_151/Y AOI21X1_70/B OAI21X1_99/Y gnd OAI22X1_7/C vdd AOI21X1
XOAI21X1_82 OAI21X1_82/A OAI21X1_82/B AOI21X1_59/A gnd AOI21X1_65/B vdd OAI21X1
XBUFX2_37 gnd gnd BUFX2_37/Y vdd BUFX2
XAOI21X1_34 AOI21X1_33/Y NAND2X1_20/Y AOI21X1_34/C gnd AOI21X1_34/Y vdd AOI21X1
XOR2X2_23 OR2X2_23/A OR2X2_23/B gnd OR2X2_23/Y vdd OR2X2
XNAND2X1_97 NOR2X1_116/Y NAND2X1_83/B gnd NAND2X1_97/Y vdd NAND2X1
XNAND2X1_100 XOR2X1_12/A BUFX4_33/Y gnd INVX1_168/A vdd NAND2X1
XOAI21X1_46 INVX1_80/Y target[5] OAI22X1_3/Y gnd OAI21X1_46/Y vdd OAI21X1
XNAND2X1_61 INVX1_107/A INVX1_127/Y gnd NAND2X1_61/Y vdd NAND2X1
XDFFPOSX1_130 NOR2X1_160/A CLKBUF1_10/Y AOI21X1_94/Y gnd vdd DFFPOSX1
XFILL_16_1_0 gnd vdd FILL
XDFFPOSX1_64 INVX1_217/A CLKBUF1_8/Y AOI22X1_16/Y gnd vdd DFFPOSX1
XDFFPOSX1_28 BUFX2_19/A CLKBUF1_4/Y NOR2X1_10/Y gnd vdd DFFPOSX1
XNOR2X1_8 INVX1_7/Y NOR2X1_6/B gnd NOR2X1_8/Y vdd NOR2X1
XAOI21X1_4 AOI21X1_4/A AOI21X1_4/B BUFX4_2/Y gnd AOI21X1_4/Y vdd AOI21X1
XOAI21X1_10 BUFX4_23/Y BUFX4_7/Y OAI22X1_6/B gnd AOI21X1_10/B vdd OAI21X1
XNAND2X1_25 AND2X2_5/A AND2X2_5/B gnd NOR2X1_48/A vdd NAND2X1
XFILL_14_3_1 gnd vdd FILL
XINVX1_2 INVX1_2/A gnd INVX1_2/Y vdd INVX1
XINVX1_204 INVX1_204/A gnd MUX2X1_5/B vdd INVX1
XINVX1_86 INVX1_86/A gnd INVX1_86/Y vdd INVX1
XNAND3X1_30 INVX1_124/A INVX1_122/A NOR3X1_3/Y gnd NAND2X1_56/B vdd NAND3X1
XFILL_3_2_0 gnd vdd FILL
XINVX1_168 INVX1_168/A gnd INVX1_168/Y vdd INVX1
XINVX1_50 target[9] gnd INVX1_50/Y vdd INVX1
XINVX1_132 OAI22X1_5/B gnd INVX1_132/Y vdd INVX1
XINVX1_14 BUFX2_23/A gnd INVX1_14/Y vdd INVX1
XAND2X2_36 AND2X2_36/A AND2X2_36/B gnd AND2X2_36/Y vdd AND2X2
XBUFX4_21 BUFX4_18/A gnd INVX8_2/A vdd BUFX4
XNOR2X1_75 NOR3X1_2/A NOR3X1_2/C gnd NOR2X1_75/Y vdd NOR2X1
XNAND3X1_4 NAND3X1_4/A BUFX4_27/Y BUFX4_13/Y gnd AOI21X1_4/A vdd NAND3X1
XNOR2X1_39 target[0] INVX1_58/Y gnd NOR2X1_39/Y vdd NOR2X1
XOR2X2_7 OR2X2_7/A OR2X2_7/B gnd OR2X2_7/Y vdd OR2X2
XNOR2X1_200 gnd INVX1_212/A gnd NOR2X1_201/A vdd NOR2X1
XOAI21X1_131 AOI21X1_79/Y OAI21X1_130/Y INVX8_3/A gnd AOI21X1_80/C vdd OAI21X1
XNOR2X1_164 NOR2X1_163/Y INVX1_182/Y gnd AOI21X1_76/B vdd NOR2X1
XNOR2X1_128 block3[0] BUFX4_34/Y gnd OAI21X1_86/B vdd NOR2X1
XNAND2X1_137 INVX8_3/A NAND2X1_137/B gnd AOI21X1_100/C vdd NAND2X1
XAOI21X1_71 NOR2X1_114/Y AOI21X1_71/B NOR2X1_142/Y gnd AOI21X1_71/Y vdd AOI21X1
XOAI21X1_83 OAI21X1_83/A OAI21X1_83/B OAI21X1_83/C gnd OAI21X1_84/C vdd OAI21X1
XBUFX2_38 gnd gnd BUFX2_38/Y vdd BUFX2
XAOI21X1_35 NOR2X1_43/Y XNOR2X1_2/Y NOR2X1_42/Y gnd OAI21X1_34/C vdd AOI21X1
XNAND2X1_101 NOR2X1_112/Y NAND2X1_83/B gnd NOR2X1_168/B vdd NAND2X1
XNAND2X1_98 XOR2X1_13/A BUFX4_33/Y gnd INVX1_167/A vdd NAND2X1
XFILL_3_1 gnd vdd FILL
XNAND2X1_62 OR2X2_15/B INVX2_9/Y gnd NAND3X1_33/B vdd NAND2X1
XOAI21X1_47 NOR2X1_65/B OAI21X1_46/Y OAI21X1_47/C gnd AOI21X1_49/C vdd OAI21X1
XDFFPOSX1_65 OR2X2_8/B CLKBUF1_8/Y AND2X2_9/Y gnd vdd DFFPOSX1
XNOR2X1_9 INVX1_8/Y NOR2X1_6/B gnd NOR2X1_9/Y vdd NOR2X1
XNAND2X1_26 XNOR2X1_5/Y XNOR2X1_6/Y gnd NOR2X1_49/A vdd NAND2X1
XOAI21X1_11 BUFX4_25/Y BUFX4_8/Y OR2X2_15/B gnd AOI21X1_11/B vdd OAI21X1
XFILL_16_1_1 gnd vdd FILL
XDFFPOSX1_29 INVX1_11/A CLKBUF1_12/Y NOR2X1_11/Y gnd vdd DFFPOSX1
XDFFPOSX1_131 AND2X2_19/B CLKBUF1_10/Y AOI21X1_93/Y gnd vdd DFFPOSX1
XAOI21X1_5 NAND3X1_5/Y AOI21X1_5/B BUFX4_2/Y gnd AOI21X1_5/Y vdd AOI21X1
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XINVX1_205 BUFX2_34/A gnd INVX1_205/Y vdd INVX1
XINVX1_87 target[3] gnd INVX1_87/Y vdd INVX1
XFILL_3_2_1 gnd vdd FILL
XFILL_5_0_0 gnd vdd FILL
XNAND3X1_31 NAND2X1_58/Y NAND3X1_31/B NAND3X1_31/C gnd NOR2X1_95/A vdd NAND3X1
XINVX1_51 target[8] gnd INVX1_51/Y vdd INVX1
XINVX1_169 INVX1_169/A gnd INVX1_169/Y vdd INVX1
XINVX1_133 INVX1_99/A gnd INVX1_133/Y vdd INVX1
XINVX1_15 INVX1_15/A gnd INVX1_15/Y vdd INVX1
XBUFX4_22 BUFX4_24/A gnd BUFX4_22/Y vdd BUFX4
XAND2X2_37 INVX1_94/A INVX1_66/A gnd AND2X2_37/Y vdd AND2X2
XNOR2X1_76 NOR2X1_75/Y NOR2X1_76/B gnd NOR2X1_76/Y vdd NOR2X1
XNOR2X1_40 gnd INVX1_59/Y gnd NOR2X1_40/Y vdd NOR2X1
XNAND3X1_5 NAND3X1_5/A BUFX4_28/Y BUFX4_15/Y gnd NAND3X1_5/Y vdd NAND3X1
XNOR2X1_201 NOR2X1_201/A INVX1_209/Y gnd AOI22X1_23/D vdd NOR2X1
XOR2X2_8 OR2X2_8/A OR2X2_8/B gnd OR2X2_8/Y vdd OR2X2
XFILL_16_1 gnd vdd FILL
XOAI21X1_132 INVX1_190/A AND2X2_30/B INVX8_3/A gnd AOI21X1_85/C vdd OAI21X1
XNOR2X1_165 AND2X2_20/B BUFX4_31/Y gnd NOR2X1_165/Y vdd NOR2X1
XNOR2X1_129 OR2X2_22/A INVX2_11/Y gnd NAND2X1_93/B vdd NOR2X1
XAOI21X1_72 AOI21X1_72/A AOI21X1_72/B BUFX4_18/Y gnd AOI21X1_72/Y vdd AOI21X1
XNAND2X1_138 INVX8_3/A NAND2X1_138/B gnd NAND2X1_138/Y vdd NAND2X1
XAOI21X1_36 NOR2X1_45/Y XNOR2X1_1/Y NOR2X1_44/Y gnd AOI21X1_36/Y vdd AOI21X1
XBUFX2_39 gnd gnd BUFX2_39/Y vdd BUFX2
XOAI21X1_84 INVX8_4/A INVX1_146/Y OAI21X1_84/C gnd OAI21X1_84/Y vdd OAI21X1
XNAND2X1_102 INVX1_200/A BUFX4_36/Y gnd INVX1_174/A vdd NAND2X1
XFILL_10_2_0 gnd vdd FILL
XNAND2X1_99 NAND2X1_93/B NOR2X1_112/Y gnd NOR2X1_149/B vdd NAND2X1
XNAND2X1_63 OAI22X1_6/B OAI22X1_6/A gnd NAND3X1_34/A vdd NAND2X1
XNAND2X1_27 NOR2X1_48/Y NOR2X1_49/Y gnd NAND2X1_27/Y vdd NAND2X1
XOAI21X1_12 BUFX4_25/Y BUFX4_8/Y INVX1_106/A gnd AOI21X1_12/B vdd OAI21X1
XOAI21X1_48 AOI21X1_43/Y AOI21X1_49/C AND2X2_7/Y gnd OAI21X1_48/Y vdd OAI21X1
XDFFPOSX1_132 XNOR2X1_24/B CLKBUF1_10/Y AOI21X1_92/Y gnd vdd DFFPOSX1
XDFFPOSX1_66 INVX1_94/A CLKBUF1_8/Y OAI21X1_57/Y gnd vdd DFFPOSX1
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XAOI21X1_6 NAND3X1_6/Y OAI21X1_6/Y BUFX4_2/Y gnd AOI21X1_6/Y vdd AOI21X1
XDFFPOSX1_30 INVX1_12/A CLKBUF1_12/Y NOR2X1_12/Y gnd vdd DFFPOSX1
XINVX1_88 target[2] gnd INVX1_88/Y vdd INVX1
XFILL_17_2_0 gnd vdd FILL
XINVX1_206 INVX1_206/A gnd INVX1_206/Y vdd INVX1
XFILL_5_0_1 gnd vdd FILL
XINVX1_170 AND2X2_34/B gnd INVX1_170/Y vdd INVX1
XINVX1_52 gnd gnd INVX1_52/Y vdd INVX1
XNAND3X1_32 NAND3X1_32/A NAND2X1_61/Y OR2X2_16/A gnd NOR2X1_95/B vdd NAND3X1
XINVX1_134 INVX1_134/A gnd INVX1_134/Y vdd INVX1
XINVX1_16 INVX1_16/A gnd INVX1_16/Y vdd INVX1
XFILL_4_3_0 gnd vdd FILL
XBUFX4_23 BUFX4_24/A gnd BUFX4_23/Y vdd BUFX4
XNOR2X1_77 NOR3X1_2/Y NOR2X1_77/B gnd NOR2X1_77/Y vdd NOR2X1
XNOR2X1_41 gnd INVX1_60/Y gnd NOR2X1_41/Y vdd NOR2X1
XNAND3X1_6 NAND3X1_6/A BUFX4_28/Y BUFX4_15/Y gnd NAND3X1_6/Y vdd NAND3X1
XOR2X2_9 OR2X2_9/A OR2X2_9/B gnd OR2X2_9/Y vdd OR2X2
XNOR2X1_202 gnd gnd gnd INVX1_211/A vdd NOR2X1
XFILL_16_2 gnd vdd FILL
XOAI21X1_133 OR2X2_22/Y OR2X2_23/Y BUFX4_20/Y gnd AOI21X1_88/B vdd OAI21X1
XNOR2X1_166 BUFX4_48/Y NAND2X1_78/Y gnd NOR2X1_166/Y vdd NOR2X1
XNOR2X1_130 BUFX4_20/Y NOR2X1_156/B gnd INVX1_161/A vdd NOR2X1
XAOI21X1_73 INVX1_175/Y INVX4_1/Y AOI21X1_73/C gnd AOI21X1_73/Y vdd AOI21X1
XNAND2X1_139 INVX1_203/Y NOR2X1_191/Y gnd AOI21X1_102/B vdd NAND2X1
XAOI21X1_37 INVX2_2/Y gnd NAND3X1_19/B gnd NOR2X1_47/B vdd AOI21X1
XOAI21X1_85 AND2X2_27/B AOI21X1_66/B BUFX2_34/A gnd AOI21X1_66/C vdd OAI21X1
XBUFX2_40 gnd gnd BUFX2_40/Y vdd BUFX2
XNAND2X1_103 BUFX4_19/Y AND2X2_15/Y gnd INVX1_176/A vdd NAND2X1
XFILL_10_2_1 gnd vdd FILL
XFILL_12_0_0 gnd vdd FILL
XDFFPOSX1_67 INVX1_40/A CLKBUF1_3/Y AOI21X1_56/Y gnd vdd DFFPOSX1
XNAND2X1_64 INVX1_103/A INVX1_131/Y gnd NAND2X1_64/Y vdd NAND2X1
XOAI21X1_49 INVX1_76/Y target[9] OAI22X1_4/Y gnd OAI21X1_50/B vdd OAI21X1
XDFFPOSX1_133 NOR2X1_163/A CLKBUF1_10/Y AOI21X1_91/Y gnd vdd DFFPOSX1
XNAND2X1_28 gnd INVX1_67/Y gnd AOI21X1_39/A vdd NAND2X1
XAOI21X1_7 AOI21X1_7/A AOI21X1_7/B BUFX4_3/Y gnd AOI21X1_7/Y vdd AOI21X1
XOAI21X1_13 BUFX4_22/Y BUFX4_6/Y INVX1_107/A gnd AOI21X1_13/B vdd OAI21X1
XDFFPOSX1_31 INVX1_13/A CLKBUF1_12/Y NOR2X1_13/Y gnd vdd DFFPOSX1
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
XFILL_17_2_1 gnd vdd FILL
XINVX1_207 INVX1_207/A gnd INVX1_207/Y vdd INVX1
XINVX1_53 gnd gnd INVX1_53/Y vdd INVX1
XNAND3X1_33 OR2X2_15/Y NAND3X1_33/B NAND3X1_33/C gnd NOR2X1_96/B vdd NAND3X1
XINVX1_89 target[7] gnd INVX1_89/Y vdd INVX1
XINVX1_17 INVX1_17/A gnd INVX1_17/Y vdd INVX1
XINVX1_171 INVX1_171/A gnd INVX1_171/Y vdd INVX1
XINVX1_135 INVX1_135/A gnd OAI22X1_5/C vdd INVX1
XNOR3X1_1 INVX2_7/Y NOR3X1_1/B NOR3X1_1/C gnd NOR3X1_1/Y vdd NOR3X1
XFILL_4_3_1 gnd vdd FILL
XFILL_6_1_0 gnd vdd FILL
XBUFX4_24 BUFX4_24/A gnd BUFX4_24/Y vdd BUFX4
XNOR2X1_78 NOR2X1_78/A INVX1_104/Y gnd NOR2X1_78/Y vdd NOR2X1
XNAND3X1_7 NAND3X1_7/A BUFX4_28/Y BUFX4_16/Y gnd AOI21X1_7/A vdd NAND3X1
XNOR2X1_42 gnd INVX1_61/Y gnd NOR2X1_42/Y vdd NOR2X1
XNOR2X1_203 NOR2X1_203/A NOR2X1_203/B gnd NOR2X1_203/Y vdd NOR2X1
XOAI21X1_134 AND2X2_28/A AND2X2_28/B BUFX2_34/A gnd AOI21X1_88/C vdd OAI21X1
XNOR2X1_167 AND2X2_21/Y NOR2X1_167/B gnd NOR2X1_167/Y vdd NOR2X1
XNOR2X1_131 block1[0] BUFX4_34/Y gnd OAI21X1_87/B vdd NOR2X1
XAOI21X1_74 AOI21X1_74/A XNOR2X1_23/Y AOI21X1_74/C gnd AOI21X1_74/Y vdd AOI21X1
XNAND2X1_140 AND2X2_34/B NOR2X1_192/Y gnd AOI21X1_103/B vdd NAND2X1
XAOI21X1_38 AND2X2_4/B OAI21X1_37/Y AOI21X1_38/C gnd OAI21X1_43/C vdd AOI21X1
XNAND2X1_104 INVX1_178/A INVX4_1/A gnd NAND3X1_37/A vdd NAND2X1
XOAI21X1_86 INVX1_154/Y OAI21X1_86/B INVX1_160/A gnd OAI21X1_92/C vdd OAI21X1
XFILL_12_0_1 gnd vdd FILL
XBUFX2_41 gnd gnd BUFX2_41/Y vdd BUFX2
XNAND2X1_65 NOR2X1_97/Y AND2X2_12/Y gnd AOI21X1_59/C vdd NAND2X1
XDFFPOSX1_68 INVX1_148/A CLKBUF1_3/Y NOR2X1_84/Y gnd vdd DFFPOSX1
XDFFPOSX1_134 AND2X2_20/B CLKBUF1_10/Y AOI21X1_90/Y gnd vdd DFFPOSX1
XOAI21X1_50 NOR2X1_52/B OAI21X1_50/B AOI21X1_45/Y gnd AOI21X1_47/B vdd OAI21X1
XDFFPOSX1_32 BUFX2_23/A CLKBUF1_6/Y NOR2X1_14/Y gnd vdd DFFPOSX1
XAOI21X1_8 AOI21X1_8/A AOI21X1_8/B BUFX4_3/Y gnd AOI21X1_8/Y vdd AOI21X1
XNAND2X1_29 OR2X2_1/B INVX1_68/Y gnd NAND2X1_29/Y vdd NAND2X1
XOAI21X1_14 BUFX4_22/Y BUFX4_6/Y INVX1_124/A gnd AOI21X1_14/B vdd OAI21X1
XFILL_11_3_0 gnd vdd FILL
XAND2X2_1 AND2X2_1/A AND2X2_1/B gnd AND2X2_1/Y vdd AND2X2
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XINVX1_208 INVX1_208/A gnd INVX1_208/Y vdd INVX1
XNAND3X1_34 NAND3X1_34/A NAND2X1_64/Y NAND3X1_34/C gnd NOR2X1_96/A vdd NAND3X1
XINVX1_90 target[6] gnd INVX1_90/Y vdd INVX1
XFILL_7_1 gnd vdd FILL
XINVX1_54 target[5] gnd INVX1_54/Y vdd INVX1
XINVX1_172 INVX1_172/A gnd MUX2X1_2/S vdd INVX1
XINVX1_136 NOR2X1_98/Y gnd INVX1_136/Y vdd INVX1
XNOR3X1_2 NOR3X1_2/A NOR3X1_2/B NOR3X1_2/C gnd NOR3X1_2/Y vdd NOR3X1
XINVX1_18 INVX1_18/A gnd INVX1_18/Y vdd INVX1
XINVX1_100 INVX1_100/A gnd NOR2X1_73/A vdd INVX1
XFILL_6_1_1 gnd vdd FILL
XBUFX4_25 BUFX4_24/A gnd BUFX4_25/Y vdd BUFX4
XNOR2X1_79 NOR2X1_79/A NOR2X1_79/B gnd NOR2X1_79/Y vdd NOR2X1
XNAND3X1_8 NAND3X1_8/A BUFX4_26/Y BUFX4_16/Y gnd AOI21X1_8/A vdd NAND3X1
XNOR2X1_43 gnd INVX1_62/Y gnd NOR2X1_43/Y vdd NOR2X1
XNOR2X1_204 gnd INVX4_5/Y gnd NOR2X1_204/Y vdd NOR2X1
XOAI21X1_135 NAND3X1_41/Y NOR2X1_177/A INVX8_3/A gnd NOR2X1_174/B vdd OAI21X1
XNOR2X1_168 BUFX4_48/Y NOR2X1_168/B gnd AOI21X1_78/C vdd NOR2X1
XNOR2X1_132 INVX1_161/A OAI21X1_90/Y gnd NOR2X1_132/Y vdd NOR2X1
XNAND2X1_141 NOR2X1_197/Y INVX1_206/A gnd MUX2X1_6/S vdd NAND2X1
XAOI21X1_75 NOR2X1_150/Y XNOR2X1_24/Y AOI21X1_75/C gnd AOI21X1_75/Y vdd AOI21X1
XAOI21X1_39 AOI21X1_39/A NAND2X1_29/Y NOR2X1_50/Y gnd OAI21X1_42/B vdd AOI21X1
XOAI21X1_87 INVX1_156/Y OAI21X1_87/B INVX1_155/Y gnd OAI21X1_87/Y vdd OAI21X1
XNAND2X1_105 NOR2X1_158/A INVX4_1/A gnd INVX1_179/A vdd NAND2X1
XDFFPOSX1_69 INVX1_110/A CLKBUF1_3/Y NOR2X1_85/Y gnd vdd DFFPOSX1
XNAND2X1_66 OR2X2_10/B INVX2_7/A gnd INVX1_145/A vdd NAND2X1
XOAI21X1_51 INVX2_4/Y gnd BUFX4_44/Y gnd NOR2X1_64/A vdd OAI21X1
XDFFPOSX1_135 AND2X2_21/B CLKBUF1_10/Y AOI21X1_89/Y gnd vdd DFFPOSX1
XAOI21X1_9 AOI21X1_9/A OAI21X1_9/Y BUFX4_3/Y gnd AOI21X1_9/Y vdd AOI21X1
XOAI21X1_15 BUFX4_22/Y BUFX4_6/Y INVX1_122/A gnd AOI21X1_15/B vdd OAI21X1
XFILL_11_3_1 gnd vdd FILL
XDFFPOSX1_33 INVX1_15/A CLKBUF1_11/Y NOR2X1_15/Y gnd vdd DFFPOSX1
XNAND2X1_30 target[15] INVX1_69/Y gnd NAND3X1_23/A vdd NAND2X1
XFILL_13_1_0 gnd vdd FILL
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XAND2X2_2 AND2X2_2/A AND2X2_3/B gnd AND2X2_2/Y vdd AND2X2
XINVX1_209 INVX1_209/A gnd INVX1_209/Y vdd INVX1
XNAND3X1_35 NAND3X1_35/A OAI21X1_88/Y INVX1_158/Y gnd OAI21X1_89/C vdd NAND3X1
XINVX1_91 target[11] gnd INVX1_91/Y vdd INVX1
XFILL_7_2 gnd vdd FILL
XINVX1_55 target[4] gnd INVX1_55/Y vdd INVX1
XINVX1_173 OR2X2_19/Y gnd INVX1_173/Y vdd INVX1
XFILL_0_2_0 gnd vdd FILL
XINVX1_137 INVX1_98/A gnd NOR2X1_99/B vdd INVX1
XNOR3X1_3 NOR3X1_3/A NOR3X1_3/B NOR3X1_3/C gnd NOR3X1_3/Y vdd NOR3X1
XINVX1_19 BUFX2_11/A gnd INVX1_19/Y vdd INVX1
XINVX1_101 NOR3X1_2/C gnd INVX1_101/Y vdd INVX1
XBUFX4_26 BUFX4_28/A gnd BUFX4_26/Y vdd BUFX4
XNAND3X1_9 NAND3X1_9/A BUFX4_26/Y BUFX4_16/Y gnd AOI21X1_9/A vdd NAND3X1
XNOR2X1_80 NOR3X1_3/A NOR3X1_3/C gnd NOR2X1_81/A vdd NOR2X1
XFILL_7_2_0 gnd vdd FILL
XNOR2X1_44 gnd INVX1_63/Y gnd NOR2X1_44/Y vdd NOR2X1
XNOR2X1_205 INVX1_204/A gnd gnd NOR2X1_205/Y vdd NOR2X1
XBUFX4_1 BUFX4_3/A gnd BUFX4_1/Y vdd BUFX4
XOAI21X1_100 AND2X2_17/Y NOR2X1_138/Y INVX1_164/A gnd OAI21X1_101/C vdd OAI21X1
XNOR2X1_169 NOR2X1_169/A BUFX4_30/Y gnd NOR2X1_170/A vdd NOR2X1
XOAI21X1_136 NAND3X1_41/Y NOR2X1_179/A AND2X2_21/B gnd AOI21X1_89/A vdd OAI21X1
XNOR2X1_133 NOR3X1_4/A NOR2X1_153/B gnd NOR2X1_133/Y vdd NOR2X1
XNAND2X1_142 INVX2_19/Y INVX2_17/A gnd NOR2X1_198/B vdd NAND2X1
XAOI21X1_76 AOI21X1_75/C AOI21X1_76/B NOR2X1_162/Y gnd AOI21X1_77/A vdd AOI21X1
XOAI21X1_88 AND2X2_14/Y NOR2X1_126/Y INVX1_159/Y gnd OAI21X1_88/Y vdd OAI21X1
XAOI21X1_40 NOR2X1_48/Y OAI21X1_42/Y AOI21X1_40/C gnd AOI21X1_40/Y vdd AOI21X1
XNAND2X1_106 OAI21X1_142/C BUFX4_36/Y gnd INVX1_180/A vdd NAND2X1
XNAND2X1_67 INVX1_110/A NOR2X1_99/B gnd OAI21X1_72/C vdd NAND2X1
XDFFPOSX1_70 XOR2X1_9/A CLKBUF1_3/Y NOR2X1_86/Y gnd vdd DFFPOSX1
XOAI21X1_52 NOR2X1_51/A OR2X2_7/Y NOR2X1_64/Y gnd AOI21X1_47/C vdd OAI21X1
XDFFPOSX1_100 NOR2X1_68/A CLKBUF1_3/Y AOI22X1_22/Y gnd vdd DFFPOSX1
XOAI21X1_16 BUFX4_22/Y BUFX4_8/Y INVX1_121/A gnd OAI21X1_16/Y vdd OAI21X1
XNAND2X1_31 target[14] INVX1_70/Y gnd NAND3X1_23/B vdd NAND2X1
XDFFPOSX1_34 INVX1_16/A CLKBUF1_12/Y NOR2X1_16/Y gnd vdd DFFPOSX1
XDFFPOSX1_136 NOR2X1_169/A CLKBUF1_10/Y AOI21X1_103/Y gnd vdd DFFPOSX1
XFILL_13_1_1 gnd vdd FILL
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XAND2X2_3 AND2X2_3/A AND2X2_3/B gnd OR2X2_2/A vdd AND2X2
XINVX1_210 INVX1_210/A gnd INVX1_210/Y vdd INVX1
XINVX1_92 OR2X2_8/A gnd INVX1_92/Y vdd INVX1
XINVX1_56 INVX1_56/A gnd INVX1_56/Y vdd INVX1
XINVX1_174 INVX1_174/A gnd INVX1_174/Y vdd INVX1
XNAND3X1_36 INVX1_169/Y NAND3X1_36/B NAND3X1_36/C gnd AOI21X1_80/B vdd NAND3X1
XFILL_0_2_1 gnd vdd FILL
XINVX1_20 INVX1_20/A gnd INVX1_20/Y vdd INVX1
XINVX1_138 INVX2_6/A gnd INVX1_138/Y vdd INVX1
XFILL_2_0_0 gnd vdd FILL
XINVX1_102 XOR2X1_7/A gnd NOR3X1_2/A vdd INVX1
XBUFX4_27 BUFX4_28/A gnd BUFX4_27/Y vdd BUFX4
XNOR3X1_4 NOR3X1_4/A OR2X2_20/B OR2X2_20/A gnd NOR3X1_5/C vdd NOR3X1
XNOR2X1_81 NOR2X1_81/A NOR2X1_81/B gnd NOR2X1_81/Y vdd NOR2X1
XFILL_11_1 gnd vdd FILL
XFILL_7_2_1 gnd vdd FILL
XFILL_9_0_0 gnd vdd FILL
XNOR2X1_45 gnd INVX2_3/Y gnd NOR2X1_45/Y vdd NOR2X1
XNOR2X1_206 INVX1_94/A INVX1_66/A gnd NOR2X1_206/Y vdd NOR2X1
XBUFX4_2 BUFX4_3/A gnd BUFX4_2/Y vdd BUFX4
XOAI21X1_137 NAND3X1_41/Y NOR2X1_180/A AND2X2_20/B gnd AOI21X1_90/A vdd OAI21X1
XNOR2X1_170 NOR2X1_170/A INVX1_183/Y gnd NOR2X1_170/Y vdd NOR2X1
XNOR2X1_134 block7[0] BUFX4_32/Y gnd NOR2X1_134/Y vdd NOR2X1
XOAI21X1_101 BUFX4_19/Y NAND2X1_97/Y OAI21X1_101/C gnd OAI22X1_7/D vdd OAI21X1
XAOI21X1_77 AOI21X1_77/A AOI21X1_77/B AOI21X1_77/C gnd AOI21X1_77/Y vdd AOI21X1
XNAND2X1_143 gnd INVX1_212/A gnd INVX1_209/A vdd NAND2X1
XAOI21X1_41 INVX1_84/Y INVX1_93/A XOR2X1_6/Y gnd AOI21X1_41/Y vdd AOI21X1
XOAI21X1_89 INVX1_157/Y INVX1_158/Y OAI21X1_89/C gnd OAI21X1_89/Y vdd OAI21X1
XNAND2X1_107 NOR2X1_160/A BUFX4_30/Y gnd INVX1_181/A vdd NAND2X1
XDFFPOSX1_71 OR2X2_10/B CLKBUF1_3/Y OR2X2_10/Y gnd vdd DFFPOSX1
XNAND2X1_68 NAND2X1_68/A AOI21X1_57/Y gnd AOI21X1_59/B vdd NAND2X1
XOAI21X1_53 INVX1_84/A INVX1_93/Y XNOR2X1_10/Y gnd NOR2X1_66/B vdd OAI21X1
XNAND2X1_32 gnd INVX1_74/Y gnd NAND3X1_24/A vdd NAND2X1
XOAI21X1_17 BUFX4_1/Y start AOI22X1_1/B gnd BUFX4_38/A vdd OAI21X1
XDFFPOSX1_137 INVX1_195/A CLKBUF1_10/Y NOR2X1_174/Y gnd vdd DFFPOSX1
XDFFPOSX1_101 OR2X2_17/B CLKBUF1_3/Y AND2X2_13/Y gnd vdd DFFPOSX1
XAOI22X1_10 AOI22X1_10/A AND2X2_6/A OAI21X1_35/Y OAI21X1_43/C gnd AOI22X1_10/Y vdd
+ AOI22X1
XDFFPOSX1_35 INVX1_1/A CLKBUF1_12/Y AOI22X1_1/Y gnd vdd DFFPOSX1
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XINVX1_93 INVX1_93/A gnd INVX1_93/Y vdd INVX1
XAND2X2_4 AND2X2_4/A AND2X2_4/B gnd AND2X2_4/Y vdd AND2X2
XINVX1_57 gnd gnd INVX1_57/Y vdd INVX1
XINVX1_211 INVX1_211/A gnd INVX1_211/Y vdd INVX1
XNAND3X1_37 NAND3X1_37/A NAND3X1_37/B INVX1_173/Y gnd NAND3X1_37/Y vdd NAND3X1
XINVX1_175 INVX1_201/A gnd INVX1_175/Y vdd INVX1
XFILL_14_2_0 gnd vdd FILL
XINVX1_139 OR2X2_10/B gnd INVX1_139/Y vdd INVX1
XFILL_2_0_1 gnd vdd FILL
XINVX1_21 INVX1_21/A gnd INVX1_21/Y vdd INVX1
XINVX1_103 INVX1_103/A gnd NOR3X1_2/B vdd INVX1
XBUFX4_28 BUFX4_28/A gnd BUFX4_28/Y vdd BUFX4
XNOR3X1_5 NOR3X1_5/A NOR3X1_5/B NOR3X1_5/C gnd NOR3X1_5/Y vdd NOR3X1
XAOI22X1_1 INVX1_1/Y AOI22X1_1/B BUFX4_39/Y AOI22X1_1/D gnd AOI22X1_1/Y vdd AOI22X1
XFILL_1_3_0 gnd vdd FILL
XFILL_11_2 gnd vdd FILL
XNOR2X1_82 NOR3X1_3/Y NOR2X1_82/B gnd NOR2X1_82/Y vdd NOR2X1
XFILL_9_0_1 gnd vdd FILL
XNOR2X1_46 target[13] INVX1_44/Y gnd OR2X2_4/B vdd NOR2X1
XNOR2X1_10 INVX1_10/Y NOR2X1_5/B gnd NOR2X1_10/Y vdd NOR2X1
XNOR2X1_207 NAND2X1_8/A NAND2X1_8/B gnd AND2X2_1/A vdd NOR2X1
XXNOR2X1_1 gnd target[11] gnd XNOR2X1_1/Y vdd XNOR2X1
XBUFX4_3 BUFX4_3/A gnd BUFX4_3/Y vdd BUFX4
XFILL_8_3_0 gnd vdd FILL
XOAI21X1_138 NOR2X1_179/B NOR2X1_177/A NOR2X1_163/A gnd AOI21X1_91/A vdd OAI21X1
XNOR2X1_171 INVX1_195/A BUFX4_30/Y gnd NOR2X1_171/Y vdd NOR2X1
XNOR2X1_135 INVX1_163/Y INVX4_1/Y gnd NOR2X1_135/Y vdd NOR2X1
XOAI21X1_102 block11[0] BUFX4_32/Y NOR2X1_140/Y gnd OAI22X1_7/B vdd OAI21X1
XAOI21X1_78 INVX1_171/A NOR2X1_170/Y AOI21X1_78/C gnd AOI21X1_78/Y vdd AOI21X1
XNAND2X1_144 INVX4_5/A NOR2X1_197/Y gnd INVX1_210/A vdd NAND2X1
XAOI21X1_42 NAND2X1_41/Y NOR2X1_58/Y NOR2X1_57/Y gnd AOI21X1_42/Y vdd AOI21X1
XOAI21X1_90 OAI21X1_89/Y INVX1_155/Y OAI21X1_87/Y gnd OAI21X1_90/Y vdd OAI21X1
XNAND2X1_108 NOR2X1_163/A BUFX4_31/Y gnd INVX1_182/A vdd NAND2X1
XDFFPOSX1_72 INVX1_135/A CLKBUF1_3/Y NOR2X1_87/Y gnd vdd DFFPOSX1
XNAND2X1_69 INVX2_7/A INVX1_139/Y gnd AOI21X1_58/A vdd NAND2X1
XDFFPOSX1_138 INVX4_5/A CLKBUF1_2/Y XNOR2X1_26/Y gnd vdd DFFPOSX1
XOAI21X1_54 OAI21X1_54/A NAND2X1_47/Y OR2X2_8/A gnd AND2X2_9/A vdd OAI21X1
XDFFPOSX1_102 OR2X2_9/B CLKBUF1_3/Y OAI21X1_84/Y gnd vdd DFFPOSX1
XOAI21X1_18 BUFX4_4/Y start AND2X2_30/B gnd AOI22X1_1/D vdd OAI21X1
XNAND2X1_33 gnd INVX1_75/Y gnd NAND2X1_33/Y vdd NAND2X1
XAOI22X1_11 INVX2_4/Y gnd INVX1_71/Y gnd gnd NAND3X1_23/C vdd AOI22X1
XDFFPOSX1_36 INVX1_2/A CLKBUF1_11/Y NOR2X1_3/Y gnd vdd DFFPOSX1
XAND2X2_5 AND2X2_5/A AND2X2_5/B gnd AND2X2_5/Y vdd AND2X2
XINVX1_212 INVX1_212/A gnd INVX1_212/Y vdd INVX1
XINVX1_58 OR2X2_1/B gnd INVX1_58/Y vdd INVX1
XNAND3X1_38 OR2X2_22/A AND2X2_24/Y AND2X2_25/Y gnd AOI21X1_82/B vdd NAND3X1
XFILL_16_0_0 gnd vdd FILL
XFILL_14_2_1 gnd vdd FILL
XINVX1_94 INVX1_94/A gnd INVX1_94/Y vdd INVX1
XINVX1_22 BUFX2_14/A gnd INVX1_22/Y vdd INVX1
XINVX1_176 INVX1_176/A gnd INVX1_176/Y vdd INVX1
XINVX1_140 XOR2X1_9/A gnd INVX1_140/Y vdd INVX1
XNOR3X1_6 NOR3X1_6/A INVX8_3/Y NOR3X1_6/C gnd NOR3X1_6/Y vdd NOR3X1
XINVX1_104 INVX1_104/A gnd INVX1_104/Y vdd INVX1
XBUFX4_29 BUFX4_28/A gnd INVX8_1/A vdd BUFX4
XFILL_1_3_1 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XNOR2X1_83 NOR2X1_83/A NOR2X1_83/B gnd NOR2X1_83/Y vdd NOR2X1
XAOI22X1_2 INVX1_9/Y AOI22X1_1/B BUFX4_39/Y AOI22X1_2/D gnd AOI22X1_2/Y vdd AOI22X1
XNOR2X1_47 NOR2X1_47/A NOR2X1_47/B gnd NOR2X1_47/Y vdd NOR2X1
XXNOR2X1_2 gnd target[7] gnd XNOR2X1_2/Y vdd XNOR2X1
XNOR2X1_208 INVX1_37/A NAND2X1_9/A gnd AND2X2_1/B vdd NOR2X1
XNOR2X1_11 INVX1_11/Y BUFX4_39/Y gnd NOR2X1_11/Y vdd NOR2X1
XNOR2X1_172 OR2X2_21/B OR2X2_21/A gnd NOR2X1_172/Y vdd NOR2X1
XBUFX4_4 BUFX4_3/A gnd BUFX4_4/Y vdd BUFX4
XFILL_8_3_1 gnd vdd FILL
XOAI21X1_139 NOR2X1_179/B NOR2X1_192/A XNOR2X1_24/B gnd AOI21X1_92/A vdd OAI21X1
XNOR2X1_136 BUFX4_18/Y NAND2X1_96/Y gnd INVX1_164/A vdd NOR2X1
XOAI21X1_103 INVX1_167/Y NOR2X1_141/Y NOR2X1_115/Y gnd OAI21X1_104/C vdd OAI21X1
XNOR2X1_100 INVX1_148/A INVX1_138/Y gnd OAI21X1_72/B vdd NOR2X1
XXNOR2X1_10 target[2] gnd gnd XNOR2X1_10/Y vdd XNOR2X1
XAOI21X1_79 AOI21X1_78/Y AOI21X1_79/B AOI21X1_79/C gnd AOI21X1_79/Y vdd AOI21X1
XNAND2X1_145 INVX4_5/A INVX1_207/A gnd OAI22X1_9/A vdd NAND2X1
XAOI21X1_43 AOI21X1_42/Y NAND2X1_40/Y AOI21X1_43/C gnd AOI21X1_43/Y vdd AOI21X1
XOAI21X1_91 INVX1_161/Y XNOR2X1_19/Y INVX1_160/Y gnd OAI21X1_92/B vdd OAI21X1
XNAND2X1_109 NOR2X1_169/A BUFX4_30/Y gnd INVX1_183/A vdd NAND2X1
XNAND2X1_70 XNOR2X1_14/Y XNOR2X1_15/Y gnd NAND2X1_70/Y vdd NAND2X1
XDFFPOSX1_73 INVX1_134/A CLKBUF1_6/Y NOR2X1_88/Y gnd vdd DFFPOSX1
XDFFPOSX1_139 XOR2X1_11/A CLKBUF1_2/Y AND2X2_36/Y gnd vdd DFFPOSX1
XOAI21X1_55 NOR2X1_66/B OAI21X1_55/B AOI21X1_42/Y gnd OAI21X1_55/Y vdd OAI21X1
XBUFX2_10 INVX1_17/A gnd nonce1[0] vdd BUFX2
XDFFPOSX1_103 INVX1_192/A CLKBUF1_4/Y AOI21X1_66/Y gnd vdd DFFPOSX1
XOAI21X1_19 BUFX4_4/Y start INVX1_86/A gnd AOI22X1_2/D vdd OAI21X1
XDFFPOSX1_37 INVX1_3/A CLKBUF1_10/Y NOR2X1_4/Y gnd vdd DFFPOSX1
XNAND2X1_34 gnd OR2X2_6/A gnd NAND3X1_25/B vdd NAND2X1
XFILL_2_1 gnd vdd FILL
XAND2X2_6 AND2X2_6/A OR2X2_5/Y gnd AND2X2_6/Y vdd AND2X2
XAOI22X1_12 INVX1_72/Y target[13] target[12] INVX1_73/Y gnd OR2X2_7/A vdd AOI22X1
XINVX1_213 OAI22X1_9/A gnd INVX1_213/Y vdd INVX1
XINVX1_95 target[1] gnd INVX1_95/Y vdd INVX1
XNAND3X1_39 OR2X2_22/A OR2X2_23/A OR2X2_23/B gnd OR2X2_20/A vdd NAND3X1
XFILL_16_0_1 gnd vdd FILL
XINVX1_59 target[3] gnd INVX1_59/Y vdd INVX1
XINVX1_177 INVX1_177/A gnd INVX1_177/Y vdd INVX1
XINVX1_141 XOR2X1_7/B gnd INVX1_141/Y vdd INVX1
XINVX1_23 INVX1_23/A gnd INVX1_23/Y vdd INVX1
XFILL_15_3_0 gnd vdd FILL
XNOR3X1_7 NOR3X1_7/A NOR3X1_7/B NOR3X1_7/C gnd NOR3X1_7/Y vdd NOR3X1
XNOR2X1_84 INVX1_109/Y BUFX4_11/Y gnd NOR2X1_84/Y vdd NOR2X1
XFILL_3_1_1 gnd vdd FILL
XINVX1_105 NOR3X1_3/C gnd NOR2X1_79/A vdd INVX1
XAOI22X1_3 INVX1_17/Y AOI22X1_1/B AOI22X1_3/C BUFX4_44/Y gnd AOI22X1_3/Y vdd AOI22X1
XBUFX4_30 BUFX4_35/A gnd BUFX4_30/Y vdd BUFX4
XNOR2X1_48 NOR2X1_48/A NOR2X1_48/B gnd NOR2X1_48/Y vdd NOR2X1
XXNOR2X1_3 target[6] gnd gnd XNOR2X1_3/Y vdd XNOR2X1
XNOR2X1_12 INVX1_12/Y NOR2X1_3/B gnd NOR2X1_12/Y vdd NOR2X1
XBUFX4_5 BUFX4_6/A gnd BUFX4_5/Y vdd BUFX4
XNOR2X1_173 INVX1_188/Y MUX2X1_4/B gnd MUX2X1_4/A vdd NOR2X1
XNOR2X1_209 INVX2_1/A NOR2X1_32/A gnd BUFX4_28/A vdd NOR2X1
XOAI21X1_140 NOR2X1_179/B NOR2X1_179/A AND2X2_19/B gnd AOI21X1_93/A vdd OAI21X1
XNOR2X1_137 block9[0] BUFX4_32/Y gnd NOR2X1_137/Y vdd NOR2X1
XOAI21X1_104 OAI22X1_7/Y NOR2X1_115/Y OAI21X1_104/C gnd OAI21X1_105/A vdd OAI21X1
XNOR2X1_101 INVX2_7/A INVX1_139/Y gnd AOI21X1_58/C vdd NOR2X1
XXNOR2X1_11 target[1] gnd gnd XNOR2X1_11/Y vdd XNOR2X1
XNAND2X1_146 MUX2X1_7/B INVX2_21/Y gnd AND2X2_33/A vdd NAND2X1
XAOI21X1_80 AOI21X1_72/Y AOI21X1_80/B AOI21X1_80/C gnd AOI21X1_80/Y vdd AOI21X1
XOAI21X1_92 NOR2X1_132/Y OAI21X1_92/B OAI21X1_92/C gnd MUX2X1_1/A vdd OAI21X1
XNAND2X1_110 INVX1_39/A INVX8_3/A gnd NOR3X1_5/B vdd NAND2X1
XAOI21X1_44 NOR2X1_60/Y XNOR2X1_8/Y NOR2X1_59/Y gnd OAI21X1_47/C vdd AOI21X1
XNAND2X1_71 NOR2X1_68/A INVX1_144/Y gnd AOI22X1_22/A vdd NAND2X1
XDFFPOSX1_74 XOR2X1_8/A CLKBUF1_6/Y NOR2X1_89/Y gnd vdd DFFPOSX1
XDFFPOSX1_140 AND2X2_34/B CLKBUF1_2/Y AOI21X1_111/Y gnd vdd DFFPOSX1
XBUFX2_11 BUFX2_11/A gnd nonce1[1] vdd BUFX2
XOAI21X1_56 AOI21X1_49/Y OAI21X1_54/A AOI22X1_16/D gnd OAI21X1_56/Y vdd OAI21X1
XDFFPOSX1_38 INVX1_4/A CLKBUF1_4/Y NOR2X1_5/Y gnd vdd DFFPOSX1
XDFFPOSX1_104 INVX1_191/A CLKBUF1_4/Y gnd gnd vdd DFFPOSX1
XNAND2X1_35 gnd INVX1_78/Y gnd NAND3X1_26/A vdd NAND2X1
XOAI21X1_20 INVX1_18/Y OR2X2_1/B start gnd AOI22X1_3/C vdd OAI21X1
XFILL_10_1_0 gnd vdd FILL
XAOI22X1_13 INVX1_76/Y target[9] target[8] INVX1_77/Y gnd NAND3X1_26/C vdd AOI22X1
XAND2X2_7 AND2X2_7/A AND2X2_7/B gnd AND2X2_7/Y vdd AND2X2
XINVX1_214 INVX1_214/A gnd INVX1_214/Y vdd INVX1
XINVX1_96 target[0] gnd INVX1_96/Y vdd INVX1
XNAND3X1_40 OR2X2_23/A OR2X2_23/B OR2X2_22/A gnd OR2X2_21/A vdd NAND3X1
XINVX1_60 target[2] gnd INVX1_60/Y vdd INVX1
XINVX1_178 INVX1_178/A gnd INVX1_178/Y vdd INVX1
XINVX1_142 XOR2X1_8/A gnd INVX1_142/Y vdd INVX1
XINVX1_24 INVX1_24/A gnd INVX1_24/Y vdd INVX1
XFILL_17_1_0 gnd vdd FILL
XFILL_15_3_1 gnd vdd FILL
XNOR3X1_8 NOR3X1_8/A NOR3X1_8/B NOR3X1_8/C gnd BUFX4_16/A vdd NOR3X1
XAND2X2_10 NOR2X1_70/Y INVX2_6/Y gnd AND2X2_10/Y vdd AND2X2
XINVX1_106 INVX1_106/A gnd NOR3X1_3/A vdd INVX1
XBUFX4_31 BUFX4_35/A gnd BUFX4_31/Y vdd BUFX4
XAOI22X1_4 INVX1_26/Y AOI22X1_1/B OR2X2_1/Y BUFX4_39/Y gnd AOI22X1_4/Y vdd AOI22X1
XNOR2X1_85 INVX1_110/Y OR2X2_10/A gnd NOR2X1_85/Y vdd NOR2X1
XNOR2X1_49 NOR2X1_49/A NOR2X1_49/B gnd NOR2X1_49/Y vdd NOR2X1
XXNOR2X1_4 target[2] gnd gnd XNOR2X1_4/Y vdd XNOR2X1
XNOR2X1_13 INVX1_13/Y NOR2X1_3/B gnd NOR2X1_13/Y vdd NOR2X1
XFILL_4_2_0 gnd vdd FILL
XINVX4_1 INVX4_1/A gnd INVX4_1/Y vdd INVX4
XBUFX4_6 BUFX4_6/A gnd BUFX4_6/Y vdd BUFX4
XOAI21X1_141 NOR2X1_179/B NOR2X1_180/A NOR2X1_160/A gnd AOI21X1_94/A vdd OAI21X1
XNOR2X1_174 INVX1_195/Y NOR2X1_174/B gnd NOR2X1_174/Y vdd NOR2X1
XOAI21X1_105 OAI21X1_105/A NOR2X1_114/Y AOI21X1_71/Y gnd NAND3X1_36/C vdd OAI21X1
XNOR2X1_102 XOR2X1_9/B INVX1_140/Y gnd AOI21X1_58/B vdd NOR2X1
XXNOR2X1_12 target[0] INVX1_86/A gnd NAND2X1_46/B vdd XNOR2X1
XNOR2X1_138 block10[0] BUFX4_33/Y gnd NOR2X1_138/Y vdd NOR2X1
XNAND2X1_147 INVX2_20/A gnd gnd AND2X2_33/B vdd NAND2X1
XAOI21X1_81 OR2X2_22/A AOI21X1_82/B NOR3X1_5/B gnd AOI21X1_81/Y vdd AOI21X1
XNAND2X1_111 OR2X2_22/A OR2X2_23/B gnd NAND2X1_112/B vdd NAND2X1
XOAI21X1_93 MUX2X1_1/Y AOI21X1_67/A AOI21X1_67/Y gnd OAI21X1_93/Y vdd OAI21X1
XAOI21X1_45 NOR2X1_62/Y XNOR2X1_7/Y NOR2X1_61/Y gnd AOI21X1_45/Y vdd AOI21X1
XBUFX2_12 INVX1_20/A gnd nonce1[2] vdd BUFX2
XDFFPOSX1_75 XOR2X1_7/B CLKBUF1_6/Y OR2X2_11/Y gnd vdd DFFPOSX1
XDFFPOSX1_141 INVX1_212/A CLKBUF1_2/Y AOI21X1_108/Y gnd vdd DFFPOSX1
XNAND2X1_72 AND2X2_11/B AND2X2_11/A gnd OAI21X1_83/B vdd NAND2X1
XOAI21X1_57 OR2X2_8/A INVX1_94/Y OAI21X1_56/Y gnd OAI21X1_57/Y vdd OAI21X1
XDFFPOSX1_39 INVX1_5/A CLKBUF1_6/Y NOR2X1_6/Y gnd vdd DFFPOSX1
XDFFPOSX1_105 INVX1_187/A CLKBUF1_7/Y AOI21X1_80/Y gnd vdd DFFPOSX1
XNAND2X1_36 gnd INVX1_79/Y gnd NAND3X1_26/B vdd NAND2X1
XOAI21X1_21 start NAND2X1_1/A BUFX4_44/Y gnd NOR2X1_24/A vdd OAI21X1
XAOI22X1_14 INVX1_80/Y target[5] target[4] INVX1_81/Y gnd AND2X2_8/A vdd AOI22X1
XAND2X2_8 AND2X2_8/A AND2X2_8/B gnd AND2X2_8/Y vdd AND2X2
XFILL_10_1_1 gnd vdd FILL
XINVX1_215 INVX1_215/A gnd INVX1_215/Y vdd INVX1
XINVX1_97 INVX8_4/A gnd INVX1_97/Y vdd INVX1
XXOR2X1_10 block10[0] AND2X2_34/B gnd XOR2X1_10/Y vdd XOR2X1
XINVX1_179 INVX1_179/A gnd INVX1_179/Y vdd INVX1
XINVX1_61 target[7] gnd INVX1_61/Y vdd INVX1
XNAND3X1_41 OR2X2_22/B OR2X2_23/A INVX4_2/Y gnd NAND3X1_41/Y vdd NAND3X1
XINVX1_25 BUFX2_17/A gnd INVX1_25/Y vdd INVX1
XINVX1_143 INVX1_143/A gnd INVX1_143/Y vdd INVX1
XFILL_17_1_1 gnd vdd FILL
XINVX1_107 INVX1_107/A gnd NOR3X1_3/B vdd INVX1
XBUFX4_32 BUFX4_35/A gnd BUFX4_32/Y vdd BUFX4
XAOI22X1_5 INVX2_2/Y gnd INVX1_43/Y gnd gnd AOI22X1_5/Y vdd AOI22X1
XNOR2X1_86 INVX1_111/Y OR2X2_10/A gnd NOR2X1_86/Y vdd NOR2X1
XAND2X2_11 AND2X2_11/A AND2X2_11/B gnd AND2X2_11/Y vdd AND2X2
XNOR2X1_50 gnd INVX1_67/Y gnd NOR2X1_50/Y vdd NOR2X1
XNOR2X1_14 INVX1_14/Y NOR2X1_6/B gnd NOR2X1_14/Y vdd NOR2X1
XXNOR2X1_5 target[1] gnd gnd XNOR2X1_5/Y vdd XNOR2X1
XFILL_4_2_1 gnd vdd FILL
XFILL_6_0_0 gnd vdd FILL
XINVX4_2 INVX8_2/A gnd INVX4_2/Y vdd INVX4
XBUFX4_7 BUFX4_6/A gnd BUFX4_7/Y vdd BUFX4
XOAI21X1_142 NAND3X1_43/Y INVX1_198/A OAI21X1_142/C gnd AOI21X1_95/A vdd OAI21X1
XNOR2X1_175 NOR2X1_179/A NAND3X1_41/Y gnd NOR2X1_175/Y vdd NOR2X1
XXNOR2X1_13 INVX1_106/A INVX1_143/A gnd NAND3X1_33/C vdd XNOR2X1
XNOR2X1_139 INVX1_166/Y INVX4_1/Y gnd OAI22X1_7/A vdd NOR2X1
XOAI21X1_106 AND2X2_18/Y NOR2X1_146/Y NOR2X1_142/Y gnd NAND3X1_36/B vdd OAI21X1
XNOR2X1_103 XOR2X1_7/A INVX1_141/Y gnd NOR2X1_103/Y vdd NOR2X1
XAOI21X1_82 AOI21X1_82/A AOI21X1_82/B NOR3X1_5/B gnd AOI21X1_82/Y vdd AOI21X1
XNAND2X1_148 INVX4_4/Y INVX1_208/A gnd OAI22X1_9/D vdd NAND2X1
XAOI21X1_46 INVX2_4/Y gnd NAND3X1_23/B gnd NOR2X1_64/B vdd AOI21X1
XNAND2X1_73 AND2X2_12/A AND2X2_12/B gnd NOR2X1_109/A vdd NAND2X1
XAOI21X1_10 NAND3X1_10/Y AOI21X1_10/B BUFX4_2/Y gnd AOI21X1_10/Y vdd AOI21X1
XNAND2X1_112 INVX1_185/Y NAND2X1_112/B gnd NAND2X1_113/B vdd NAND2X1
XOAI21X1_94 block6[0] BUFX4_34/Y NOR2X1_133/Y gnd OAI21X1_94/Y vdd OAI21X1
XBUFX2_13 INVX1_21/A gnd nonce1[3] vdd BUFX2
XDFFPOSX1_142 XOR2X1_13/A CLKBUF1_2/Y NOR2X1_203/Y gnd vdd DFFPOSX1
XOAI21X1_58 INVX2_6/Y INVX1_98/Y NOR2X1_70/Y gnd OAI21X1_58/Y vdd OAI21X1
XDFFPOSX1_76 OR2X2_12/B CLKBUF1_1/Y OR2X2_12/Y gnd vdd DFFPOSX1
XNAND2X1_37 NOR2X1_53/Y AND2X2_8/Y gnd AOI21X1_43/C vdd NAND2X1
XOAI21X1_22 INVX1_35/Y NAND2X1_6/A BUFX4_44/Y gnd NOR2X1_28/B vdd OAI21X1
XDFFPOSX1_106 OR2X2_22/A CLKBUF1_7/Y AOI21X1_81/Y gnd vdd DFFPOSX1
XAOI22X1_15 INVX1_82/Y gnd INVX1_83/Y gnd gnd AND2X2_8/B vdd AOI22X1
XDFFPOSX1_40 INVX1_6/A CLKBUF1_10/Y NOR2X1_7/Y gnd vdd DFFPOSX1
XINVX1_98 INVX1_98/A gnd INVX1_98/Y vdd INVX1
XAND2X2_9 AND2X2_9/A OR2X2_8/Y gnd AND2X2_9/Y vdd AND2X2
XCLKBUF1_1 clk gnd CLKBUF1_1/Y vdd CLKBUF1
XXOR2X1_11 XOR2X1_11/A block9[0] gnd XOR2X1_11/Y vdd XOR2X1
XINVX1_62 target[6] gnd INVX1_62/Y vdd INVX1
XINVX1_180 INVX1_180/A gnd INVX1_180/Y vdd INVX1
XNAND3X1_42 OR2X2_22/B INVX4_2/Y INVX1_196/Y gnd NOR2X1_179/B vdd NAND3X1
XINVX1_216 INVX1_216/A gnd INVX1_216/Y vdd INVX1
XINVX1_144 INVX8_4/A gnd INVX1_144/Y vdd INVX1
XFILL_11_2_0 gnd vdd FILL
XINVX1_26 BUFX2_2/A gnd INVX1_26/Y vdd INVX1
XINVX1_108 INVX1_121/A gnd INVX1_108/Y vdd INVX1
XAOI22X1_6 INVX1_44/Y target[13] target[12] INVX1_45/Y gnd OR2X2_4/A vdd AOI22X1
XBUFX4_33 BUFX4_35/A gnd BUFX4_33/Y vdd BUFX4
XAND2X2_12 AND2X2_12/A AND2X2_12/B gnd AND2X2_12/Y vdd AND2X2
XNOR2X1_87 INVX1_112/Y OR2X2_10/A gnd NOR2X1_87/Y vdd NOR2X1
XFILL_6_1 gnd vdd FILL
XNOR2X1_51 NOR2X1_51/A NOR2X1_51/B gnd AND2X2_7/B vdd NOR2X1
XXNOR2X1_6 target[0] OR2X2_1/B gnd XNOR2X1_6/Y vdd XNOR2X1
XINVX4_3 INVX4_3/A gnd INVX4_3/Y vdd INVX4
XFILL_6_0_1 gnd vdd FILL
XNOR2X1_15 INVX1_15/Y NOR2X1_3/B gnd NOR2X1_15/Y vdd NOR2X1
XBUFX4_8 BUFX4_6/A gnd BUFX4_8/Y vdd BUFX4
XOAI21X1_143 NOR2X1_182/B INVX1_198/A XNOR2X1_23/B gnd AOI21X1_96/A vdd OAI21X1
XNOR2X1_176 NOR2X1_180/A NAND3X1_41/Y gnd NOR2X1_176/Y vdd NOR2X1
XFILL_5_3_0 gnd vdd FILL
XOAI21X1_107 AND2X2_14/Y NOR2X1_126/Y INVX1_170/Y gnd AOI21X1_72/A vdd OAI21X1
XNOR2X1_140 BUFX4_20/Y NAND2X1_97/Y gnd NOR2X1_140/Y vdd NOR2X1
XNOR2X1_104 XOR2X1_8/B INVX1_142/Y gnd AOI21X1_60/A vdd NOR2X1
XXNOR2X1_14 XOR2X1_7/A XOR2X1_7/B gnd XNOR2X1_14/Y vdd XNOR2X1
XAOI21X1_83 AOI21X1_82/B AOI21X1_83/B NOR3X1_5/B gnd AOI21X1_83/Y vdd AOI21X1
XNAND2X1_149 INVX1_208/A NAND2X1_149/B gnd AND2X2_36/B vdd NAND2X1
XAOI21X1_47 AND2X2_7/B AOI21X1_47/B AOI21X1_47/C gnd AOI22X1_16/D vdd AOI21X1
XBUFX2_14 BUFX2_14/A gnd nonce1[4] vdd BUFX2
XAOI21X1_11 AOI21X1_11/A AOI21X1_11/B BUFX4_3/Y gnd AOI21X1_11/Y vdd AOI21X1
XNAND2X1_113 OR2X2_20/A NAND2X1_113/B gnd AOI21X1_83/B vdd NAND2X1
XOAI21X1_95 INVX1_162/Y OAI21X1_94/Y OAI21X1_93/Y gnd OAI21X1_97/A vdd OAI21X1
XNAND2X1_74 NAND2X1_74/A NAND2X1_74/B gnd NOR2X1_110/A vdd NAND2X1
XOAI21X1_59 INVX2_7/Y NOR3X1_1/C NOR2X1_70/Y gnd OAI21X1_59/Y vdd OAI21X1
XDFFPOSX1_143 XOR2X1_12/A CLKBUF1_2/Y AND2X2_32/Y gnd vdd DFFPOSX1
XDFFPOSX1_77 OR2X2_13/B CLKBUF1_1/Y OR2X2_13/Y gnd vdd DFFPOSX1
XDFFPOSX1_41 INVX1_7/A CLKBUF1_6/Y NOR2X1_8/Y gnd vdd DFFPOSX1
XNAND2X1_38 target[3] gnd gnd INVX1_93/A vdd NAND2X1
XDFFPOSX1_107 OR2X2_23/B CLKBUF1_4/Y AOI21X1_82/Y gnd vdd DFFPOSX1
XOAI21X1_23 AND2X2_3/A AND2X2_3/B BUFX4_45/Y gnd OR2X2_2/B vdd OAI21X1
XAOI22X1_16 AOI22X1_16/A AND2X2_9/A OAI21X1_48/Y AOI22X1_16/D gnd AOI22X1_16/Y vdd
+ AOI22X1
XINVX1_99 INVX1_99/A gnd NOR3X1_1/B vdd INVX1
XXOR2X1_12 XOR2X1_12/A block8[0] gnd XOR2X1_12/Y vdd XOR2X1
XNAND3X1_43 OR2X2_23/B OR2X2_22/A INVX4_2/Y gnd NAND3X1_43/Y vdd NAND3X1
XMUX2X1_1 MUX2X1_1/A MUX2X1_1/B MUX2X1_1/S gnd MUX2X1_1/Y vdd MUX2X1
XINVX1_63 target[11] gnd INVX1_63/Y vdd INVX1
XINVX1_217 INVX1_217/A gnd INVX1_217/Y vdd INVX1
XCLKBUF1_2 clk gnd CLKBUF1_2/Y vdd CLKBUF1
XFILL_11_2_1 gnd vdd FILL
XINVX1_181 INVX1_181/A gnd INVX1_181/Y vdd INVX1
XINVX1_27 BUFX2_3/A gnd INVX1_27/Y vdd INVX1
XFILL_13_0_0 gnd vdd FILL
XINVX1_145 INVX1_145/A gnd INVX1_145/Y vdd INVX1
XINVX1_109 INVX1_148/A gnd INVX1_109/Y vdd INVX1
XBUFX4_34 BUFX4_35/A gnd BUFX4_34/Y vdd BUFX4
XNOR2X1_88 NOR2X1_88/A OR2X2_11/A gnd NOR2X1_88/Y vdd NOR2X1
XAND2X2_13 AND2X2_13/A OR2X2_17/Y gnd AND2X2_13/Y vdd AND2X2
XAOI22X1_7 INVX1_48/Y target[9] target[8] INVX1_49/Y gnd AOI22X1_7/Y vdd AOI22X1
XFILL_0_1_0 gnd vdd FILL
XNOR2X1_52 NOR2X1_52/A NOR2X1_52/B gnd AND2X2_7/A vdd NOR2X1
XINVX4_4 gnd gnd INVX4_4/Y vdd INVX4
XXNOR2X1_7 gnd target[11] gnd XNOR2X1_7/Y vdd XNOR2X1
XNOR2X1_16 INVX1_16/Y NOR2X1_3/B gnd NOR2X1_16/Y vdd NOR2X1
XBUFX4_9 BUFX4_9/A gnd BUFX4_9/Y vdd BUFX4
XOAI21X1_144 NOR2X1_189/B INVX1_198/A XNOR2X1_22/B gnd AOI21X1_97/A vdd OAI21X1
XNOR2X1_177 NOR2X1_177/A NOR2X1_179/B gnd NOR2X1_177/Y vdd NOR2X1
XFILL_5_3_1 gnd vdd FILL
XFILL_7_1_0 gnd vdd FILL
XOAI21X1_108 INVX1_174/Y NOR2X1_157/Y INVX1_177/A gnd OAI21X1_108/Y vdd OAI21X1
XNOR2X1_141 XOR2X1_13/A BUFX4_33/Y gnd NOR2X1_141/Y vdd NOR2X1
XXNOR2X1_15 XOR2X1_8/A XOR2X1_8/B gnd XNOR2X1_15/Y vdd XNOR2X1
XNOR2X1_105 INVX1_106/A INVX1_143/Y gnd NOR2X1_105/Y vdd NOR2X1
XAOI21X1_84 INVX1_186/Y OR2X2_20/Y NOR3X1_5/B gnd AOI21X1_84/Y vdd AOI21X1
XNAND2X1_150 INVX2_18/Y NOR2X1_204/Y gnd NAND2X1_150/Y vdd NAND2X1
XAOI21X1_48 AOI21X1_48/A AOI21X1_48/B NOR2X1_67/Y gnd OAI21X1_55/B vdd AOI21X1
XOAI21X1_1 BUFX4_23/Y BUFX4_7/Y INVX2_6/A gnd OAI21X1_1/Y vdd OAI21X1
XNAND2X1_114 BUFX4_19/Y OR2X2_22/B gnd OR2X2_21/B vdd NAND2X1
XINVX8_1 INVX8_1/A gnd BUFX4_6/A vdd INVX8
XAOI21X1_12 AOI21X1_12/A AOI21X1_12/B BUFX4_3/Y gnd AOI21X1_12/Y vdd AOI21X1
XOAI21X1_96 NOR2X1_135/Y NOR2X1_134/Y NOR2X1_121/Y gnd OAI21X1_96/Y vdd OAI21X1
XDFFPOSX1_144 INVX2_20/A CLKBUF1_2/Y MUX2X1_7/Y gnd vdd DFFPOSX1
XNAND2X1_75 NOR2X1_109/Y NOR2X1_110/Y gnd NAND2X1_75/Y vdd NAND2X1
XDFFPOSX1_78 INVX2_9/A CLKBUF1_6/Y NOR2X1_90/Y gnd vdd DFFPOSX1
XOAI21X1_60 NOR3X1_1/C INVX2_7/Y NOR3X1_1/B gnd NAND2X1_53/A vdd OAI21X1
XBUFX2_15 INVX1_23/A gnd nonce1[5] vdd BUFX2
XDFFPOSX1_42 INVX1_8/A CLKBUF1_6/Y NOR2X1_9/Y gnd vdd DFFPOSX1
XNAND2X1_39 target[1] INVX1_85/Y gnd NAND2X1_39/Y vdd NAND2X1
XDFFPOSX1_108 OR2X2_23/A CLKBUF1_7/Y AOI21X1_83/Y gnd vdd DFFPOSX1
XOAI21X1_24 OR2X2_2/A NAND2X1_8/B BUFX4_45/Y gnd AOI21X1_25/C vdd OAI21X1
XAOI22X1_17 INVX2_8/Y INVX1_121/A INVX1_123/Y INVX1_122/A gnd NAND3X1_31/C vdd AOI22X1
XXOR2X1_13 XOR2X1_13/A block7[0] gnd XOR2X1_13/Y vdd XOR2X1
XMUX2X1_2 MUX2X1_2/A MUX2X1_2/B MUX2X1_2/S gnd MUX2X1_2/Y vdd MUX2X1
XNAND3X1_44 OR2X2_23/B INVX4_2/Y INVX2_15/Y gnd NOR2X1_182/B vdd NAND3X1
XINVX1_218 OR2X2_8/B gnd INVX1_218/Y vdd INVX1
XCLKBUF1_3 clk gnd CLKBUF1_3/Y vdd CLKBUF1
XINVX1_64 OR2X2_8/A gnd INVX1_64/Y vdd INVX1
XINVX1_182 INVX1_182/A gnd INVX1_182/Y vdd INVX1
XFILL_13_0_1 gnd vdd FILL
XINVX1_146 OR2X2_9/B gnd INVX1_146/Y vdd INVX1
XINVX1_28 BUFX2_4/A gnd INVX1_28/Y vdd INVX1
XINVX1_110 INVX1_110/A gnd INVX1_110/Y vdd INVX1
XNOR2X1_89 NOR2X1_89/A OR2X2_11/A gnd NOR2X1_89/Y vdd NOR2X1
XAND2X2_14 AND2X2_14/A AND2X2_14/B gnd AND2X2_14/Y vdd AND2X2
XBUFX4_35 BUFX4_35/A gnd INVX4_1/A vdd BUFX4
XAOI22X1_8 INVX1_52/Y target[5] target[4] INVX1_53/Y gnd AND2X2_5/A vdd AOI22X1
XFILL_12_3_0 gnd vdd FILL
XFILL_0_1_1 gnd vdd FILL
XNOR2X1_53 XOR2X1_4/Y XOR2X1_5/Y gnd NOR2X1_53/Y vdd NOR2X1
XXNOR2X1_8 gnd target[7] gnd XNOR2X1_8/Y vdd XNOR2X1
XNOR2X1_17 INVX1_19/Y NOR2X1_6/B gnd NOR2X1_17/Y vdd NOR2X1
XINVX4_5 INVX4_5/A gnd INVX4_5/Y vdd INVX4
XOAI21X1_145 INVX1_199/A INVX1_198/A NOR2X1_158/A gnd AOI21X1_98/A vdd OAI21X1
XNOR2X1_178 NOR2X1_192/A NOR2X1_179/B gnd NOR2X1_178/Y vdd NOR2X1
XFILL_7_1_1 gnd vdd FILL
XOAI21X1_109 INVX1_175/Y INVX4_1/Y INVX1_176/Y gnd AOI21X1_73/C vdd OAI21X1
XFILL_10_1 gnd vdd FILL
XNOR2X1_142 INVX8_2/A NOR2X1_149/B gnd NOR2X1_142/Y vdd NOR2X1
XXNOR2X1_16 XOR2X1_9/A XOR2X1_9/B gnd XNOR2X1_16/Y vdd XNOR2X1
XNOR2X1_106 OR2X2_15/B INVX2_9/Y gnd AOI21X1_61/A vdd NOR2X1
XAOI21X1_85 INVX1_187/Y INVX1_190/A AOI21X1_85/C gnd AOI21X1_85/Y vdd AOI21X1
XNAND2X1_151 AND2X2_1/A AND2X2_1/B gnd NOR3X1_8/C vdd NAND2X1
XOAI21X1_2 BUFX4_23/Y BUFX4_7/Y INVX1_98/A gnd OAI21X1_2/Y vdd OAI21X1
XNAND2X1_115 INVX8_3/A NOR2X1_172/Y gnd NAND2X1_115/Y vdd NAND2X1
XAOI21X1_49 NOR2X1_65/Y OAI21X1_55/Y AOI21X1_49/C gnd AOI21X1_49/Y vdd AOI21X1
XOAI21X1_97 OAI21X1_97/A NOR2X1_121/Y OAI21X1_96/Y gnd AOI21X1_69/B vdd OAI21X1
XINVX8_2 INVX8_2/A gnd INVX8_2/Y vdd INVX8
XAOI21X1_13 NAND3X1_13/Y AOI21X1_13/B BUFX4_1/Y gnd AOI21X1_13/Y vdd AOI21X1
XNAND2X1_76 INVX1_98/A INVX1_147/Y gnd AOI21X1_64/A vdd NAND2X1
XDFFPOSX1_145 INVX2_18/A CLKBUF1_4/Y MUX2X1_6/Y gnd vdd DFFPOSX1
XOAI21X1_61 OAI22X1_5/B NOR3X1_1/Y NOR2X1_70/Y gnd NOR2X1_73/B vdd OAI21X1
XDFFPOSX1_79 INVX1_143/A CLKBUF1_8/Y NOR2X1_91/Y gnd vdd DFFPOSX1
XBUFX2_16 INVX1_24/A gnd nonce1[6] vdd BUFX2
XNAND2X1_40 NAND2X1_40/A AOI21X1_41/Y gnd NAND2X1_40/Y vdd NAND2X1
XDFFPOSX1_109 OR2X2_22/B CLKBUF1_7/Y NOR3X1_5/Y gnd vdd DFFPOSX1
XOAI21X1_25 NAND2X1_7/Y INVX1_36/A BUFX4_45/Y gnd NOR2X1_30/A vdd OAI21X1
XDFFPOSX1_43 INVX2_1/A CLKBUF1_9/Y AOI21X1_17/Y gnd vdd DFFPOSX1
XAOI22X1_18 INVX1_124/Y INVX1_117/A OR2X2_14/B INVX1_125/Y gnd OR2X2_16/A vdd AOI22X1
XMUX2X1_3 MUX2X1_4/A MUX2X1_4/B MUX2X1_3/S gnd MUX2X1_3/Y vdd MUX2X1
XXOR2X1_14 block11[0] block6[0] gnd XOR2X1_14/Y vdd XOR2X1
XNAND3X1_45 OR2X2_22/A INVX4_2/Y INVX2_14/Y gnd NOR2X1_189/B vdd NAND3X1
XINVX1_219 OR2X2_5/B gnd INVX1_219/Y vdd INVX1
XCLKBUF1_4 clk gnd CLKBUF1_4/Y vdd CLKBUF1
XINVX1_65 INVX1_65/A gnd INVX1_65/Y vdd INVX1
XINVX1_183 INVX1_183/A gnd INVX1_183/Y vdd INVX1
XINVX1_147 INVX1_110/A gnd INVX1_147/Y vdd INVX1
XINVX1_29 BUFX2_5/A gnd INVX1_29/Y vdd INVX1
XINVX1_111 XOR2X1_9/A gnd INVX1_111/Y vdd INVX1
XAOI22X1_9 INVX1_54/Y gnd INVX1_55/Y gnd gnd AND2X2_5/B vdd AOI22X1
XBUFX4_36 BUFX4_35/A gnd BUFX4_36/Y vdd BUFX4
XAND2X2_15 AND2X2_15/A AND2X2_15/B gnd AND2X2_15/Y vdd AND2X2
XFILL_12_3_1 gnd vdd FILL
XFILL_14_1_0 gnd vdd FILL
XNOR2X1_90 INVX1_115/Y OR2X2_11/A gnd NOR2X1_90/Y vdd NOR2X1
XNOR2X1_18 INVX1_20/Y NOR2X1_6/B gnd NOR2X1_18/Y vdd NOR2X1
XNOR2X1_54 target[3] gnd gnd INVX1_84/A vdd NOR2X1
XXNOR2X1_9 target[6] gnd gnd XNOR2X1_9/Y vdd XNOR2X1
XFILL_1_2_0 gnd vdd FILL
XOAI21X1_146 NAND3X1_43/Y INVX4_3/Y INVX1_178/A gnd AOI21X1_99/A vdd OAI21X1
XOAI21X1_110 INVX1_176/Y INVX1_157/Y INVX1_177/Y gnd OAI21X1_111/B vdd OAI21X1
XNOR2X1_179 NOR2X1_179/A NOR2X1_179/B gnd NOR2X1_179/Y vdd NOR2X1
XXNOR2X1_17 INVX1_110/A INVX1_98/A gnd NAND2X1_74/A vdd XNOR2X1
XNOR2X1_107 INVX1_117/A INVX1_124/Y gnd OR2X2_16/B vdd NOR2X1
XNOR2X1_143 XOR2X1_12/A BUFX4_33/Y gnd NOR2X1_143/Y vdd NOR2X1
XAOI21X1_86 MUX2X1_3/Y AOI21X1_86/B INVX1_189/Y gnd AOI21X1_86/Y vdd AOI21X1
XNAND2X1_152 AND2X2_3/B AND2X2_2/A gnd NOR3X1_8/B vdd NAND2X1
XOAI21X1_3 BUFX4_24/Y BUFX4_5/Y XOR2X1_9/B gnd OAI21X1_3/Y vdd OAI21X1
XAOI21X1_50 INVX2_6/Y INVX1_98/Y OAI21X1_58/Y gnd AOI21X1_50/Y vdd AOI21X1
XNAND2X1_116 INVX1_188/Y NOR2X1_172/Y gnd INVX1_190/A vdd NAND2X1
XFILL_8_2_0 gnd vdd FILL
XINVX8_3 INVX8_3/A gnd INVX8_3/Y vdd INVX8
XOAI21X1_98 INVX1_165/Y INVX4_1/Y INVX1_151/A gnd OAI21X1_98/Y vdd OAI21X1
XBUFX2_17 BUFX2_17/A gnd nonce1[7] vdd BUFX2
XDFFPOSX1_146 INVX1_204/A CLKBUF1_2/Y MUX2X1_5/Y gnd vdd DFFPOSX1
XNAND2X1_77 INVX2_6/A INVX1_148/Y gnd AOI21X1_64/B vdd NAND2X1
XOAI21X1_62 NOR2X1_73/A XOR2X1_8/B NOR2X1_70/Y gnd NOR2X1_74/B vdd OAI21X1
XAOI21X1_14 AOI21X1_14/A AOI21X1_14/B BUFX4_1/Y gnd AOI21X1_14/Y vdd AOI21X1
XDFFPOSX1_80 OR2X2_14/B CLKBUF1_8/Y OR2X2_14/Y gnd vdd DFFPOSX1
XNAND2X1_41 gnd INVX1_87/Y gnd NAND2X1_41/Y vdd NAND2X1
XDFFPOSX1_44 INVX2_6/A CLKBUF1_5/Y AOI21X1_1/Y gnd vdd DFFPOSX1
XOAI21X1_26 NAND2X1_7/Y INVX1_38/A BUFX4_45/Y gnd NOR2X1_31/A vdd OAI21X1
XDFFPOSX1_110 BUFX4_18/A CLKBUF1_7/Y AOI21X1_84/Y gnd vdd DFFPOSX1
XAOI22X1_19 INVX1_128/Y OR2X2_13/B OR2X2_12/B INVX1_129/Y gnd NAND3X1_34/C vdd AOI22X1
XMUX2X1_4 MUX2X1_4/A MUX2X1_4/B MUX2X1_4/S gnd MUX2X1_4/Y vdd MUX2X1
XXOR2X1_15 block10[0] block5[0] gnd XOR2X1_15/Y vdd XOR2X1
XINVX1_220 NOR2X1_1/A gnd NAND2X1_4/A vdd INVX1
XNAND3X1_46 INVX1_198/Y XOR2X1_14/Y INVX1_199/Y gnd AOI21X1_98/B vdd NAND3X1
XNAND3X1_10 NAND3X1_10/A BUFX4_27/Y BUFX4_15/Y gnd NAND3X1_10/Y vdd NAND3X1
XCLKBUF1_5 clk gnd CLKBUF1_5/Y vdd CLKBUF1
XINVX1_66 INVX1_66/A gnd INVX1_66/Y vdd INVX1
XINVX1_184 AND2X2_16/Y gnd INVX1_184/Y vdd INVX1
XINVX1_148 INVX1_148/A gnd INVX1_148/Y vdd INVX1
XINVX1_30 BUFX2_6/A gnd INVX1_30/Y vdd INVX1
XINVX1_112 INVX1_135/A gnd INVX1_112/Y vdd INVX1
XAOI21X1_100 NOR2X1_187/Y XOR2X1_16/Y AOI21X1_100/C gnd AOI21X1_100/Y vdd AOI21X1
XBUFX4_37 BUFX4_38/A gnd NOR2X1_5/B vdd BUFX4
XFILL_14_1_1 gnd vdd FILL
XNOR2X1_91 INVX1_116/Y BUFX4_9/Y gnd NOR2X1_91/Y vdd NOR2X1
XAND2X2_16 INVX2_12/Y AND2X2_15/B gnd AND2X2_16/Y vdd AND2X2
XNOR2X1_55 target[1] INVX1_85/Y gnd NOR2X1_55/Y vdd NOR2X1
XFILL_3_0_0 gnd vdd FILL
XNOR2X1_19 INVX1_21/Y NOR2X1_3/B gnd NOR2X1_19/Y vdd NOR2X1
XFILL_1_2_1 gnd vdd FILL
XOAI21X1_147 NOR2X1_182/B INVX4_3/Y INVX1_200/Y gnd NAND2X1_137/B vdd OAI21X1
XNOR2X1_180 NOR2X1_180/A NOR2X1_179/B gnd NOR2X1_180/Y vdd NOR2X1
XXNOR2X1_18 INVX1_148/A INVX2_6/A gnd NAND2X1_74/B vdd XNOR2X1
XOAI21X1_111 AOI21X1_73/Y OAI21X1_111/B OAI21X1_108/Y gnd OAI21X1_113/A vdd OAI21X1
XNOR2X1_144 NOR2X1_143/Y INVX1_168/Y gnd AOI21X1_71/B vdd NOR2X1
XAOI21X1_87 MUX2X1_4/Y AOI21X1_87/B INVX1_189/Y gnd AOI21X1_87/Y vdd AOI21X1
XNOR2X1_108 NOR2X1_108/A AOI21X1_62/Y gnd OAI21X1_79/C vdd NOR2X1
XAOI21X1_51 INVX2_6/A INVX1_98/A XOR2X1_9/B gnd NOR2X1_71/A vdd AOI21X1
XINVX8_4 INVX8_4/A gnd BUFX4_3/A vdd INVX8
XOAI21X1_4 BUFX4_23/Y BUFX4_7/Y INVX2_7/A gnd AOI21X1_4/B vdd OAI21X1
XFILL_8_2_1 gnd vdd FILL
XNAND2X1_117 INVX1_86/A INVX1_190/Y gnd AOI21X1_86/B vdd NAND2X1
XAOI21X1_15 AOI21X1_15/A AOI21X1_15/B BUFX4_1/Y gnd AOI21X1_15/Y vdd AOI21X1
XOAI21X1_99 OAI21X1_98/Y NOR2X1_137/Y INVX1_164/Y gnd OAI21X1_99/Y vdd OAI21X1
XNAND2X1_78 AND2X2_15/A NOR2X1_112/Y gnd NAND2X1_78/Y vdd NAND2X1
XBUFX2_18 INVX1_9/A gnd nonce2[0] vdd BUFX2
XOAI21X1_63 INVX1_101/Y XOR2X1_7/A NOR2X1_70/Y gnd NOR2X1_76/B vdd OAI21X1
XDFFPOSX1_45 INVX1_98/A CLKBUF1_9/Y AOI21X1_2/Y gnd vdd DFFPOSX1
XDFFPOSX1_81 INVX1_117/A CLKBUF1_9/Y NOR2X1_92/Y gnd vdd DFFPOSX1
XNAND2X1_42 XNOR2X1_8/Y XNOR2X1_9/Y gnd NOR2X1_65/B vdd NAND2X1
XOAI21X1_27 NAND2X1_7/Y INVX1_38/A INVX1_37/A gnd OAI21X1_27/Y vdd OAI21X1
XDFFPOSX1_147 INVX1_18/A CLKBUF1_11/Y NOR3X1_7/Y gnd vdd DFFPOSX1
XAOI22X1_20 INVX1_132/Y INVX1_134/A INVX1_135/A INVX1_133/Y gnd AND2X2_12/A vdd AOI22X1
XDFFPOSX1_111 OR2X2_1/B CLKBUF1_3/Y AOI21X1_87/Y gnd vdd DFFPOSX1
XMUX2X1_5 MUX2X1_7/A MUX2X1_5/B MUX2X1_5/S gnd MUX2X1_5/Y vdd MUX2X1
XCLKBUF1_6 clk gnd CLKBUF1_6/Y vdd CLKBUF1
XINVX1_67 target[1] gnd INVX1_67/Y vdd INVX1
XNAND3X1_47 INVX4_2/Y NOR2X1_184/Y INVX4_3/A gnd AND2X2_31/A vdd NAND3X1
XINVX1_185 OR2X2_23/A gnd INVX1_185/Y vdd INVX1
XXOR2X1_16 XOR2X1_16/A block4[0] gnd XOR2X1_16/Y vdd XOR2X1
XINVX1_221 NAND2X1_6/A gnd AND2X2_2/A vdd INVX1
XFILL_1_1 gnd vdd FILL
XNAND3X1_11 NAND3X1_11/A BUFX4_26/Y BUFX4_16/Y gnd AOI21X1_11/A vdd NAND3X1
XINVX1_149 OR2X2_22/B gnd INVX1_149/Y vdd INVX1
XINVX1_31 BUFX2_7/A gnd INVX1_31/Y vdd INVX1
XINVX1_113 INVX1_134/A gnd NOR2X1_88/A vdd INVX1
XAOI21X1_101 NOR2X1_189/Y XOR2X1_17/Y NAND2X1_138/Y gnd AOI21X1_101/Y vdd AOI21X1
XBUFX4_38 BUFX4_38/A gnd NOR2X1_6/B vdd BUFX4
XNOR2X1_92 INVX1_117/Y BUFX4_11/Y gnd NOR2X1_92/Y vdd NOR2X1
XAND2X2_17 BUFX4_32/Y block10[0] gnd AND2X2_17/Y vdd AND2X2
XNOR2X1_56 target[0] INVX1_86/Y gnd NOR2X1_56/Y vdd NOR2X1
XFILL_15_2_0 gnd vdd FILL
XNOR2X1_20 INVX1_22/Y NOR2X1_5/B gnd NOR2X1_20/Y vdd NOR2X1
XFILL_3_0_1 gnd vdd FILL
XOAI21X1_148 NOR2X1_189/B INVX4_3/Y INVX1_201/Y gnd NAND2X1_138/B vdd OAI21X1
XNOR2X1_181 INVX1_198/A NAND3X1_43/Y gnd NOR2X1_181/Y vdd NOR2X1
XOAI21X1_112 AND2X2_14/Y NOR2X1_126/Y INVX1_178/Y gnd NAND3X1_37/B vdd OAI21X1
XNOR2X1_145 NOR3X1_4/A NOR2X1_168/B gnd INVX1_169/A vdd NOR2X1
XNOR2X1_109 NOR2X1_109/A NAND2X1_70/Y gnd NOR2X1_109/Y vdd NOR2X1
XFILL_2_3_0 gnd vdd FILL
XAOI21X1_88 AND2X2_28/Y AOI21X1_88/B AOI21X1_88/C gnd AOI21X1_88/Y vdd AOI21X1
XXNOR2X1_19 INVX4_1/A block2[0] gnd XNOR2X1_19/Y vdd XNOR2X1
XAOI21X1_52 INVX2_7/Y NOR3X1_1/C OAI21X1_59/Y gnd AOI21X1_52/Y vdd AOI21X1
XBUFX2_19 BUFX2_19/A gnd nonce2[1] vdd BUFX2
XOAI21X1_5 BUFX4_24/Y BUFX4_5/Y INVX1_99/A gnd AOI21X1_5/B vdd OAI21X1
XNAND2X1_118 OR2X2_1/B INVX1_190/Y gnd AOI21X1_87/B vdd NAND2X1
XAOI21X1_16 AOI21X1_16/A OAI21X1_16/Y BUFX4_1/Y gnd AOI21X1_16/Y vdd AOI21X1
XFILL_14_1 gnd vdd FILL
XOAI21X1_64 NOR2X1_75/Y INVX1_103/A NOR2X1_70/Y gnd NOR2X1_77/B vdd OAI21X1
XFILL_9_3_0 gnd vdd FILL
XDFFPOSX1_82 INVX1_118/A CLKBUF1_8/Y NOR2X1_93/Y gnd vdd DFFPOSX1
XNAND2X1_79 INVX2_11/Y INVX2_10/Y gnd INVX2_12/A vdd NAND2X1
XAOI22X1_21 INVX1_134/Y OAI22X1_5/B OAI22X1_5/C INVX1_99/A gnd AND2X2_12/B vdd AOI22X1
XDFFPOSX1_46 XOR2X1_9/B CLKBUF1_1/Y AOI21X1_3/Y gnd vdd DFFPOSX1
XDFFPOSX1_112 INVX1_86/A CLKBUF1_4/Y AOI21X1_86/Y gnd vdd DFFPOSX1
XOAI21X1_28 start NAND2X1_1/B BUFX4_45/Y gnd NOR2X1_33/A vdd OAI21X1
XNAND2X1_43 INVX1_217/A INVX1_92/Y gnd AOI22X1_16/A vdd NAND2X1
XDFFPOSX1_10 INVX1_37/A CLKBUF1_9/Y AOI21X1_28/Y gnd vdd DFFPOSX1
XMUX2X1_6 INVX2_18/Y MUX2X1_7/A MUX2X1_6/S gnd MUX2X1_6/Y vdd MUX2X1
XINVX1_68 target[0] gnd INVX1_68/Y vdd INVX1
XXOR2X1_17 XOR2X1_17/A block3[0] gnd XOR2X1_17/Y vdd XOR2X1
XINVX1_222 start gnd NOR2X1_32/A vdd INVX1
XNAND3X1_48 NAND2X1_1/A NAND2X1_1/B NAND2X1_4/A gnd NOR3X1_8/A vdd NAND3X1
XCLKBUF1_7 clk gnd CLKBUF1_7/Y vdd CLKBUF1
XNAND3X1_12 NAND3X1_12/A BUFX4_26/Y BUFX4_14/Y gnd AOI21X1_12/A vdd NAND3X1
XINVX1_186 BUFX4_18/Y gnd INVX1_186/Y vdd INVX1
XFILL_10_0_0 gnd vdd FILL
XINVX1_32 BUFX2_8/A gnd INVX1_32/Y vdd INVX1
XINVX1_114 XOR2X1_8/A gnd NOR2X1_89/A vdd INVX1
XAOI21X1_102 AOI21X1_102/A AOI21X1_102/B AND2X2_31/A gnd NOR3X1_6/A vdd AOI21X1
XINVX1_150 OR2X2_23/A gnd INVX1_150/Y vdd INVX1
XBUFX4_39 BUFX4_38/A gnd BUFX4_39/Y vdd BUFX4
XNOR2X1_93 NOR2X1_93/A BUFX4_9/Y gnd NOR2X1_93/Y vdd NOR2X1
XAND2X2_18 BUFX4_33/Y XOR2X1_11/A gnd AND2X2_18/Y vdd AND2X2
XNOR2X1_57 gnd INVX1_87/Y gnd NOR2X1_57/Y vdd NOR2X1
XNOR2X1_21 INVX1_23/Y NOR2X1_5/B gnd NOR2X1_21/Y vdd NOR2X1
XFILL_17_0_0 gnd vdd FILL
XFILL_15_2_1 gnd vdd FILL
XOAI21X1_149 XOR2X1_12/A block7[0] block2[0] gnd AOI21X1_102/A vdd OAI21X1
XNOR2X1_182 INVX1_198/A NOR2X1_182/B gnd NOR2X1_182/Y vdd NOR2X1
XOAI21X1_113 OAI21X1_113/A INVX1_173/Y NAND3X1_37/Y gnd OAI21X1_113/Y vdd OAI21X1
XNOR2X1_146 XOR2X1_11/A BUFX4_33/Y gnd NOR2X1_146/Y vdd NOR2X1
XNOR2X1_110 NOR2X1_110/A OAI21X1_82/A gnd NOR2X1_110/Y vdd NOR2X1
XFILL_2_3_1 gnd vdd FILL
XFILL_4_1_0 gnd vdd FILL
XXNOR2X1_20 BUFX4_34/Y block4[0] gnd MUX2X1_1/B vdd XNOR2X1
XAOI21X1_89 AOI21X1_89/A AOI21X1_89/B INVX8_3/Y gnd AOI21X1_89/Y vdd AOI21X1
XAOI21X1_53 INVX1_124/A NOR3X1_3/Y OAI21X1_69/Y gnd AOI21X1_53/Y vdd AOI21X1
XOAI21X1_6 BUFX4_24/Y BUFX4_5/Y OAI22X1_5/B gnd OAI21X1_6/Y vdd OAI21X1
XNAND2X1_119 INVX1_39/A INVX1_193/Y gnd NAND2X1_119/Y vdd NAND2X1
XAOI21X1_17 INVX2_1/Y AOI22X1_1/B OR2X2_1/A gnd AOI21X1_17/Y vdd AOI21X1
XOAI21X1_65 NOR3X1_2/Y OAI22X1_6/B NOR2X1_70/Y gnd NOR2X1_78/A vdd OAI21X1
XDFFPOSX1_83 INVX2_8/A CLKBUF1_5/Y NOR2X1_94/Y gnd vdd DFFPOSX1
XFILL_9_3_1 gnd vdd FILL
XFILL_14_2 gnd vdd FILL
XNAND2X1_80 NOR2X1_112/Y INVX2_12/Y gnd NAND2X1_80/Y vdd NAND2X1
XBUFX2_20 INVX1_11/A gnd nonce2[2] vdd BUFX2
XDFFPOSX1_47 INVX2_7/A CLKBUF1_1/Y AOI21X1_4/Y gnd vdd DFFPOSX1
XDFFPOSX1_113 AND2X2_30/B CLKBUF1_7/Y AOI21X1_85/Y gnd vdd DFFPOSX1
XOAI21X1_29 INVX2_1/Y INVX1_39/Y NOR2X1_33/B gnd OAI21X1_29/Y vdd OAI21X1
XNAND2X1_44 AND2X2_7/B AND2X2_7/A gnd OAI21X1_54/A vdd NAND2X1
XAOI22X1_22 AOI22X1_22/A AND2X2_13/A OAI21X1_75/Y OAI21X1_83/C gnd AOI22X1_22/Y vdd
+ AOI22X1
XDFFPOSX1_11 BUFX2_2/A CLKBUF1_12/Y AOI22X1_4/Y gnd vdd DFFPOSX1
XMUX2X1_7 MUX2X1_7/A MUX2X1_7/B MUX2X1_7/S gnd MUX2X1_7/Y vdd MUX2X1
XNAND3X1_49 NAND3X1_49/A BUFX4_27/Y BUFX4_13/Y gnd AOI21X1_1/A vdd NAND3X1
XINVX1_187 INVX1_187/A gnd INVX1_187/Y vdd INVX1
XNAND3X1_13 NAND3X1_13/A BUFX4_26/Y BUFX4_14/Y gnd NAND3X1_13/Y vdd NAND3X1
XCLKBUF1_8 clk gnd CLKBUF1_8/Y vdd CLKBUF1
XINVX1_69 gnd gnd INVX1_69/Y vdd INVX1
XFILL_10_0_1 gnd vdd FILL
XINVX1_151 INVX1_151/A gnd INVX1_151/Y vdd INVX1
XINVX1_33 BUFX2_9/A gnd INVX1_33/Y vdd INVX1
XAOI21X1_103 AOI21X1_103/A AOI21X1_103/B INVX8_3/Y gnd AOI21X1_103/Y vdd AOI21X1
XINVX1_115 INVX2_9/A gnd INVX1_115/Y vdd INVX1
XNOR2X1_94 NOR2X1_94/A BUFX4_11/Y gnd NOR2X1_94/Y vdd NOR2X1
XAND2X2_19 BUFX4_31/Y AND2X2_19/B gnd OAI22X1_8/A vdd AND2X2
XBUFX4_40 BUFX4_38/A gnd NOR2X1_3/B vdd BUFX4
XNOR2X1_58 gnd INVX1_88/Y gnd NOR2X1_58/Y vdd NOR2X1
XNOR2X1_22 INVX1_24/Y NOR2X1_5/B gnd NOR2X1_22/Y vdd NOR2X1
XFILL_17_0_1 gnd vdd FILL
XNOR2X1_183 INVX1_198/A NOR2X1_189/B gnd NOR2X1_183/Y vdd NOR2X1
XCLKBUF1_10 clk gnd CLKBUF1_10/Y vdd CLKBUF1
XOAI21X1_150 NAND3X1_41/Y NOR2X1_192/A NOR2X1_169/A gnd AOI21X1_103/A vdd OAI21X1
XOAI21X1_114 INVX1_179/Y NOR2X1_158/Y NOR2X1_155/Y gnd OAI21X1_115/C vdd OAI21X1
XNOR2X1_147 INVX1_170/Y INVX4_1/Y gnd NOR2X1_147/Y vdd NOR2X1
XFILL_16_3_0 gnd vdd FILL
XNOR2X1_111 INVX1_98/A INVX1_147/Y gnd AOI21X1_64/C vdd NOR2X1
XFILL_4_1_1 gnd vdd FILL
XXNOR2X1_21 BUFX4_34/Y block5[0] gnd XNOR2X1_21/Y vdd XNOR2X1
XAOI21X1_54 INVX1_124/A NOR3X1_3/Y INVX1_122/A gnd NOR2X1_83/A vdd AOI21X1
XAOI21X1_90 AOI21X1_90/A AOI21X1_90/B INVX8_3/Y gnd AOI21X1_90/Y vdd AOI21X1
XOAI21X1_7 BUFX4_24/Y BUFX4_5/Y XOR2X1_8/B gnd AOI21X1_7/B vdd OAI21X1
XNAND2X1_120 INVX1_39/A INVX1_194/Y gnd NAND2X1_120/Y vdd NAND2X1
XAOI21X1_18 INVX1_27/Y AOI22X1_1/B OR2X2_1/A gnd AOI21X1_18/Y vdd AOI21X1
XDFFPOSX1_84 NAND3X1_49/A CLKBUF1_9/Y AND2X2_10/Y gnd vdd DFFPOSX1
XOAI21X1_66 INVX1_104/Y OR2X2_15/B NOR2X1_70/Y gnd NOR2X1_79/B vdd OAI21X1
XNAND2X1_81 AND2X2_15/A NOR2X1_116/Y gnd NOR2X1_117/B vdd NAND2X1
XBUFX2_21 INVX1_12/A gnd nonce2[3] vdd BUFX2
XDFFPOSX1_48 INVX1_99/A CLKBUF1_6/Y AOI21X1_5/Y gnd vdd DFFPOSX1
XDFFPOSX1_114 INVX1_188/A CLKBUF1_7/Y NAND2X1_115/Y gnd vdd DFFPOSX1
XOAI21X1_30 start INVX1_39/A BUFX4_45/Y gnd AOI21X1_30/C vdd OAI21X1
XNAND2X1_45 AND2X2_8/A AND2X2_8/B gnd NOR2X1_65/A vdd NAND2X1
XAOI22X1_23 XOR2X1_12/A AOI22X1_23/B INVX1_210/Y AOI22X1_23/D gnd AOI22X1_23/Y vdd
+ AOI22X1
XDFFPOSX1_12 BUFX2_3/A CLKBUF1_12/Y AOI21X1_18/Y gnd vdd DFFPOSX1
XINVX1_188 INVX1_188/A gnd INVX1_188/Y vdd INVX1
XCLKBUF1_9 clk gnd CLKBUF1_9/Y vdd CLKBUF1
XNAND3X1_14 NAND3X1_14/A INVX8_1/A BUFX4_14/Y gnd AOI21X1_14/A vdd NAND3X1
XINVX1_70 gnd gnd INVX1_70/Y vdd INVX1
XAOI21X1_104 OAI21X1_158/C INVX1_215/A XOR2X1_13/A gnd NOR2X1_203/A vdd AOI21X1
XINVX1_152 INVX1_152/A gnd INVX1_152/Y vdd INVX1
XINVX1_34 INVX1_34/A gnd INVX1_34/Y vdd INVX1
XBUFX4_41 reset gnd BUFX2_34/A vdd BUFX4
XINVX1_116 INVX1_143/A gnd INVX1_116/Y vdd INVX1
XAND2X2_20 BUFX4_31/Y AND2X2_20/B gnd AND2X2_20/Y vdd AND2X2
XNOR2X1_95 NOR2X1_95/A NOR2X1_95/B gnd AND2X2_11/B vdd NOR2X1
XFILL_11_1_0 gnd vdd FILL
XNOR2X1_23 INVX1_25/Y NOR2X1_5/B gnd NOR2X1_23/Y vdd NOR2X1
XNOR2X1_59 gnd INVX1_89/Y gnd NOR2X1_59/Y vdd NOR2X1
XOAI21X1_151 INVX2_19/Y INVX4_4/Y INVX4_5/A gnd AOI22X1_23/B vdd OAI21X1
XFILL_5_1 gnd vdd FILL
XCLKBUF1_11 clk gnd CLKBUF1_11/Y vdd CLKBUF1
XNOR2X1_184 OR2X2_23/B OR2X2_22/A gnd NOR2X1_184/Y vdd NOR2X1
XOAI21X1_115 OAI21X1_113/Y NOR2X1_155/Y OAI21X1_115/C gnd MUX2X1_2/A vdd OAI21X1
XNOR2X1_148 NOR2X1_168/B NOR2X1_147/Y gnd AOI21X1_72/B vdd NOR2X1
XFILL_16_3_1 gnd vdd FILL
XXNOR2X1_22 BUFX4_36/Y XNOR2X1_22/B gnd MUX2X1_2/B vdd XNOR2X1
XNOR2X1_112 INVX1_149/Y INVX1_150/Y gnd NOR2X1_112/Y vdd NOR2X1
XAOI21X1_91 AOI21X1_91/A AOI21X1_91/B INVX8_3/Y gnd AOI21X1_91/Y vdd AOI21X1
XFILL_5_2_0 gnd vdd FILL
XOAI21X1_8 BUFX4_25/Y BUFX4_5/Y XOR2X1_7/A gnd AOI21X1_8/B vdd OAI21X1
XAOI21X1_55 INVX1_108/Y NAND2X1_56/B OAI21X1_70/Y gnd AOI21X1_55/Y vdd AOI21X1
XNAND2X1_121 OR2X2_23/B OR2X2_22/A gnd NOR2X1_177/A vdd NAND2X1
XDFFPOSX1_85 NAND3X1_2/A CLKBUF1_9/Y AOI21X1_50/Y gnd vdd DFFPOSX1
XOAI21X1_67 NOR2X1_79/A INVX1_106/A NOR2X1_70/Y gnd NOR2X1_81/B vdd OAI21X1
XNAND2X1_82 NOR2X1_116/Y INVX2_12/Y gnd NOR2X1_118/B vdd NAND2X1
XBUFX2_22 INVX1_13/A gnd nonce2[4] vdd BUFX2
XAOI21X1_19 INVX1_28/Y AOI22X1_1/B OR2X2_1/A gnd AOI21X1_19/Y vdd AOI21X1
XDFFPOSX1_115 AND2X2_28/B CLKBUF1_4/Y AND2X2_29/Y gnd vdd DFFPOSX1
XOAI21X1_31 start INVX1_120/A INVX8_4/A gnd AOI21X1_31/C vdd OAI21X1
XDFFPOSX1_49 OAI22X1_5/B CLKBUF1_1/Y AOI21X1_6/Y gnd vdd DFFPOSX1
XNAND2X1_46 XNOR2X1_11/Y NAND2X1_46/B gnd NOR2X1_66/A vdd NAND2X1
XNAND2X1_10 target[15] INVX1_41/Y gnd NAND3X1_19/A vdd NAND2X1
XDFFPOSX1_13 BUFX2_4/A CLKBUF1_11/Y AOI21X1_19/Y gnd vdd DFFPOSX1
XINVX1_189 BUFX2_34/A gnd INVX1_189/Y vdd INVX1
XNAND3X1_15 NAND3X1_15/A INVX8_1/A BUFX4_14/Y gnd AOI21X1_15/A vdd NAND3X1
XFILL_18_1 gnd vdd FILL
XINVX1_71 target[14] gnd INVX1_71/Y vdd INVX1
XINVX1_153 INVX1_153/A gnd MUX2X1_1/S vdd INVX1
XINVX1_35 INVX1_35/A gnd INVX1_35/Y vdd INVX1
XAOI21X1_105 INVX1_213/Y INVX1_214/Y INVX2_17/Y gnd AOI21X1_105/Y vdd AOI21X1
XINVX1_117 INVX1_117/A gnd INVX1_117/Y vdd INVX1
XBUFX4_42 reset gnd INVX8_3/A vdd BUFX4
XNOR2X1_96 NOR2X1_96/A NOR2X1_96/B gnd AND2X2_11/A vdd NOR2X1
XFILL_11_1_1 gnd vdd FILL
XAND2X2_21 BUFX4_30/Y AND2X2_21/B gnd AND2X2_21/Y vdd AND2X2
XNOR2X1_60 gnd INVX1_90/Y gnd NOR2X1_60/Y vdd NOR2X1
XCLKBUF1_12 clk gnd CLKBUF1_12/Y vdd CLKBUF1
XNOR2X1_24 NOR2X1_24/A INVX1_34/Y gnd NOR2X1_24/Y vdd NOR2X1
XFILL_0_0_0 gnd vdd FILL
XOAI21X1_152 MUX2X1_7/B INVX1_208/Y AOI22X1_23/Y gnd AND2X2_32/A vdd OAI21X1
XNOR2X1_185 OR2X2_22/B OR2X2_23/A gnd INVX4_3/A vdd NOR2X1
XOAI21X1_116 MUX2X1_2/Y AOI21X1_74/A AOI21X1_74/Y gnd OAI21X1_116/Y vdd OAI21X1
XXNOR2X1_23 BUFX4_36/Y XNOR2X1_23/B gnd XNOR2X1_23/Y vdd XNOR2X1
XNOR2X1_149 BUFX4_48/Y NOR2X1_149/B gnd INVX1_171/A vdd NOR2X1
XNOR2X1_113 OR2X2_23/B INVX2_10/Y gnd AND2X2_15/A vdd NOR2X1
XAOI21X1_92 AOI21X1_92/A AOI21X1_92/B INVX8_3/Y gnd AOI21X1_92/Y vdd AOI21X1
XAOI21X1_56 INVX1_120/Y NAND2X1_57/Y AOI21X1_56/C gnd AOI21X1_56/Y vdd AOI21X1
XOAI21X1_9 BUFX4_25/Y BUFX4_8/Y INVX1_103/A gnd OAI21X1_9/Y vdd OAI21X1
XFILL_7_0_0 gnd vdd FILL
XNAND2X1_122 OR2X2_22/A INVX2_14/Y gnd NOR2X1_179/A vdd NAND2X1
XBUFX2_23 BUFX2_23/A gnd nonce2[5] vdd BUFX2
XFILL_5_2_1 gnd vdd FILL
XNAND2X1_83 NOR2X1_120/Y NAND2X1_83/B gnd NOR2X1_159/B vdd NAND2X1
XAOI21X1_20 INVX1_29/Y AOI22X1_1/B OR2X2_1/A gnd AOI21X1_20/Y vdd AOI21X1
XOAI21X1_32 NOR2X1_38/Y NOR2X1_39/Y OAI21X1_32/C gnd NAND2X1_20/A vdd OAI21X1
XDFFPOSX1_50 XOR2X1_8/B CLKBUF1_1/Y AOI21X1_7/Y gnd vdd DFFPOSX1
XDFFPOSX1_86 NAND3X1_3/A CLKBUF1_1/Y NOR2X1_71/Y gnd vdd DFFPOSX1
XOAI21X1_68 NOR2X1_81/A INVX1_107/A NOR2X1_70/Y gnd NOR2X1_82/B vdd OAI21X1
XNAND2X1_47 NOR2X1_65/Y NOR2X1_66/Y gnd NAND2X1_47/Y vdd NAND2X1
XBUFX2_1 INVX2_1/A gnd finish vdd BUFX2
XDFFPOSX1_116 AND2X2_14/B CLKBUF1_4/Y AOI21X1_88/Y gnd vdd DFFPOSX1
XDFFPOSX1_14 BUFX2_5/A CLKBUF1_11/Y AOI21X1_20/Y gnd vdd DFFPOSX1
XNAND2X1_11 target[14] INVX1_42/Y gnd NAND3X1_19/B vdd NAND2X1
XINVX1_190 INVX1_190/A gnd INVX1_190/Y vdd INVX1
XINVX1_72 gnd gnd INVX1_72/Y vdd INVX1
XINVX1_154 INVX1_154/A gnd INVX1_154/Y vdd INVX1
XNAND3X1_16 NAND3X1_16/A INVX8_1/A BUFX4_13/Y gnd AOI21X1_16/A vdd NAND3X1
XINVX1_36 INVX1_36/A gnd INVX1_36/Y vdd INVX1
XAOI21X1_106 INVX4_4/Y INVX2_17/A INVX1_212/A gnd AOI21X1_106/Y vdd AOI21X1
XINVX1_118 INVX1_118/A gnd NOR2X1_93/A vdd INVX1
XBUFX4_43 reset gnd OR2X2_8/A vdd BUFX4
XNOR2X1_97 XOR2X1_7/Y XOR2X1_8/Y gnd NOR2X1_97/Y vdd NOR2X1
XAND2X2_22 BUFX4_30/Y INVX1_195/A gnd AND2X2_22/Y vdd AND2X2
XNOR2X1_61 gnd INVX1_91/Y gnd NOR2X1_61/Y vdd NOR2X1
XINVX2_10 OR2X2_22/A gnd INVX2_10/Y vdd INVX2
XFILL_12_2_0 gnd vdd FILL
XNOR2X1_25 BUFX4_6/Y BUFX4_22/Y gnd NOR2X1_25/Y vdd NOR2X1
XFILL_0_0_1 gnd vdd FILL
XOAI21X1_153 INVX4_5/Y gnd gnd gnd OAI21X1_158/C vdd OAI21X1
XNOR2X1_186 INVX4_3/Y NAND3X1_43/Y gnd NOR2X1_186/Y vdd NOR2X1
XOAI21X1_117 OAI21X1_142/C BUFX4_36/Y AOI21X1_74/C gnd OAI21X1_117/Y vdd OAI21X1
XNOR2X1_150 BUFX4_47/Y NAND2X1_96/Y gnd NOR2X1_150/Y vdd NOR2X1
XAOI21X1_93 AOI21X1_93/A AOI21X1_93/B INVX8_3/Y gnd AOI21X1_93/Y vdd AOI21X1
XXNOR2X1_24 BUFX4_31/Y XNOR2X1_24/B gnd XNOR2X1_24/Y vdd XNOR2X1
XNOR2X1_114 NOR3X1_4/A NAND2X1_78/Y gnd NOR2X1_114/Y vdd NOR2X1
XAOI21X1_57 INVX1_136/Y INVX1_145/A XOR2X1_9/Y gnd AOI21X1_57/Y vdd AOI21X1
XOR2X2_10 OR2X2_10/A OR2X2_10/B gnd OR2X2_10/Y vdd OR2X2
XDFFPOSX1_1 INVX1_120/A CLKBUF1_3/Y DFFPOSX1_1/D gnd vdd DFFPOSX1
XFILL_7_0_1 gnd vdd FILL
XBUFX2_24 INVX1_15/A gnd nonce2[6] vdd BUFX2
XAOI21X1_21 INVX1_30/Y AOI22X1_1/B OR2X2_1/A gnd AOI21X1_21/Y vdd AOI21X1
XNAND2X1_123 XOR2X1_11/A NOR2X1_175/Y gnd AOI21X1_89/B vdd NAND2X1
XDFFPOSX1_87 NAND3X1_4/A CLKBUF1_3/Y AOI21X1_52/Y gnd vdd DFFPOSX1
XOAI21X1_69 NOR3X1_3/Y INVX1_124/A NOR2X1_70/Y gnd OAI21X1_69/Y vdd OAI21X1
XNAND2X1_84 AND2X2_15/A NOR2X1_120/Y gnd NAND2X1_84/Y vdd NAND2X1
XBUFX2_2 BUFX2_2/A gnd nonce0[0] vdd BUFX2
XDFFPOSX1_117 AND2X2_14/A CLKBUF1_2/Y BUFX2_34/Y gnd vdd DFFPOSX1
XDFFPOSX1_51 XOR2X1_7/A CLKBUF1_1/Y AOI21X1_8/Y gnd vdd DFFPOSX1
XNAND2X1_48 gnd INVX1_95/Y gnd AOI21X1_48/A vdd NAND2X1
XFILL_6_3_0 gnd vdd FILL
XOAI21X1_33 INVX1_52/Y target[5] OAI22X1_1/Y gnd OAI21X1_33/Y vdd OAI21X1
XNAND2X1_12 gnd INVX1_46/Y gnd NAND3X1_20/A vdd NAND2X1
XDFFPOSX1_15 BUFX2_6/A CLKBUF1_11/Y AOI21X1_21/Y gnd vdd DFFPOSX1
XINVX1_73 gnd gnd INVX1_73/Y vdd INVX1
XNAND2X1_1 NAND2X1_1/A NAND2X1_1/B gnd NOR2X1_1/B vdd NAND2X1
XINVX1_191 INVX1_191/A gnd MUX2X1_3/S vdd INVX1
XINVX1_155 INVX1_155/A gnd INVX1_155/Y vdd INVX1
XINVX1_37 INVX1_37/A gnd INVX1_37/Y vdd INVX1
XNAND3X1_17 BUFX4_44/Y NAND2X1_4/Y INVX1_35/A gnd NOR2X1_26/A vdd NAND3X1
XAOI21X1_107 gnd INVX4_5/Y INVX2_17/Y gnd AOI21X1_107/Y vdd AOI21X1
XINVX1_119 INVX2_8/A gnd NOR2X1_94/A vdd INVX1
XBUFX4_44 reset gnd BUFX4_44/Y vdd BUFX4
XNOR2X1_98 OR2X2_10/B INVX2_7/A gnd NOR2X1_98/Y vdd NOR2X1
XAND2X2_23 BUFX4_36/Y INVX1_202/A gnd AND2X2_23/Y vdd AND2X2
.ends

