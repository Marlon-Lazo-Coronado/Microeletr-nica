module area_sys (clk, reset, block0, block1, block2, block3, block4, block5, block6, block7, block8, block9, block10, block11, start, target, nonce0, nonce1, nonce2, nonce3, finish);

input clk;
input reset;
input start;
output finish;
input [7:0] block0;
input [7:0] block1;
input [7:0] block2;
input [7:0] block3;
input [7:0] block4;
input [7:0] block5;
input [7:0] block6;
input [7:0] block7;
input [7:0] block8;
input [7:0] block9;
input [7:0] block10;
input [7:0] block11;
input [15:0] target;
output [7:0] nonce0;
output [7:0] nonce1;
output [7:0] nonce2;
output [7:0] nonce3;

wire vdd = 1'b1;
wire gnd = 1'b0;

BUFX4 BUFX4_1 ( .A(_10_), .Y(_10__bF_buf3) );
BUFX4 BUFX4_2 ( .A(_10_), .Y(_10__bF_buf2) );
BUFX4 BUFX4_3 ( .A(_10_), .Y(_10__bF_buf1) );
BUFX4 BUFX4_4 ( .A(_10_), .Y(_10__bF_buf0) );
CLKBUF1 CLKBUF1_1 ( .A(clk), .Y(clk_bF_buf11) );
CLKBUF1 CLKBUF1_2 ( .A(clk), .Y(clk_bF_buf10) );
CLKBUF1 CLKBUF1_3 ( .A(clk), .Y(clk_bF_buf9) );
CLKBUF1 CLKBUF1_4 ( .A(clk), .Y(clk_bF_buf8) );
CLKBUF1 CLKBUF1_5 ( .A(clk), .Y(clk_bF_buf7) );
CLKBUF1 CLKBUF1_6 ( .A(clk), .Y(clk_bF_buf6) );
CLKBUF1 CLKBUF1_7 ( .A(clk), .Y(clk_bF_buf5) );
CLKBUF1 CLKBUF1_8 ( .A(clk), .Y(clk_bF_buf4) );
CLKBUF1 CLKBUF1_9 ( .A(clk), .Y(clk_bF_buf3) );
CLKBUF1 CLKBUF1_10 ( .A(clk), .Y(clk_bF_buf2) );
CLKBUF1 CLKBUF1_11 ( .A(clk), .Y(clk_bF_buf1) );
CLKBUF1 CLKBUF1_12 ( .A(clk), .Y(clk_bF_buf0) );
BUFX4 BUFX4_5 ( .A(_27_), .Y(_27__bF_buf3) );
BUFX4 BUFX4_6 ( .A(_27_), .Y(_27__bF_buf2) );
BUFX4 BUFX4_7 ( .A(_27_), .Y(_27__bF_buf1) );
BUFX4 BUFX4_8 ( .A(_27_), .Y(_27__bF_buf0) );
BUFX4 BUFX4_9 ( .A(_417_), .Y(_417__bF_buf3) );
BUFX4 BUFX4_10 ( .A(_417_), .Y(_417__bF_buf2) );
BUFX4 BUFX4_11 ( .A(_417_), .Y(_417__bF_buf1) );
BUFX4 BUFX4_12 ( .A(_417_), .Y(_417__bF_buf0) );
BUFX4 BUFX4_13 ( .A(_18_), .Y(_18__bF_buf3) );
BUFX4 BUFX4_14 ( .A(_18_), .Y(_18__bF_buf2) );
BUFX4 BUFX4_15 ( .A(_18_), .Y(_18__bF_buf1) );
BUFX4 BUFX4_16 ( .A(_18_), .Y(_18__bF_buf0) );
BUFX4 BUFX4_17 ( .A(micro_abc_calculation_ints_counter_4_), .Y(micro_abc_calculation_ints_counter_4_bF_buf4_) );
BUFX4 BUFX4_18 ( .A(micro_abc_calculation_ints_counter_4_), .Y(micro_abc_calculation_ints_counter_4_bF_buf3_) );
BUFX4 BUFX4_19 ( .A(micro_abc_calculation_ints_counter_4_), .Y(micro_abc_calculation_ints_counter_4_bF_buf2_) );
BUFX4 BUFX4_20 ( .A(micro_abc_calculation_ints_counter_4_), .Y(micro_abc_calculation_ints_counter_4_bF_buf1_) );
BUFX4 BUFX4_21 ( .A(micro_abc_calculation_ints_counter_4_), .Y(micro_abc_calculation_ints_counter_4_bF_buf0_) );
BUFX4 BUFX4_22 ( .A(_26_), .Y(_26__bF_buf3) );
BUFX4 BUFX4_23 ( .A(_26_), .Y(_26__bF_buf2) );
BUFX4 BUFX4_24 ( .A(_26_), .Y(_26__bF_buf1) );
BUFX4 BUFX4_25 ( .A(_26_), .Y(_26__bF_buf0) );
BUFX4 BUFX4_26 ( .A(_20_), .Y(_20__bF_buf3) );
BUFX4 BUFX4_27 ( .A(_20_), .Y(_20__bF_buf2) );
BUFX4 BUFX4_28 ( .A(_20_), .Y(_20__bF_buf1) );
BUFX4 BUFX4_29 ( .A(_20_), .Y(_20__bF_buf0) );
BUFX4 BUFX4_30 ( .A(_583_), .Y(_583__bF_buf6) );
BUFX4 BUFX4_31 ( .A(_583_), .Y(_583__bF_buf5) );
BUFX4 BUFX4_32 ( .A(_583_), .Y(_583__bF_buf4) );
BUFX4 BUFX4_33 ( .A(_583_), .Y(_583__bF_buf3) );
BUFX4 BUFX4_34 ( .A(_583_), .Y(_583__bF_buf2) );
BUFX4 BUFX4_35 ( .A(_583_), .Y(_583__bF_buf1) );
BUFX4 BUFX4_36 ( .A(_583_), .Y(_583__bF_buf0) );
BUFX4 BUFX4_37 ( .A(_63_), .Y(_63__bF_buf3) );
BUFX4 BUFX4_38 ( .A(_63_), .Y(_63__bF_buf2) );
BUFX4 BUFX4_39 ( .A(_63_), .Y(_63__bF_buf1) );
BUFX4 BUFX4_40 ( .A(_63_), .Y(_63__bF_buf0) );
BUFX4 BUFX4_41 ( .A(reset), .Y(reset_bF_buf5) );
BUFX4 BUFX4_42 ( .A(reset), .Y(reset_bF_buf4) );
BUFX4 BUFX4_43 ( .A(reset), .Y(reset_bF_buf3) );
BUFX4 BUFX4_44 ( .A(reset), .Y(reset_bF_buf2) );
BUFX4 BUFX4_45 ( .A(reset), .Y(reset_bF_buf1) );
BUFX4 BUFX4_46 ( .A(reset), .Y(reset_bF_buf0) );
BUFX4 BUFX4_47 ( .A(_591_), .Y(_591__bF_buf3) );
BUFX4 BUFX4_48 ( .A(_591_), .Y(_591__bF_buf2) );
BUFX4 BUFX4_49 ( .A(_591_), .Y(_591__bF_buf1) );
BUFX4 BUFX4_50 ( .A(_591_), .Y(_591__bF_buf0) );
NAND2X1 NAND2X1_1 ( .A(counter_0_), .B(invalid_nonce), .Y(_22_) );
NOR2X1 NOR2X1_1 ( .A(counter_1_), .B(_22_), .Y(_23_) );
AND2X2 AND2X2_1 ( .A(_13_), .B(_14_), .Y(_24_) );
AND2X2 AND2X2_2 ( .A(_16_), .B(counter_3_), .Y(_25_) );
NAND3X1 NAND3X1_1 ( .A(_23_), .B(_25_), .C(_24_), .Y(_26_) );
INVX8 INVX8_1 ( .A(_20__bF_buf3), .Y(_27_) );
OAI21X1 OAI21X1_1 ( .A(_26__bF_buf3), .B(_27__bF_buf3), .C(loop_limit_inst_compare_inst_number0_0_), .Y(_28_) );
AOI21X1 AOI21X1_1 ( .A(_21_), .B(_28_), .C(_10__bF_buf3), .Y(_3__0_) );
NAND3X1 NAND3X1_2 ( .A(current_loop_actualize_1_), .B(_20__bF_buf2), .C(_18__bF_buf3), .Y(_29_) );
OAI21X1 OAI21X1_2 ( .A(_26__bF_buf2), .B(_27__bF_buf2), .C(loop_limit_inst_compare_inst_number0_1_), .Y(_30_) );
AOI21X1 AOI21X1_2 ( .A(_29_), .B(_30_), .C(_10__bF_buf2), .Y(_3__1_) );
NAND3X1 NAND3X1_3 ( .A(current_loop_actualize_2_), .B(_20__bF_buf1), .C(_18__bF_buf2), .Y(_31_) );
OAI21X1 OAI21X1_3 ( .A(_26__bF_buf1), .B(_27__bF_buf1), .C(loop_limit_inst_compare_inst_number0_2_), .Y(_32_) );
AOI21X1 AOI21X1_3 ( .A(_31_), .B(_32_), .C(_10__bF_buf1), .Y(_3__2_) );
NAND3X1 NAND3X1_4 ( .A(current_loop_actualize_3_), .B(_20__bF_buf0), .C(_18__bF_buf1), .Y(_33_) );
OAI21X1 OAI21X1_4 ( .A(_26__bF_buf0), .B(_27__bF_buf0), .C(loop_limit_inst_compare_inst_number0_3_), .Y(_34_) );
AOI21X1 AOI21X1_4 ( .A(_33_), .B(_34_), .C(_10__bF_buf0), .Y(_3__3_) );
NAND3X1 NAND3X1_5 ( .A(current_loop_actualize_4_), .B(_20__bF_buf3), .C(_18__bF_buf0), .Y(_35_) );
OAI21X1 OAI21X1_5 ( .A(_26__bF_buf3), .B(_27__bF_buf3), .C(loop_limit_inst_compare_inst_number0_4_), .Y(_36_) );
AOI21X1 AOI21X1_5 ( .A(_35_), .B(_36_), .C(_10__bF_buf3), .Y(_3__4_) );
NAND3X1 NAND3X1_6 ( .A(current_loop_actualize_5_), .B(_20__bF_buf2), .C(_18__bF_buf3), .Y(_37_) );
OAI21X1 OAI21X1_6 ( .A(_26__bF_buf2), .B(_27__bF_buf2), .C(loop_limit_inst_compare_inst_number0_5_), .Y(_38_) );
AOI21X1 AOI21X1_6 ( .A(_37_), .B(_38_), .C(_10__bF_buf2), .Y(_3__5_) );
NAND3X1 NAND3X1_7 ( .A(current_loop_actualize_6_), .B(_20__bF_buf1), .C(_18__bF_buf2), .Y(_39_) );
OAI21X1 OAI21X1_7 ( .A(_26__bF_buf1), .B(_27__bF_buf1), .C(loop_limit_inst_compare_inst_number0_6_), .Y(_40_) );
AOI21X1 AOI21X1_7 ( .A(_39_), .B(_40_), .C(_10__bF_buf1), .Y(_3__6_) );
NAND3X1 NAND3X1_8 ( .A(current_loop_actualize_7_), .B(_20__bF_buf0), .C(_18__bF_buf1), .Y(_41_) );
OAI21X1 OAI21X1_8 ( .A(_26__bF_buf0), .B(_27__bF_buf0), .C(loop_limit_inst_compare_inst_number0_7_), .Y(_42_) );
AOI21X1 AOI21X1_8 ( .A(_41_), .B(_42_), .C(_10__bF_buf0), .Y(_3__7_) );
NAND3X1 NAND3X1_9 ( .A(current_loop_actualize_8_), .B(_20__bF_buf3), .C(_18__bF_buf0), .Y(_43_) );
OAI21X1 OAI21X1_9 ( .A(_26__bF_buf3), .B(_27__bF_buf3), .C(loop_limit_inst_compare_inst_number0_8_), .Y(_44_) );
AOI21X1 AOI21X1_9 ( .A(_43_), .B(_44_), .C(_10__bF_buf3), .Y(_3__8_) );
NAND3X1 NAND3X1_10 ( .A(current_loop_actualize_9_), .B(_20__bF_buf2), .C(_18__bF_buf3), .Y(_45_) );
OAI21X1 OAI21X1_10 ( .A(_26__bF_buf2), .B(_27__bF_buf2), .C(loop_limit_inst_compare_inst_number0_9_), .Y(_46_) );
AOI21X1 AOI21X1_10 ( .A(_45_), .B(_46_), .C(_10__bF_buf2), .Y(_3__9_) );
NAND3X1 NAND3X1_11 ( .A(current_loop_actualize_10_), .B(_20__bF_buf1), .C(_18__bF_buf2), .Y(_47_) );
OAI21X1 OAI21X1_11 ( .A(_26__bF_buf1), .B(_27__bF_buf1), .C(loop_limit_inst_compare_inst_number0_10_), .Y(_48_) );
AOI21X1 AOI21X1_11 ( .A(_47_), .B(_48_), .C(_10__bF_buf1), .Y(_3__10_) );
NAND3X1 NAND3X1_12 ( .A(current_loop_actualize_11_), .B(_20__bF_buf0), .C(_18__bF_buf1), .Y(_49_) );
OAI21X1 OAI21X1_12 ( .A(_26__bF_buf0), .B(_27__bF_buf0), .C(loop_limit_inst_compare_inst_number0_11_), .Y(_50_) );
AOI21X1 AOI21X1_12 ( .A(_49_), .B(_50_), .C(_10__bF_buf0), .Y(_3__11_) );
NAND3X1 NAND3X1_13 ( .A(current_loop_actualize_12_), .B(_20__bF_buf3), .C(_18__bF_buf0), .Y(_51_) );
OAI21X1 OAI21X1_13 ( .A(_26__bF_buf3), .B(_27__bF_buf3), .C(loop_limit_inst_compare_inst_number0_12_), .Y(_52_) );
AOI21X1 AOI21X1_13 ( .A(_51_), .B(_52_), .C(_10__bF_buf3), .Y(_3__12_) );
NAND3X1 NAND3X1_14 ( .A(current_loop_actualize_13_), .B(_20__bF_buf2), .C(_18__bF_buf3), .Y(_53_) );
OAI21X1 OAI21X1_14 ( .A(_26__bF_buf2), .B(_27__bF_buf2), .C(loop_limit_inst_compare_inst_number0_13_), .Y(_54_) );
AOI21X1 AOI21X1_14 ( .A(_53_), .B(_54_), .C(_10__bF_buf2), .Y(_3__13_) );
NAND3X1 NAND3X1_15 ( .A(current_loop_actualize_14_), .B(_20__bF_buf1), .C(_18__bF_buf2), .Y(_55_) );
OAI21X1 OAI21X1_15 ( .A(_26__bF_buf1), .B(_27__bF_buf1), .C(loop_limit_inst_compare_inst_number0_14_), .Y(_56_) );
AOI21X1 AOI21X1_15 ( .A(_55_), .B(_56_), .C(_10__bF_buf1), .Y(_3__14_) );
NAND3X1 NAND3X1_16 ( .A(current_loop_actualize_15_), .B(_20__bF_buf0), .C(_18__bF_buf1), .Y(_57_) );
OAI21X1 OAI21X1_16 ( .A(_26__bF_buf0), .B(_27__bF_buf0), .C(loop_limit_inst_compare_inst_number0_15_), .Y(_58_) );
AOI21X1 AOI21X1_16 ( .A(_57_), .B(_58_), .C(_10__bF_buf0), .Y(_3__15_) );
INVX2 INVX2_1 ( .A(_135_), .Y(_59_) );
NAND2X1 NAND2X1_2 ( .A(reset_bF_buf5), .B(validity_validity_reg), .Y(_60_) );
NOR2X1 NOR2X1_2 ( .A(start), .B(_10__bF_buf3), .Y(_61_) );
AOI21X1 AOI21X1_17 ( .A(_59_), .B(_60_), .C(_61_), .Y(_1_) );
INVX1 INVX1_1 ( .A(_139__0_), .Y(_62_) );
OAI21X1 OAI21X1_17 ( .A(_10__bF_buf2), .B(start), .C(_60_), .Y(_63_) );
OAI21X1 OAI21X1_18 ( .A(_10__bF_buf1), .B(start), .C(hash_array2_2), .Y(_64_) );
AOI22X1 AOI22X1_1 ( .A(_62_), .B(_60_), .C(_63__bF_buf3), .D(_64_), .Y(_7__0_) );
INVX1 INVX1_2 ( .A(_139__1_), .Y(_65_) );
NOR2X1 NOR2X1_3 ( .A(_65_), .B(_63__bF_buf2), .Y(_7__1_) );
INVX1 INVX1_3 ( .A(_139__2_), .Y(_66_) );
NOR2X1 NOR2X1_4 ( .A(_66_), .B(_63__bF_buf1), .Y(_7__2_) );
INVX1 INVX1_4 ( .A(_139__3_), .Y(_67_) );
NOR2X1 NOR2X1_5 ( .A(_67_), .B(_63__bF_buf0), .Y(_7__3_) );
INVX1 INVX1_5 ( .A(_139__4_), .Y(_68_) );
NOR2X1 NOR2X1_6 ( .A(_68_), .B(_63__bF_buf3), .Y(_7__4_) );
INVX1 INVX1_6 ( .A(_139__5_), .Y(_69_) );
NOR2X1 NOR2X1_7 ( .A(_69_), .B(_63__bF_buf2), .Y(_7__5_) );
INVX1 INVX1_7 ( .A(_139__6_), .Y(_70_) );
NOR2X1 NOR2X1_8 ( .A(_70_), .B(_63__bF_buf1), .Y(_7__6_) );
INVX1 INVX1_8 ( .A(_139__7_), .Y(_71_) );
NOR2X1 NOR2X1_9 ( .A(_71_), .B(_63__bF_buf0), .Y(_7__7_) );
INVX1 INVX1_9 ( .A(_138__0_), .Y(_72_) );
OAI21X1 OAI21X1_19 ( .A(_10__bF_buf0), .B(start), .C(hash_array2_1), .Y(_73_) );
AOI22X1 AOI22X1_2 ( .A(_72_), .B(_60_), .C(_63__bF_buf3), .D(_73_), .Y(_6__0_) );
INVX1 INVX1_10 ( .A(_138__1_), .Y(_74_) );
NOR2X1 NOR2X1_10 ( .A(_74_), .B(_63__bF_buf2), .Y(_6__1_) );
INVX1 INVX1_11 ( .A(_138__2_), .Y(_75_) );
NOR2X1 NOR2X1_11 ( .A(_75_), .B(_63__bF_buf1), .Y(_6__2_) );
INVX1 INVX1_12 ( .A(_138__3_), .Y(_76_) );
NOR2X1 NOR2X1_12 ( .A(_76_), .B(_63__bF_buf0), .Y(_6__3_) );
INVX1 INVX1_13 ( .A(_138__4_), .Y(_77_) );
NOR2X1 NOR2X1_13 ( .A(_77_), .B(_63__bF_buf3), .Y(_6__4_) );
INVX1 INVX1_14 ( .A(_138__5_), .Y(_78_) );
NOR2X1 NOR2X1_14 ( .A(_78_), .B(_63__bF_buf2), .Y(_6__5_) );
INVX1 INVX1_15 ( .A(_138__6_), .Y(_79_) );
NOR2X1 NOR2X1_15 ( .A(_79_), .B(_63__bF_buf1), .Y(_6__6_) );
INVX1 INVX1_16 ( .A(_138__7_), .Y(_80_) );
NOR2X1 NOR2X1_16 ( .A(_80_), .B(_63__bF_buf0), .Y(_6__7_) );
INVX1 INVX1_17 ( .A(_137__0_), .Y(_81_) );
INVX1 INVX1_18 ( .A(validity_validity_reg), .Y(_82_) );
OAI21X1 OAI21X1_20 ( .A(_82_), .B(hash_array2_0), .C(start), .Y(_83_) );
AOI22X1 AOI22X1_3 ( .A(_81_), .B(_60_), .C(_83_), .D(reset_bF_buf4), .Y(_5__0_) );
INVX1 INVX1_19 ( .A(_137__1_), .Y(_84_) );
NOR2X1 NOR2X1_17 ( .A(_84_), .B(_63__bF_buf3), .Y(_5__1_) );
INVX1 INVX1_20 ( .A(_137__2_), .Y(_85_) );
NOR2X1 NOR2X1_18 ( .A(_85_), .B(_63__bF_buf2), .Y(_5__2_) );
INVX1 INVX1_21 ( .A(_137__3_), .Y(_86_) );
NOR2X1 NOR2X1_19 ( .A(_86_), .B(_63__bF_buf1), .Y(_5__3_) );
INVX1 INVX1_22 ( .A(_137__4_), .Y(_87_) );
NOR2X1 NOR2X1_20 ( .A(_87_), .B(_63__bF_buf0), .Y(_5__4_) );
INVX1 INVX1_23 ( .A(_137__5_), .Y(_88_) );
NOR2X1 NOR2X1_21 ( .A(_88_), .B(_63__bF_buf3), .Y(_5__5_) );
INVX1 INVX1_24 ( .A(_137__6_), .Y(_89_) );
NOR2X1 NOR2X1_22 ( .A(_89_), .B(_63__bF_buf2), .Y(_5__6_) );
INVX1 INVX1_25 ( .A(_137__7_), .Y(_90_) );
NOR2X1 NOR2X1_23 ( .A(_90_), .B(_63__bF_buf1), .Y(_5__7_) );
INVX1 INVX1_26 ( .A(_136__0_), .Y(_91_) );
OR2X2 OR2X2_1 ( .A(_61_), .B(hash_array2_0), .Y(_92_) );
AOI22X1 AOI22X1_4 ( .A(_91_), .B(_60_), .C(_92_), .D(_63__bF_buf0), .Y(_4__0_) );
INVX1 INVX1_27 ( .A(_136__1_), .Y(_93_) );
AOI21X1 AOI21X1_18 ( .A(_93_), .B(_60_), .C(_61_), .Y(_4__1_) );
INVX1 INVX1_28 ( .A(_136__2_), .Y(_94_) );
AOI21X1 AOI21X1_19 ( .A(_94_), .B(_60_), .C(_61_), .Y(_4__2_) );
INVX1 INVX1_29 ( .A(_136__3_), .Y(_95_) );
AOI21X1 AOI21X1_20 ( .A(_95_), .B(_60_), .C(_61_), .Y(_4__3_) );
INVX1 INVX1_30 ( .A(_136__4_), .Y(_96_) );
AOI21X1 AOI21X1_21 ( .A(_96_), .B(_60_), .C(_61_), .Y(_4__4_) );
INVX1 INVX1_31 ( .A(_136__5_), .Y(_97_) );
AOI21X1 AOI21X1_22 ( .A(_97_), .B(_60_), .C(_61_), .Y(_4__5_) );
INVX1 INVX1_32 ( .A(_136__6_), .Y(_98_) );
AOI21X1 AOI21X1_23 ( .A(_98_), .B(_60_), .C(_61_), .Y(_4__6_) );
INVX1 INVX1_33 ( .A(_136__7_), .Y(_99_) );
AOI21X1 AOI21X1_24 ( .A(_99_), .B(_60_), .C(_61_), .Y(_4__7_) );
NAND2X1 NAND2X1_3 ( .A(start), .B(counter_0_), .Y(_100_) );
INVX1 INVX1_34 ( .A(_100_), .Y(_101_) );
OAI21X1 OAI21X1_21 ( .A(start), .B(counter_0_), .C(reset_bF_buf3), .Y(_102_) );
NOR2X1 NOR2X1_24 ( .A(_102_), .B(_101_), .Y(_0__0_) );
NOR2X1 NOR2X1_25 ( .A(_27__bF_buf3), .B(_26__bF_buf3), .Y(_103_) );
NAND2X1 NAND2X1_4 ( .A(_11_), .B(_100_), .Y(_104_) );
NAND2X1 NAND2X1_5 ( .A(counter_1_), .B(_101_), .Y(_105_) );
NAND3X1 NAND3X1_17 ( .A(reset_bF_buf2), .B(_104_), .C(_105_), .Y(_106_) );
NOR2X1 NOR2X1_26 ( .A(_106_), .B(_103_), .Y(_0__1_) );
NAND2X1 NAND2X1_6 ( .A(counter_2_), .B(counter_1_), .Y(_107_) );
NOR2X1 NOR2X1_27 ( .A(_100_), .B(_107_), .Y(_108_) );
INVX1 INVX1_35 ( .A(_105_), .Y(_109_) );
OAI21X1 OAI21X1_22 ( .A(_109_), .B(counter_2_), .C(reset_bF_buf1), .Y(_110_) );
NOR2X1 NOR2X1_28 ( .A(_108_), .B(_110_), .Y(_0__2_) );
AND2X2 AND2X2_3 ( .A(_108_), .B(counter_3_), .Y(_111_) );
OAI21X1 OAI21X1_23 ( .A(_108_), .B(counter_3_), .C(reset_bF_buf0), .Y(_112_) );
OR2X2 OR2X2_2 ( .A(_111_), .B(_112_), .Y(_113_) );
NOR2X1 NOR2X1_29 ( .A(_103_), .B(_113_), .Y(_0__3_) );
OAI21X1 OAI21X1_24 ( .A(_111_), .B(counter_4_), .C(reset_bF_buf5), .Y(_114_) );
AOI21X1 AOI21X1_25 ( .A(counter_4_), .B(_111_), .C(_114_), .Y(_0__4_) );
AOI21X1 AOI21X1_26 ( .A(counter_4_), .B(_111_), .C(counter_5_), .Y(_115_) );
NAND2X1 NAND2X1_7 ( .A(counter_3_), .B(_108_), .Y(_116_) );
NAND2X1 NAND2X1_8 ( .A(counter_5_), .B(counter_4_), .Y(_117_) );
OAI21X1 OAI21X1_25 ( .A(_116_), .B(_117_), .C(reset_bF_buf4), .Y(_118_) );
NOR2X1 NOR2X1_30 ( .A(_118_), .B(_115_), .Y(_0__5_) );
INVX1 INVX1_36 ( .A(_117_), .Y(_119_) );
AOI21X1 AOI21X1_27 ( .A(_119_), .B(_111_), .C(counter_6_), .Y(_120_) );
NAND2X1 NAND2X1_9 ( .A(counter_6_), .B(_119_), .Y(_121_) );
OAI21X1 OAI21X1_26 ( .A(_116_), .B(_121_), .C(reset_bF_buf3), .Y(_122_) );
NOR2X1 NOR2X1_31 ( .A(_122_), .B(_120_), .Y(_0__6_) );
OAI21X1 OAI21X1_27 ( .A(_116_), .B(_121_), .C(counter_7_), .Y(_123_) );
INVX1 INVX1_37 ( .A(counter_7_), .Y(_124_) );
INVX1 INVX1_38 ( .A(_121_), .Y(_125_) );
NAND3X1 NAND3X1_18 ( .A(_124_), .B(_111_), .C(_125_), .Y(_126_) );
AOI21X1 AOI21X1_28 ( .A(_123_), .B(_126_), .C(_10__bF_buf3), .Y(_0__7_) );
NOR2X1 NOR2X1_32 ( .A(_19_), .B(_82_), .Y(_127_) );
OAI21X1 OAI21X1_28 ( .A(start), .B(invalid_nonce), .C(reset_bF_buf2), .Y(_128_) );
NOR2X1 NOR2X1_33 ( .A(_128_), .B(_127_), .Y(_2_) );
INVX1 INVX1_39 ( .A(micro_counter_inst_ready), .Y(_129_) );
OAI21X1 OAI21X1_29 ( .A(_59_), .B(_129_), .C(_127_), .Y(_130_) );
AOI21X1 AOI21X1_29 ( .A(_59_), .B(_129_), .C(_130_), .Y(_131_) );
OAI21X1 OAI21X1_30 ( .A(start), .B(micro_counter_inst_ready), .C(reset_bF_buf1), .Y(_132_) );
AOI21X1 AOI21X1_30 ( .A(_18__bF_buf0), .B(_131_), .C(_132_), .Y(_8_) );
INVX1 INVX1_40 ( .A(fail), .Y(_133_) );
OAI21X1 OAI21X1_31 ( .A(start), .B(loop_limit_inst_stop), .C(reset_bF_buf0), .Y(_134_) );
AOI21X1 AOI21X1_31 ( .A(_133_), .B(_20__bF_buf3), .C(_134_), .Y(_9_) );
BUFX2 BUFX2_1 ( .A(_135_), .Y(finish) );
BUFX2 BUFX2_2 ( .A(_136__0_), .Y(nonce0[0]) );
BUFX2 BUFX2_3 ( .A(_136__1_), .Y(nonce0[1]) );
BUFX2 BUFX2_4 ( .A(_136__2_), .Y(nonce0[2]) );
BUFX2 BUFX2_5 ( .A(_136__3_), .Y(nonce0[3]) );
BUFX2 BUFX2_6 ( .A(_136__4_), .Y(nonce0[4]) );
BUFX2 BUFX2_7 ( .A(_136__5_), .Y(nonce0[5]) );
BUFX2 BUFX2_8 ( .A(_136__6_), .Y(nonce0[6]) );
BUFX2 BUFX2_9 ( .A(_136__7_), .Y(nonce0[7]) );
BUFX2 BUFX2_10 ( .A(_137__0_), .Y(nonce1[0]) );
BUFX2 BUFX2_11 ( .A(_137__1_), .Y(nonce1[1]) );
BUFX2 BUFX2_12 ( .A(_137__2_), .Y(nonce1[2]) );
BUFX2 BUFX2_13 ( .A(_137__3_), .Y(nonce1[3]) );
BUFX2 BUFX2_14 ( .A(_137__4_), .Y(nonce1[4]) );
BUFX2 BUFX2_15 ( .A(_137__5_), .Y(nonce1[5]) );
BUFX2 BUFX2_16 ( .A(_137__6_), .Y(nonce1[6]) );
BUFX2 BUFX2_17 ( .A(_137__7_), .Y(nonce1[7]) );
BUFX2 BUFX2_18 ( .A(_138__0_), .Y(nonce2[0]) );
BUFX2 BUFX2_19 ( .A(_138__1_), .Y(nonce2[1]) );
BUFX2 BUFX2_20 ( .A(_138__2_), .Y(nonce2[2]) );
BUFX2 BUFX2_21 ( .A(_138__3_), .Y(nonce2[3]) );
BUFX2 BUFX2_22 ( .A(_138__4_), .Y(nonce2[4]) );
BUFX2 BUFX2_23 ( .A(_138__5_), .Y(nonce2[5]) );
BUFX2 BUFX2_24 ( .A(_138__6_), .Y(nonce2[6]) );
BUFX2 BUFX2_25 ( .A(_138__7_), .Y(nonce2[7]) );
BUFX2 BUFX2_26 ( .A(_139__0_), .Y(nonce3[0]) );
BUFX2 BUFX2_27 ( .A(_139__1_), .Y(nonce3[1]) );
BUFX2 BUFX2_28 ( .A(_139__2_), .Y(nonce3[2]) );
BUFX2 BUFX2_29 ( .A(_139__3_), .Y(nonce3[3]) );
BUFX2 BUFX2_30 ( .A(_139__4_), .Y(nonce3[4]) );
BUFX2 BUFX2_31 ( .A(_139__5_), .Y(nonce3[5]) );
BUFX2 BUFX2_32 ( .A(_139__6_), .Y(nonce3[6]) );
BUFX2 BUFX2_33 ( .A(_139__7_), .Y(nonce3[7]) );
DFFPOSX1 DFFPOSX1_1 ( .CLK(clk_bF_buf11), .D(_9_), .Q(loop_limit_inst_stop) );
DFFPOSX1 DFFPOSX1_2 ( .CLK(clk_bF_buf10), .D(_8_), .Q(micro_counter_inst_ready) );
DFFPOSX1 DFFPOSX1_3 ( .CLK(clk_bF_buf9), .D(_0__0_), .Q(counter_0_) );
DFFPOSX1 DFFPOSX1_4 ( .CLK(clk_bF_buf8), .D(_0__1_), .Q(counter_1_) );
DFFPOSX1 DFFPOSX1_5 ( .CLK(clk_bF_buf7), .D(_0__2_), .Q(counter_2_) );
DFFPOSX1 DFFPOSX1_6 ( .CLK(clk_bF_buf6), .D(_0__3_), .Q(counter_3_) );
DFFPOSX1 DFFPOSX1_7 ( .CLK(clk_bF_buf5), .D(_0__4_), .Q(counter_4_) );
DFFPOSX1 DFFPOSX1_8 ( .CLK(clk_bF_buf4), .D(_0__5_), .Q(counter_5_) );
DFFPOSX1 DFFPOSX1_9 ( .CLK(clk_bF_buf3), .D(_0__6_), .Q(counter_6_) );
DFFPOSX1 DFFPOSX1_10 ( .CLK(clk_bF_buf2), .D(_0__7_), .Q(counter_7_) );
DFFPOSX1 DFFPOSX1_11 ( .CLK(clk_bF_buf1), .D(_4__0_), .Q(_136__0_) );
DFFPOSX1 DFFPOSX1_12 ( .CLK(clk_bF_buf0), .D(_4__1_), .Q(_136__1_) );
DFFPOSX1 DFFPOSX1_13 ( .CLK(clk_bF_buf11), .D(_4__2_), .Q(_136__2_) );
DFFPOSX1 DFFPOSX1_14 ( .CLK(clk_bF_buf10), .D(_4__3_), .Q(_136__3_) );
DFFPOSX1 DFFPOSX1_15 ( .CLK(clk_bF_buf9), .D(_4__4_), .Q(_136__4_) );
DFFPOSX1 DFFPOSX1_16 ( .CLK(clk_bF_buf8), .D(_4__5_), .Q(_136__5_) );
DFFPOSX1 DFFPOSX1_17 ( .CLK(clk_bF_buf7), .D(_4__6_), .Q(_136__6_) );
DFFPOSX1 DFFPOSX1_18 ( .CLK(clk_bF_buf6), .D(_4__7_), .Q(_136__7_) );
DFFPOSX1 DFFPOSX1_19 ( .CLK(clk_bF_buf5), .D(_5__0_), .Q(_137__0_) );
DFFPOSX1 DFFPOSX1_20 ( .CLK(clk_bF_buf4), .D(_5__1_), .Q(_137__1_) );
DFFPOSX1 DFFPOSX1_21 ( .CLK(clk_bF_buf3), .D(_5__2_), .Q(_137__2_) );
DFFPOSX1 DFFPOSX1_22 ( .CLK(clk_bF_buf2), .D(_5__3_), .Q(_137__3_) );
DFFPOSX1 DFFPOSX1_23 ( .CLK(clk_bF_buf1), .D(_5__4_), .Q(_137__4_) );
DFFPOSX1 DFFPOSX1_24 ( .CLK(clk_bF_buf0), .D(_5__5_), .Q(_137__5_) );
DFFPOSX1 DFFPOSX1_25 ( .CLK(clk_bF_buf11), .D(_5__6_), .Q(_137__6_) );
DFFPOSX1 DFFPOSX1_26 ( .CLK(clk_bF_buf10), .D(_5__7_), .Q(_137__7_) );
DFFPOSX1 DFFPOSX1_27 ( .CLK(clk_bF_buf9), .D(_6__0_), .Q(_138__0_) );
DFFPOSX1 DFFPOSX1_28 ( .CLK(clk_bF_buf8), .D(_6__1_), .Q(_138__1_) );
DFFPOSX1 DFFPOSX1_29 ( .CLK(clk_bF_buf7), .D(_6__2_), .Q(_138__2_) );
DFFPOSX1 DFFPOSX1_30 ( .CLK(clk_bF_buf6), .D(_6__3_), .Q(_138__3_) );
DFFPOSX1 DFFPOSX1_31 ( .CLK(clk_bF_buf5), .D(_6__4_), .Q(_138__4_) );
DFFPOSX1 DFFPOSX1_32 ( .CLK(clk_bF_buf4), .D(_6__5_), .Q(_138__5_) );
DFFPOSX1 DFFPOSX1_33 ( .CLK(clk_bF_buf3), .D(_6__6_), .Q(_138__6_) );
DFFPOSX1 DFFPOSX1_34 ( .CLK(clk_bF_buf2), .D(_6__7_), .Q(_138__7_) );
DFFPOSX1 DFFPOSX1_35 ( .CLK(clk_bF_buf1), .D(_7__0_), .Q(_139__0_) );
DFFPOSX1 DFFPOSX1_36 ( .CLK(clk_bF_buf0), .D(_7__1_), .Q(_139__1_) );
DFFPOSX1 DFFPOSX1_37 ( .CLK(clk_bF_buf11), .D(_7__2_), .Q(_139__2_) );
DFFPOSX1 DFFPOSX1_38 ( .CLK(clk_bF_buf10), .D(_7__3_), .Q(_139__3_) );
DFFPOSX1 DFFPOSX1_39 ( .CLK(clk_bF_buf9), .D(_7__4_), .Q(_139__4_) );
DFFPOSX1 DFFPOSX1_40 ( .CLK(clk_bF_buf8), .D(_7__5_), .Q(_139__5_) );
DFFPOSX1 DFFPOSX1_41 ( .CLK(clk_bF_buf7), .D(_7__6_), .Q(_139__6_) );
DFFPOSX1 DFFPOSX1_42 ( .CLK(clk_bF_buf6), .D(_7__7_), .Q(_139__7_) );
DFFPOSX1 DFFPOSX1_43 ( .CLK(clk_bF_buf5), .D(_1_), .Q(_135_) );
DFFPOSX1 DFFPOSX1_44 ( .CLK(clk_bF_buf4), .D(_3__0_), .Q(loop_limit_inst_compare_inst_number0_0_) );
DFFPOSX1 DFFPOSX1_45 ( .CLK(clk_bF_buf3), .D(_3__1_), .Q(loop_limit_inst_compare_inst_number0_1_) );
DFFPOSX1 DFFPOSX1_46 ( .CLK(clk_bF_buf2), .D(_3__2_), .Q(loop_limit_inst_compare_inst_number0_2_) );
DFFPOSX1 DFFPOSX1_47 ( .CLK(clk_bF_buf1), .D(_3__3_), .Q(loop_limit_inst_compare_inst_number0_3_) );
DFFPOSX1 DFFPOSX1_48 ( .CLK(clk_bF_buf0), .D(_3__4_), .Q(loop_limit_inst_compare_inst_number0_4_) );
DFFPOSX1 DFFPOSX1_49 ( .CLK(clk_bF_buf11), .D(_3__5_), .Q(loop_limit_inst_compare_inst_number0_5_) );
DFFPOSX1 DFFPOSX1_50 ( .CLK(clk_bF_buf10), .D(_3__6_), .Q(loop_limit_inst_compare_inst_number0_6_) );
DFFPOSX1 DFFPOSX1_51 ( .CLK(clk_bF_buf9), .D(_3__7_), .Q(loop_limit_inst_compare_inst_number0_7_) );
DFFPOSX1 DFFPOSX1_52 ( .CLK(clk_bF_buf8), .D(_3__8_), .Q(loop_limit_inst_compare_inst_number0_8_) );
DFFPOSX1 DFFPOSX1_53 ( .CLK(clk_bF_buf7), .D(_3__9_), .Q(loop_limit_inst_compare_inst_number0_9_) );
DFFPOSX1 DFFPOSX1_54 ( .CLK(clk_bF_buf6), .D(_3__10_), .Q(loop_limit_inst_compare_inst_number0_10_) );
DFFPOSX1 DFFPOSX1_55 ( .CLK(clk_bF_buf5), .D(_3__11_), .Q(loop_limit_inst_compare_inst_number0_11_) );
DFFPOSX1 DFFPOSX1_56 ( .CLK(clk_bF_buf4), .D(_3__12_), .Q(loop_limit_inst_compare_inst_number0_12_) );
DFFPOSX1 DFFPOSX1_57 ( .CLK(clk_bF_buf3), .D(_3__13_), .Q(loop_limit_inst_compare_inst_number0_13_) );
DFFPOSX1 DFFPOSX1_58 ( .CLK(clk_bF_buf2), .D(_3__14_), .Q(loop_limit_inst_compare_inst_number0_14_) );
DFFPOSX1 DFFPOSX1_59 ( .CLK(clk_bF_buf1), .D(_3__15_), .Q(loop_limit_inst_compare_inst_number0_15_) );
DFFPOSX1 DFFPOSX1_60 ( .CLK(clk_bF_buf0), .D(_2_), .Q(invalid_nonce) );
INVX1 INVX1_41 ( .A(gnd), .Y(_194_) );
NAND2X1 NAND2X1_10 ( .A(target[15]), .B(_194_), .Y(_195_) );
INVX1 INVX1_42 ( .A(gnd), .Y(_196_) );
NAND2X1 NAND2X1_11 ( .A(target[14]), .B(_196_), .Y(_197_) );
INVX2 INVX2_2 ( .A(target[15]), .Y(_198_) );
INVX1 INVX1_43 ( .A(target[14]), .Y(_199_) );
AOI22X1 AOI22X1_5 ( .A(_198_), .B(gnd), .C(_199_), .D(gnd), .Y(_200_) );
NAND3X1 NAND3X1_19 ( .A(_195_), .B(_197_), .C(_200_), .Y(_201_) );
INVX1 INVX1_44 ( .A(gnd), .Y(_202_) );
INVX1 INVX1_45 ( .A(gnd), .Y(_203_) );
AOI22X1 AOI22X1_6 ( .A(_202_), .B(target[13]), .C(target[12]), .D(_203_), .Y(_204_) );
INVX1 INVX1_46 ( .A(target[13]), .Y(_205_) );
NAND2X1 NAND2X1_12 ( .A(gnd), .B(_205_), .Y(_206_) );
INVX1 INVX1_47 ( .A(target[12]), .Y(_207_) );
NAND2X1 NAND2X1_13 ( .A(gnd), .B(_207_), .Y(_208_) );
NAND3X1 NAND3X1_20 ( .A(_206_), .B(_208_), .C(_204_), .Y(_209_) );
NOR2X1 NOR2X1_34 ( .A(_201_), .B(_209_), .Y(_210_) );
XNOR2X1 XNOR2X1_1 ( .A(gnd), .B(target[11]), .Y(_211_) );
INVX2 INVX2_3 ( .A(target[10]), .Y(_212_) );
OR2X2 OR2X2_3 ( .A(_212_), .B(gnd), .Y(_213_) );
NAND2X1 NAND2X1_14 ( .A(gnd), .B(_212_), .Y(_214_) );
NAND3X1 NAND3X1_21 ( .A(_213_), .B(_214_), .C(_211_), .Y(_215_) );
INVX1 INVX1_48 ( .A(gnd), .Y(_216_) );
INVX1 INVX1_49 ( .A(gnd), .Y(_217_) );
AOI22X1 AOI22X1_7 ( .A(_216_), .B(target[9]), .C(target[8]), .D(_217_), .Y(_218_) );
INVX1 INVX1_50 ( .A(target[9]), .Y(_219_) );
NAND2X1 NAND2X1_15 ( .A(gnd), .B(_219_), .Y(_220_) );
INVX1 INVX1_51 ( .A(target[8]), .Y(_221_) );
NAND2X1 NAND2X1_16 ( .A(gnd), .B(_221_), .Y(_222_) );
NAND3X1 NAND3X1_22 ( .A(_220_), .B(_222_), .C(_218_), .Y(_223_) );
NOR2X1 NOR2X1_35 ( .A(_223_), .B(_215_), .Y(_224_) );
AND2X2 AND2X2_4 ( .A(_224_), .B(_210_), .Y(_225_) );
XOR2X1 XOR2X1_1 ( .A(gnd), .B(target[7]), .Y(_226_) );
XOR2X1 XOR2X1_2 ( .A(target[6]), .B(gnd), .Y(_227_) );
NOR2X1 NOR2X1_36 ( .A(_226_), .B(_227_), .Y(_228_) );
INVX1 INVX1_52 ( .A(gnd), .Y(_229_) );
INVX1 INVX1_53 ( .A(gnd), .Y(_230_) );
AOI22X1 AOI22X1_8 ( .A(_229_), .B(target[5]), .C(target[4]), .D(_230_), .Y(_231_) );
INVX1 INVX1_54 ( .A(target[5]), .Y(_232_) );
INVX1 INVX1_55 ( .A(target[4]), .Y(_233_) );
AOI22X1 AOI22X1_9 ( .A(_232_), .B(gnd), .C(_233_), .D(gnd), .Y(_234_) );
AND2X2 AND2X2_5 ( .A(_231_), .B(_234_), .Y(_235_) );
NAND2X1 NAND2X1_17 ( .A(_228_), .B(_235_), .Y(_236_) );
NOR2X1 NOR2X1_37 ( .A(target[3]), .B(gnd), .Y(_237_) );
INVX1 INVX1_56 ( .A(_237_), .Y(_238_) );
NAND2X1 NAND2X1_18 ( .A(target[3]), .B(gnd), .Y(_239_) );
XOR2X1 XOR2X1_3 ( .A(target[2]), .B(gnd), .Y(_240_) );
AOI21X1 AOI21X1_32 ( .A(_238_), .B(_239_), .C(_240_), .Y(_241_) );
INVX1 INVX1_57 ( .A(gnd), .Y(_242_) );
NAND2X1 NAND2X1_19 ( .A(target[1]), .B(_242_), .Y(_243_) );
NOR2X1 NOR2X1_38 ( .A(target[1]), .B(_242_), .Y(_244_) );
INVX1 INVX1_58 ( .A(hash_array2_0), .Y(_245_) );
NOR2X1 NOR2X1_39 ( .A(target[0]), .B(_245_), .Y(_246_) );
OAI21X1 OAI21X1_32 ( .A(_244_), .B(_246_), .C(_243_), .Y(_247_) );
NAND2X1 NAND2X1_20 ( .A(_247_), .B(_241_), .Y(_248_) );
INVX1 INVX1_59 ( .A(target[3]), .Y(_249_) );
NOR2X1 NOR2X1_40 ( .A(gnd), .B(_249_), .Y(_250_) );
NAND2X1 NAND2X1_21 ( .A(gnd), .B(_249_), .Y(_251_) );
INVX1 INVX1_60 ( .A(target[2]), .Y(_252_) );
NOR2X1 NOR2X1_41 ( .A(gnd), .B(_252_), .Y(_253_) );
AOI21X1 AOI21X1_33 ( .A(_251_), .B(_253_), .C(_250_), .Y(_141_) );
AOI21X1 AOI21X1_34 ( .A(_141_), .B(_248_), .C(_236_), .Y(_142_) );
XNOR2X1 XNOR2X1_2 ( .A(gnd), .B(target[7]), .Y(_143_) );
XNOR2X1 XNOR2X1_3 ( .A(target[6]), .B(gnd), .Y(_144_) );
NAND2X1 NAND2X1_22 ( .A(_143_), .B(_144_), .Y(_145_) );
OAI22X1 OAI22X1_1 ( .A(_232_), .B(gnd), .C(_233_), .D(gnd), .Y(_146_) );
OAI21X1 OAI21X1_33 ( .A(_229_), .B(target[5]), .C(_146_), .Y(_147_) );
INVX1 INVX1_61 ( .A(target[7]), .Y(_148_) );
NOR2X1 NOR2X1_42 ( .A(gnd), .B(_148_), .Y(_149_) );
INVX1 INVX1_62 ( .A(target[6]), .Y(_150_) );
NOR2X1 NOR2X1_43 ( .A(gnd), .B(_150_), .Y(_151_) );
AOI21X1 AOI21X1_35 ( .A(_151_), .B(_143_), .C(_149_), .Y(_152_) );
OAI21X1 OAI21X1_34 ( .A(_145_), .B(_147_), .C(_152_), .Y(_153_) );
OAI21X1 OAI21X1_35 ( .A(_142_), .B(_153_), .C(_225_), .Y(_154_) );
INVX1 INVX1_63 ( .A(target[11]), .Y(_155_) );
NOR2X1 NOR2X1_44 ( .A(gnd), .B(_155_), .Y(_156_) );
NOR2X1 NOR2X1_45 ( .A(gnd), .B(_212_), .Y(_157_) );
AOI21X1 AOI21X1_36 ( .A(_157_), .B(_211_), .C(_156_), .Y(_158_) );
OAI22X1 OAI22X1_2 ( .A(_219_), .B(gnd), .C(_221_), .D(gnd), .Y(_159_) );
OAI21X1 OAI21X1_36 ( .A(_216_), .B(target[9]), .C(_159_), .Y(_160_) );
OAI21X1 OAI21X1_37 ( .A(_215_), .B(_160_), .C(_158_), .Y(_161_) );
NOR2X1 NOR2X1_46 ( .A(target[13]), .B(_202_), .Y(_162_) );
OR2X2 OR2X2_4 ( .A(_204_), .B(_162_), .Y(_163_) );
AOI21X1 AOI21X1_37 ( .A(_198_), .B(gnd), .C(_197_), .Y(_164_) );
OAI21X1 OAI21X1_38 ( .A(_198_), .B(gnd), .C(reset_bF_buf5), .Y(_165_) );
NOR2X1 NOR2X1_47 ( .A(_165_), .B(_164_), .Y(_166_) );
OAI21X1 OAI21X1_39 ( .A(_201_), .B(_163_), .C(_166_), .Y(_167_) );
AOI21X1 AOI21X1_38 ( .A(_210_), .B(_161_), .C(_167_), .Y(_168_) );
INVX1 INVX1_64 ( .A(reset_bF_buf4), .Y(_169_) );
NAND2X1 NAND2X1_23 ( .A(compare_hash_0_compare_var_0_), .B(_169_), .Y(_170_) );
NAND2X1 NAND2X1_24 ( .A(_210_), .B(_224_), .Y(_171_) );
NAND2X1 NAND2X1_25 ( .A(_231_), .B(_234_), .Y(_172_) );
NOR2X1 NOR2X1_48 ( .A(_172_), .B(_145_), .Y(_173_) );
INVX1 INVX1_65 ( .A(_239_), .Y(_174_) );
XNOR2X1 XNOR2X1_4 ( .A(target[2]), .B(gnd), .Y(_175_) );
OAI21X1 OAI21X1_40 ( .A(_237_), .B(_174_), .C(_175_), .Y(_176_) );
XNOR2X1 XNOR2X1_5 ( .A(target[1]), .B(gnd), .Y(_177_) );
XNOR2X1 XNOR2X1_6 ( .A(target[0]), .B(hash_array2_0), .Y(_178_) );
NAND2X1 NAND2X1_26 ( .A(_177_), .B(_178_), .Y(_179_) );
NOR2X1 NOR2X1_49 ( .A(_179_), .B(_176_), .Y(_180_) );
NAND2X1 NAND2X1_27 ( .A(_173_), .B(_180_), .Y(_181_) );
OAI21X1 OAI21X1_41 ( .A(_171_), .B(_181_), .C(reset_bF_buf3), .Y(_182_) );
AOI22X1 AOI22X1_10 ( .A(_170_), .B(_182_), .C(_154_), .D(_168_), .Y(_140__0_) );
OR2X2 OR2X2_5 ( .A(reset_bF_buf2), .B(compare_hash_0_compare_var_1_), .Y(_183_) );
AND2X2 AND2X2_6 ( .A(_182_), .B(_183_), .Y(_140__1_) );
INVX1 INVX1_66 ( .A(compare_hash_0_compare_var_2_), .Y(_184_) );
INVX1 INVX1_67 ( .A(target[1]), .Y(_185_) );
NOR2X1 NOR2X1_50 ( .A(gnd), .B(_185_), .Y(_186_) );
NAND2X1 NAND2X1_28 ( .A(gnd), .B(_185_), .Y(_187_) );
INVX1 INVX1_68 ( .A(target[0]), .Y(_188_) );
NAND2X1 NAND2X1_29 ( .A(hash_array2_0), .B(_188_), .Y(_189_) );
AOI21X1 AOI21X1_39 ( .A(_187_), .B(_189_), .C(_186_), .Y(_190_) );
OAI21X1 OAI21X1_42 ( .A(_176_), .B(_190_), .C(_141_), .Y(_191_) );
AOI21X1 AOI21X1_40 ( .A(_173_), .B(_191_), .C(_153_), .Y(_192_) );
OAI21X1 OAI21X1_43 ( .A(_192_), .B(_171_), .C(_168_), .Y(_193_) );
OAI21X1 OAI21X1_44 ( .A(reset_bF_buf1), .B(_184_), .C(_193_), .Y(_140__2_) );
DFFPOSX1 DFFPOSX1_61 ( .CLK(clk_bF_buf11), .D(_140__0_), .Q(compare_hash_0_compare_var_0_) );
DFFPOSX1 DFFPOSX1_62 ( .CLK(clk_bF_buf10), .D(_140__1_), .Q(compare_hash_0_compare_var_1_) );
DFFPOSX1 DFFPOSX1_63 ( .CLK(clk_bF_buf9), .D(_140__2_), .Q(compare_hash_0_compare_var_2_) );
INVX1 INVX1_69 ( .A(gnd), .Y(_308_) );
NAND2X1 NAND2X1_30 ( .A(target[15]), .B(_308_), .Y(_309_) );
INVX1 INVX1_70 ( .A(gnd), .Y(_310_) );
NAND2X1 NAND2X1_31 ( .A(target[14]), .B(_310_), .Y(_311_) );
INVX2 INVX2_4 ( .A(target[15]), .Y(_312_) );
INVX1 INVX1_71 ( .A(target[14]), .Y(_313_) );
AOI22X1 AOI22X1_11 ( .A(_312_), .B(gnd), .C(_313_), .D(gnd), .Y(_314_) );
NAND3X1 NAND3X1_23 ( .A(_309_), .B(_311_), .C(_314_), .Y(_315_) );
INVX1 INVX1_72 ( .A(gnd), .Y(_316_) );
INVX1 INVX1_73 ( .A(gnd), .Y(_317_) );
AOI22X1 AOI22X1_12 ( .A(_316_), .B(target[13]), .C(target[12]), .D(_317_), .Y(_318_) );
INVX1 INVX1_74 ( .A(target[13]), .Y(_319_) );
NAND2X1 NAND2X1_32 ( .A(gnd), .B(_319_), .Y(_320_) );
INVX1 INVX1_75 ( .A(target[12]), .Y(_321_) );
NAND2X1 NAND2X1_33 ( .A(gnd), .B(_321_), .Y(_322_) );
NAND3X1 NAND3X1_24 ( .A(_320_), .B(_322_), .C(_318_), .Y(_323_) );
NOR2X1 NOR2X1_51 ( .A(_315_), .B(_323_), .Y(_324_) );
XNOR2X1 XNOR2X1_7 ( .A(gnd), .B(target[11]), .Y(_325_) );
INVX2 INVX2_5 ( .A(target[10]), .Y(_326_) );
OR2X2 OR2X2_6 ( .A(_326_), .B(gnd), .Y(_327_) );
NAND2X1 NAND2X1_34 ( .A(gnd), .B(_326_), .Y(_328_) );
NAND3X1 NAND3X1_25 ( .A(_327_), .B(_328_), .C(_325_), .Y(_329_) );
INVX1 INVX1_76 ( .A(gnd), .Y(_330_) );
INVX1 INVX1_77 ( .A(gnd), .Y(_331_) );
AOI22X1 AOI22X1_13 ( .A(_330_), .B(target[9]), .C(target[8]), .D(_331_), .Y(_332_) );
INVX1 INVX1_78 ( .A(target[9]), .Y(_333_) );
NAND2X1 NAND2X1_35 ( .A(gnd), .B(_333_), .Y(_334_) );
INVX1 INVX1_79 ( .A(target[8]), .Y(_335_) );
NAND2X1 NAND2X1_36 ( .A(gnd), .B(_335_), .Y(_336_) );
NAND3X1 NAND3X1_26 ( .A(_334_), .B(_336_), .C(_332_), .Y(_337_) );
NOR2X1 NOR2X1_52 ( .A(_337_), .B(_329_), .Y(_338_) );
AND2X2 AND2X2_7 ( .A(_338_), .B(_324_), .Y(_339_) );
XOR2X1 XOR2X1_4 ( .A(gnd), .B(target[7]), .Y(_340_) );
XOR2X1 XOR2X1_5 ( .A(target[6]), .B(gnd), .Y(_341_) );
NOR2X1 NOR2X1_53 ( .A(_340_), .B(_341_), .Y(_342_) );
INVX1 INVX1_80 ( .A(gnd), .Y(_343_) );
INVX1 INVX1_81 ( .A(gnd), .Y(_344_) );
AOI22X1 AOI22X1_14 ( .A(_343_), .B(target[5]), .C(target[4]), .D(_344_), .Y(_345_) );
INVX1 INVX1_82 ( .A(target[5]), .Y(_346_) );
INVX1 INVX1_83 ( .A(target[4]), .Y(_347_) );
AOI22X1 AOI22X1_15 ( .A(_346_), .B(gnd), .C(_347_), .D(gnd), .Y(_348_) );
AND2X2 AND2X2_8 ( .A(_345_), .B(_348_), .Y(_349_) );
NAND2X1 NAND2X1_37 ( .A(_342_), .B(_349_), .Y(_350_) );
NOR2X1 NOR2X1_54 ( .A(target[3]), .B(gnd), .Y(_351_) );
INVX1 INVX1_84 ( .A(_351_), .Y(_352_) );
NAND2X1 NAND2X1_38 ( .A(target[3]), .B(gnd), .Y(_353_) );
XOR2X1 XOR2X1_6 ( .A(target[2]), .B(gnd), .Y(_354_) );
AOI21X1 AOI21X1_41 ( .A(_352_), .B(_353_), .C(_354_), .Y(_355_) );
INVX1 INVX1_85 ( .A(gnd), .Y(_356_) );
NAND2X1 NAND2X1_39 ( .A(target[1]), .B(_356_), .Y(_357_) );
NOR2X1 NOR2X1_55 ( .A(target[1]), .B(_356_), .Y(_358_) );
INVX1 INVX1_86 ( .A(hash_array2_1), .Y(_359_) );
NOR2X1 NOR2X1_56 ( .A(target[0]), .B(_359_), .Y(_360_) );
OAI21X1 OAI21X1_45 ( .A(_358_), .B(_360_), .C(_357_), .Y(_361_) );
NAND2X1 NAND2X1_40 ( .A(_361_), .B(_355_), .Y(_362_) );
INVX1 INVX1_87 ( .A(target[3]), .Y(_363_) );
NOR2X1 NOR2X1_57 ( .A(gnd), .B(_363_), .Y(_364_) );
NAND2X1 NAND2X1_41 ( .A(gnd), .B(_363_), .Y(_365_) );
INVX1 INVX1_88 ( .A(target[2]), .Y(_366_) );
NOR2X1 NOR2X1_58 ( .A(gnd), .B(_366_), .Y(_367_) );
AOI21X1 AOI21X1_42 ( .A(_365_), .B(_367_), .C(_364_), .Y(_255_) );
AOI21X1 AOI21X1_43 ( .A(_255_), .B(_362_), .C(_350_), .Y(_256_) );
XNOR2X1 XNOR2X1_8 ( .A(gnd), .B(target[7]), .Y(_257_) );
XNOR2X1 XNOR2X1_9 ( .A(target[6]), .B(gnd), .Y(_258_) );
NAND2X1 NAND2X1_42 ( .A(_257_), .B(_258_), .Y(_259_) );
OAI22X1 OAI22X1_3 ( .A(_346_), .B(gnd), .C(_347_), .D(gnd), .Y(_260_) );
OAI21X1 OAI21X1_46 ( .A(_343_), .B(target[5]), .C(_260_), .Y(_261_) );
INVX1 INVX1_89 ( .A(target[7]), .Y(_262_) );
NOR2X1 NOR2X1_59 ( .A(gnd), .B(_262_), .Y(_263_) );
INVX1 INVX1_90 ( .A(target[6]), .Y(_264_) );
NOR2X1 NOR2X1_60 ( .A(gnd), .B(_264_), .Y(_265_) );
AOI21X1 AOI21X1_44 ( .A(_265_), .B(_257_), .C(_263_), .Y(_266_) );
OAI21X1 OAI21X1_47 ( .A(_259_), .B(_261_), .C(_266_), .Y(_267_) );
OAI21X1 OAI21X1_48 ( .A(_256_), .B(_267_), .C(_339_), .Y(_268_) );
INVX1 INVX1_91 ( .A(target[11]), .Y(_269_) );
NOR2X1 NOR2X1_61 ( .A(gnd), .B(_269_), .Y(_270_) );
NOR2X1 NOR2X1_62 ( .A(gnd), .B(_326_), .Y(_271_) );
AOI21X1 AOI21X1_45 ( .A(_271_), .B(_325_), .C(_270_), .Y(_272_) );
OAI22X1 OAI22X1_4 ( .A(_333_), .B(gnd), .C(_335_), .D(gnd), .Y(_273_) );
OAI21X1 OAI21X1_49 ( .A(_330_), .B(target[9]), .C(_273_), .Y(_274_) );
OAI21X1 OAI21X1_50 ( .A(_329_), .B(_274_), .C(_272_), .Y(_275_) );
NOR2X1 NOR2X1_63 ( .A(target[13]), .B(_316_), .Y(_276_) );
OR2X2 OR2X2_7 ( .A(_318_), .B(_276_), .Y(_277_) );
AOI21X1 AOI21X1_46 ( .A(_312_), .B(gnd), .C(_311_), .Y(_278_) );
OAI21X1 OAI21X1_51 ( .A(_312_), .B(gnd), .C(reset_bF_buf0), .Y(_279_) );
NOR2X1 NOR2X1_64 ( .A(_279_), .B(_278_), .Y(_280_) );
OAI21X1 OAI21X1_52 ( .A(_315_), .B(_277_), .C(_280_), .Y(_281_) );
AOI21X1 AOI21X1_47 ( .A(_324_), .B(_275_), .C(_281_), .Y(_282_) );
INVX1 INVX1_92 ( .A(reset_bF_buf5), .Y(_283_) );
NAND2X1 NAND2X1_43 ( .A(compare_hash_1_compare_var_0_), .B(_283_), .Y(_284_) );
NAND2X1 NAND2X1_44 ( .A(_324_), .B(_338_), .Y(_285_) );
NAND2X1 NAND2X1_45 ( .A(_345_), .B(_348_), .Y(_286_) );
NOR2X1 NOR2X1_65 ( .A(_286_), .B(_259_), .Y(_287_) );
INVX1 INVX1_93 ( .A(_353_), .Y(_288_) );
XNOR2X1 XNOR2X1_10 ( .A(target[2]), .B(gnd), .Y(_289_) );
OAI21X1 OAI21X1_53 ( .A(_351_), .B(_288_), .C(_289_), .Y(_290_) );
XNOR2X1 XNOR2X1_11 ( .A(target[1]), .B(gnd), .Y(_291_) );
XNOR2X1 XNOR2X1_12 ( .A(target[0]), .B(hash_array2_1), .Y(_292_) );
NAND2X1 NAND2X1_46 ( .A(_291_), .B(_292_), .Y(_293_) );
NOR2X1 NOR2X1_66 ( .A(_293_), .B(_290_), .Y(_294_) );
NAND2X1 NAND2X1_47 ( .A(_287_), .B(_294_), .Y(_295_) );
OAI21X1 OAI21X1_54 ( .A(_285_), .B(_295_), .C(reset_bF_buf4), .Y(_296_) );
AOI22X1 AOI22X1_16 ( .A(_284_), .B(_296_), .C(_268_), .D(_282_), .Y(_254__0_) );
OR2X2 OR2X2_8 ( .A(reset_bF_buf3), .B(compare_hash_1_compare_var_1_), .Y(_297_) );
AND2X2 AND2X2_9 ( .A(_296_), .B(_297_), .Y(_254__1_) );
INVX1 INVX1_94 ( .A(compare_hash_1_compare_var_2_), .Y(_298_) );
INVX1 INVX1_95 ( .A(target[1]), .Y(_299_) );
NOR2X1 NOR2X1_67 ( .A(gnd), .B(_299_), .Y(_300_) );
NAND2X1 NAND2X1_48 ( .A(gnd), .B(_299_), .Y(_301_) );
INVX1 INVX1_96 ( .A(target[0]), .Y(_302_) );
NAND2X1 NAND2X1_49 ( .A(hash_array2_1), .B(_302_), .Y(_303_) );
AOI21X1 AOI21X1_48 ( .A(_301_), .B(_303_), .C(_300_), .Y(_304_) );
OAI21X1 OAI21X1_55 ( .A(_290_), .B(_304_), .C(_255_), .Y(_305_) );
AOI21X1 AOI21X1_49 ( .A(_287_), .B(_305_), .C(_267_), .Y(_306_) );
OAI21X1 OAI21X1_56 ( .A(_306_), .B(_285_), .C(_282_), .Y(_307_) );
OAI21X1 OAI21X1_57 ( .A(reset_bF_buf2), .B(_298_), .C(_307_), .Y(_254__2_) );
DFFPOSX1 DFFPOSX1_64 ( .CLK(clk_bF_buf8), .D(_254__0_), .Q(compare_hash_1_compare_var_0_) );
DFFPOSX1 DFFPOSX1_65 ( .CLK(clk_bF_buf7), .D(_254__1_), .Q(compare_hash_1_compare_var_1_) );
DFFPOSX1 DFFPOSX1_66 ( .CLK(clk_bF_buf6), .D(_254__2_), .Q(compare_hash_1_compare_var_2_) );
INVX2 INVX2_6 ( .A(loop_limit_inst_compare_inst_number0_0_), .Y(_412_) );
NOR2X1 NOR2X1_68 ( .A(loop_limit_inst_compare_inst_compare_var_0_), .B(loop_limit_inst_compare_inst_compare_var_1_), .Y(_413_) );
OR2X2 OR2X2_9 ( .A(_413_), .B(loop_limit_inst_compare_inst_compare_var_2_), .Y(_414_) );
NAND2X1 NAND2X1_50 ( .A(loop_limit_inst_compare_inst_compare_var_0_), .B(loop_limit_inst_compare_inst_compare_var_1_), .Y(_415_) );
INVX1 INVX1_97 ( .A(reset_bF_buf1), .Y(_416_) );
NOR2X1 NOR2X1_69 ( .A(loop_limit_inst_stop), .B(_416_), .Y(_417_) );
NAND2X1 NAND2X1_51 ( .A(_415_), .B(_417__bF_buf3), .Y(_418_) );
NOR2X1 NOR2X1_70 ( .A(_414_), .B(_418_), .Y(_419_) );
AND2X2 AND2X2_10 ( .A(_419_), .B(_412_), .Y(_368__0_) );
INVX1 INVX1_98 ( .A(loop_limit_inst_compare_inst_number0_1_), .Y(_420_) );
OAI21X1 OAI21X1_58 ( .A(_412_), .B(_420_), .C(_419_), .Y(_421_) );
AOI21X1 AOI21X1_50 ( .A(_412_), .B(_420_), .C(_421_), .Y(_368__1_) );
AOI21X1 AOI21X1_51 ( .A(loop_limit_inst_compare_inst_number0_0_), .B(loop_limit_inst_compare_inst_number0_1_), .C(loop_limit_inst_compare_inst_number0_2_), .Y(_422_) );
NAND3X1 NAND3X1_27 ( .A(loop_limit_inst_compare_inst_number0_0_), .B(loop_limit_inst_compare_inst_number0_1_), .C(loop_limit_inst_compare_inst_number0_2_), .Y(_423_) );
NAND2X1 NAND2X1_52 ( .A(_423_), .B(_419_), .Y(_424_) );
NOR2X1 NOR2X1_71 ( .A(_422_), .B(_424_), .Y(_368__2_) );
INVX2 INVX2_7 ( .A(loop_limit_inst_compare_inst_number0_3_), .Y(_425_) );
OAI21X1 OAI21X1_59 ( .A(_425_), .B(_423_), .C(_419_), .Y(_426_) );
AOI21X1 AOI21X1_52 ( .A(_425_), .B(_423_), .C(_426_), .Y(_368__3_) );
INVX1 INVX1_99 ( .A(loop_limit_inst_compare_inst_number0_4_), .Y(_427_) );
NOR3X1 NOR3X1_1 ( .A(_425_), .B(_427_), .C(_423_), .Y(_428_) );
OAI21X1 OAI21X1_60 ( .A(_423_), .B(_425_), .C(_427_), .Y(_429_) );
NAND2X1 NAND2X1_53 ( .A(_429_), .B(_419_), .Y(_430_) );
NOR2X1 NOR2X1_72 ( .A(_428_), .B(_430_), .Y(_368__4_) );
NAND2X1 NAND2X1_54 ( .A(loop_limit_inst_compare_inst_number0_5_), .B(_428_), .Y(_431_) );
INVX1 INVX1_100 ( .A(_431_), .Y(_432_) );
OAI21X1 OAI21X1_61 ( .A(loop_limit_inst_compare_inst_number0_5_), .B(_428_), .C(_419_), .Y(_433_) );
NOR2X1 NOR2X1_73 ( .A(_432_), .B(_433_), .Y(_368__5_) );
NAND3X1 NAND3X1_28 ( .A(loop_limit_inst_compare_inst_number0_5_), .B(loop_limit_inst_compare_inst_number0_6_), .C(_428_), .Y(_371_) );
INVX1 INVX1_101 ( .A(_371_), .Y(_372_) );
OAI21X1 OAI21X1_62 ( .A(_432_), .B(loop_limit_inst_compare_inst_number0_6_), .C(_419_), .Y(_373_) );
NOR2X1 NOR2X1_74 ( .A(_372_), .B(_373_), .Y(_368__6_) );
INVX1 INVX1_102 ( .A(loop_limit_inst_compare_inst_number0_7_), .Y(_374_) );
NOR2X1 NOR2X1_75 ( .A(_374_), .B(_371_), .Y(_375_) );
OAI21X1 OAI21X1_63 ( .A(_372_), .B(loop_limit_inst_compare_inst_number0_7_), .C(_419_), .Y(_376_) );
NOR2X1 NOR2X1_76 ( .A(_375_), .B(_376_), .Y(_368__7_) );
INVX1 INVX1_103 ( .A(loop_limit_inst_compare_inst_number0_8_), .Y(_377_) );
NOR3X1 NOR3X1_2 ( .A(_374_), .B(_377_), .C(_371_), .Y(_378_) );
OAI21X1 OAI21X1_64 ( .A(_375_), .B(loop_limit_inst_compare_inst_number0_8_), .C(_419_), .Y(_379_) );
NOR2X1 NOR2X1_77 ( .A(_378_), .B(_379_), .Y(_368__8_) );
NAND2X1 NAND2X1_55 ( .A(loop_limit_inst_compare_inst_number0_9_), .B(_378_), .Y(_380_) );
INVX1 INVX1_104 ( .A(_380_), .Y(_381_) );
OAI21X1 OAI21X1_65 ( .A(_378_), .B(loop_limit_inst_compare_inst_number0_9_), .C(_419_), .Y(_382_) );
NOR2X1 NOR2X1_78 ( .A(_382_), .B(_381_), .Y(_368__9_) );
NAND3X1 NAND3X1_29 ( .A(loop_limit_inst_compare_inst_number0_9_), .B(loop_limit_inst_compare_inst_number0_10_), .C(_378_), .Y(_383_) );
INVX1 INVX1_105 ( .A(_383_), .Y(_384_) );
OAI21X1 OAI21X1_66 ( .A(_381_), .B(loop_limit_inst_compare_inst_number0_10_), .C(_419_), .Y(_385_) );
NOR2X1 NOR2X1_79 ( .A(_384_), .B(_385_), .Y(_368__10_) );
INVX1 INVX1_106 ( .A(loop_limit_inst_compare_inst_number0_11_), .Y(_386_) );
NOR2X1 NOR2X1_80 ( .A(_386_), .B(_383_), .Y(_387_) );
OAI21X1 OAI21X1_67 ( .A(_384_), .B(loop_limit_inst_compare_inst_number0_11_), .C(_419_), .Y(_388_) );
NOR2X1 NOR2X1_81 ( .A(_387_), .B(_388_), .Y(_368__11_) );
INVX1 INVX1_107 ( .A(loop_limit_inst_compare_inst_number0_12_), .Y(_389_) );
NOR3X1 NOR3X1_3 ( .A(_386_), .B(_389_), .C(_383_), .Y(_390_) );
OAI21X1 OAI21X1_68 ( .A(_387_), .B(loop_limit_inst_compare_inst_number0_12_), .C(_419_), .Y(_391_) );
NOR2X1 NOR2X1_82 ( .A(_390_), .B(_391_), .Y(_368__12_) );
OAI21X1 OAI21X1_69 ( .A(_390_), .B(loop_limit_inst_compare_inst_number0_13_), .C(_419_), .Y(_392_) );
AOI21X1 AOI21X1_53 ( .A(loop_limit_inst_compare_inst_number0_13_), .B(_390_), .C(_392_), .Y(_368__13_) );
AOI21X1 AOI21X1_54 ( .A(loop_limit_inst_compare_inst_number0_13_), .B(_390_), .C(loop_limit_inst_compare_inst_number0_14_), .Y(_393_) );
NAND3X1 NAND3X1_30 ( .A(loop_limit_inst_compare_inst_number0_13_), .B(loop_limit_inst_compare_inst_number0_14_), .C(_390_), .Y(_394_) );
NAND2X1 NAND2X1_56 ( .A(_419_), .B(_394_), .Y(_395_) );
NOR2X1 NOR2X1_83 ( .A(_393_), .B(_395_), .Y(_368__14_) );
INVX1 INVX1_108 ( .A(loop_limit_inst_compare_inst_number0_15_), .Y(_396_) );
OAI21X1 OAI21X1_70 ( .A(_394_), .B(_396_), .C(_419_), .Y(_397_) );
AOI21X1 AOI21X1_55 ( .A(_396_), .B(_394_), .C(_397_), .Y(_368__15_) );
INVX1 INVX1_109 ( .A(loop_limit_inst_compare_inst_number1_0_), .Y(_398_) );
NOR2X1 NOR2X1_84 ( .A(_398_), .B(_417__bF_buf2), .Y(_370__0_) );
INVX1 INVX1_110 ( .A(loop_limit_inst_compare_inst_number1_1_), .Y(_399_) );
NOR2X1 NOR2X1_85 ( .A(_399_), .B(_417__bF_buf1), .Y(_370__1_) );
INVX1 INVX1_111 ( .A(loop_limit_inst_compare_inst_number1_2_), .Y(_400_) );
NOR2X1 NOR2X1_86 ( .A(_400_), .B(_417__bF_buf0), .Y(_370__2_) );
OR2X2 OR2X2_10 ( .A(_417__bF_buf3), .B(loop_limit_inst_compare_inst_number1_3_), .Y(_370__3_) );
INVX1 INVX1_112 ( .A(loop_limit_inst_compare_inst_number1_4_), .Y(_401_) );
NOR2X1 NOR2X1_87 ( .A(_401_), .B(_417__bF_buf2), .Y(_370__4_) );
INVX1 INVX1_113 ( .A(loop_limit_inst_compare_inst_number1_5_), .Y(_402_) );
NOR2X1 NOR2X1_88 ( .A(_402_), .B(_417__bF_buf1), .Y(_370__5_) );
INVX1 INVX1_114 ( .A(loop_limit_inst_compare_inst_number1_6_), .Y(_403_) );
NOR2X1 NOR2X1_89 ( .A(_403_), .B(_417__bF_buf0), .Y(_370__6_) );
OR2X2 OR2X2_11 ( .A(_417__bF_buf3), .B(loop_limit_inst_compare_inst_number1_7_), .Y(_370__7_) );
OR2X2 OR2X2_12 ( .A(_417__bF_buf2), .B(loop_limit_inst_compare_inst_number1_8_), .Y(_370__8_) );
OR2X2 OR2X2_13 ( .A(_417__bF_buf1), .B(loop_limit_inst_compare_inst_number1_9_), .Y(_370__9_) );
INVX1 INVX1_115 ( .A(loop_limit_inst_compare_inst_number1_10_), .Y(_404_) );
NOR2X1 NOR2X1_90 ( .A(_404_), .B(_417__bF_buf0), .Y(_370__10_) );
INVX1 INVX1_116 ( .A(loop_limit_inst_compare_inst_number1_11_), .Y(_405_) );
NOR2X1 NOR2X1_91 ( .A(_405_), .B(_417__bF_buf3), .Y(_370__11_) );
OR2X2 OR2X2_14 ( .A(_417__bF_buf2), .B(loop_limit_inst_compare_inst_number1_12_), .Y(_370__12_) );
INVX1 INVX1_117 ( .A(loop_limit_inst_compare_inst_number1_13_), .Y(_406_) );
NOR2X1 NOR2X1_92 ( .A(_406_), .B(_417__bF_buf1), .Y(_370__13_) );
INVX1 INVX1_118 ( .A(loop_limit_inst_compare_inst_number1_14_), .Y(_407_) );
NOR2X1 NOR2X1_93 ( .A(_407_), .B(_417__bF_buf0), .Y(_370__14_) );
INVX1 INVX1_119 ( .A(loop_limit_inst_compare_inst_number1_15_), .Y(_408_) );
NOR2X1 NOR2X1_94 ( .A(_408_), .B(_417__bF_buf3), .Y(_370__15_) );
INVX1 INVX1_120 ( .A(loop_limit_inst_stop), .Y(_409_) );
NAND2X1 NAND2X1_57 ( .A(loop_limit_inst_compare_inst_compare_var_2_), .B(_413_), .Y(_410_) );
OAI21X1 OAI21X1_71 ( .A(_409_), .B(fail), .C(reset_bF_buf0), .Y(_411_) );
AOI21X1 AOI21X1_56 ( .A(_409_), .B(_410_), .C(_411_), .Y(_369_) );
DFFPOSX1 DFFPOSX1_67 ( .CLK(clk_bF_buf5), .D(_369_), .Q(fail) );
DFFPOSX1 DFFPOSX1_68 ( .CLK(clk_bF_buf4), .D(_370__0_), .Q(loop_limit_inst_compare_inst_number1_0_) );
DFFPOSX1 DFFPOSX1_69 ( .CLK(clk_bF_buf3), .D(_370__1_), .Q(loop_limit_inst_compare_inst_number1_1_) );
DFFPOSX1 DFFPOSX1_70 ( .CLK(clk_bF_buf2), .D(_370__2_), .Q(loop_limit_inst_compare_inst_number1_2_) );
DFFPOSX1 DFFPOSX1_71 ( .CLK(clk_bF_buf1), .D(_370__3_), .Q(loop_limit_inst_compare_inst_number1_3_) );
DFFPOSX1 DFFPOSX1_72 ( .CLK(clk_bF_buf0), .D(_370__4_), .Q(loop_limit_inst_compare_inst_number1_4_) );
DFFPOSX1 DFFPOSX1_73 ( .CLK(clk_bF_buf11), .D(_370__5_), .Q(loop_limit_inst_compare_inst_number1_5_) );
DFFPOSX1 DFFPOSX1_74 ( .CLK(clk_bF_buf10), .D(_370__6_), .Q(loop_limit_inst_compare_inst_number1_6_) );
DFFPOSX1 DFFPOSX1_75 ( .CLK(clk_bF_buf9), .D(_370__7_), .Q(loop_limit_inst_compare_inst_number1_7_) );
DFFPOSX1 DFFPOSX1_76 ( .CLK(clk_bF_buf8), .D(_370__8_), .Q(loop_limit_inst_compare_inst_number1_8_) );
DFFPOSX1 DFFPOSX1_77 ( .CLK(clk_bF_buf7), .D(_370__9_), .Q(loop_limit_inst_compare_inst_number1_9_) );
DFFPOSX1 DFFPOSX1_78 ( .CLK(clk_bF_buf6), .D(_370__10_), .Q(loop_limit_inst_compare_inst_number1_10_) );
DFFPOSX1 DFFPOSX1_79 ( .CLK(clk_bF_buf5), .D(_370__11_), .Q(loop_limit_inst_compare_inst_number1_11_) );
DFFPOSX1 DFFPOSX1_80 ( .CLK(clk_bF_buf4), .D(_370__12_), .Q(loop_limit_inst_compare_inst_number1_12_) );
DFFPOSX1 DFFPOSX1_81 ( .CLK(clk_bF_buf3), .D(_370__13_), .Q(loop_limit_inst_compare_inst_number1_13_) );
DFFPOSX1 DFFPOSX1_82 ( .CLK(clk_bF_buf2), .D(_370__14_), .Q(loop_limit_inst_compare_inst_number1_14_) );
DFFPOSX1 DFFPOSX1_83 ( .CLK(clk_bF_buf1), .D(_370__15_), .Q(loop_limit_inst_compare_inst_number1_15_) );
DFFPOSX1 DFFPOSX1_84 ( .CLK(clk_bF_buf0), .D(_368__0_), .Q(current_loop_actualize_0_) );
DFFPOSX1 DFFPOSX1_85 ( .CLK(clk_bF_buf11), .D(_368__1_), .Q(current_loop_actualize_1_) );
DFFPOSX1 DFFPOSX1_86 ( .CLK(clk_bF_buf10), .D(_368__2_), .Q(current_loop_actualize_2_) );
DFFPOSX1 DFFPOSX1_87 ( .CLK(clk_bF_buf9), .D(_368__3_), .Q(current_loop_actualize_3_) );
DFFPOSX1 DFFPOSX1_88 ( .CLK(clk_bF_buf8), .D(_368__4_), .Q(current_loop_actualize_4_) );
DFFPOSX1 DFFPOSX1_89 ( .CLK(clk_bF_buf7), .D(_368__5_), .Q(current_loop_actualize_5_) );
DFFPOSX1 DFFPOSX1_90 ( .CLK(clk_bF_buf6), .D(_368__6_), .Q(current_loop_actualize_6_) );
DFFPOSX1 DFFPOSX1_91 ( .CLK(clk_bF_buf5), .D(_368__7_), .Q(current_loop_actualize_7_) );
DFFPOSX1 DFFPOSX1_92 ( .CLK(clk_bF_buf4), .D(_368__8_), .Q(current_loop_actualize_8_) );
DFFPOSX1 DFFPOSX1_93 ( .CLK(clk_bF_buf3), .D(_368__9_), .Q(current_loop_actualize_9_) );
DFFPOSX1 DFFPOSX1_94 ( .CLK(clk_bF_buf2), .D(_368__10_), .Q(current_loop_actualize_10_) );
DFFPOSX1 DFFPOSX1_95 ( .CLK(clk_bF_buf1), .D(_368__11_), .Q(current_loop_actualize_11_) );
DFFPOSX1 DFFPOSX1_96 ( .CLK(clk_bF_buf0), .D(_368__12_), .Q(current_loop_actualize_12_) );
DFFPOSX1 DFFPOSX1_97 ( .CLK(clk_bF_buf11), .D(_368__13_), .Q(current_loop_actualize_13_) );
DFFPOSX1 DFFPOSX1_98 ( .CLK(clk_bF_buf10), .D(_368__14_), .Q(current_loop_actualize_14_) );
DFFPOSX1 DFFPOSX1_99 ( .CLK(clk_bF_buf9), .D(_368__15_), .Q(current_loop_actualize_15_) );
INVX1 INVX1_121 ( .A(loop_limit_inst_compare_inst_number0_15_), .Y(_488_) );
NAND2X1 NAND2X1_58 ( .A(loop_limit_inst_compare_inst_number1_15_), .B(_488_), .Y(_489_) );
INVX1 INVX1_122 ( .A(loop_limit_inst_compare_inst_number0_14_), .Y(_490_) );
NAND2X1 NAND2X1_59 ( .A(loop_limit_inst_compare_inst_number1_14_), .B(_490_), .Y(_491_) );
INVX2 INVX2_8 ( .A(loop_limit_inst_compare_inst_number1_15_), .Y(_492_) );
INVX1 INVX1_123 ( .A(loop_limit_inst_compare_inst_number1_14_), .Y(_493_) );
AOI22X1 AOI22X1_17 ( .A(_492_), .B(loop_limit_inst_compare_inst_number0_15_), .C(_493_), .D(loop_limit_inst_compare_inst_number0_14_), .Y(_494_) );
NAND3X1 NAND3X1_31 ( .A(_489_), .B(_491_), .C(_494_), .Y(_495_) );
INVX1 INVX1_124 ( .A(loop_limit_inst_compare_inst_number0_13_), .Y(_496_) );
INVX1 INVX1_125 ( .A(loop_limit_inst_compare_inst_number0_12_), .Y(_497_) );
AOI22X1 AOI22X1_18 ( .A(_496_), .B(loop_limit_inst_compare_inst_number1_13_), .C(loop_limit_inst_compare_inst_number1_12_), .D(_497_), .Y(_498_) );
INVX1 INVX1_126 ( .A(loop_limit_inst_compare_inst_number1_13_), .Y(_499_) );
NAND2X1 NAND2X1_60 ( .A(loop_limit_inst_compare_inst_number0_13_), .B(_499_), .Y(_500_) );
INVX1 INVX1_127 ( .A(loop_limit_inst_compare_inst_number1_12_), .Y(_501_) );
NAND2X1 NAND2X1_61 ( .A(loop_limit_inst_compare_inst_number0_12_), .B(_501_), .Y(_502_) );
NAND3X1 NAND3X1_32 ( .A(_500_), .B(_502_), .C(_498_), .Y(_503_) );
NOR2X1 NOR2X1_95 ( .A(_495_), .B(_503_), .Y(_504_) );
XNOR2X1 XNOR2X1_13 ( .A(loop_limit_inst_compare_inst_number0_11_), .B(loop_limit_inst_compare_inst_number1_11_), .Y(_505_) );
INVX2 INVX2_9 ( .A(loop_limit_inst_compare_inst_number1_10_), .Y(_506_) );
OR2X2 OR2X2_15 ( .A(_506_), .B(loop_limit_inst_compare_inst_number0_10_), .Y(_507_) );
NAND2X1 NAND2X1_62 ( .A(loop_limit_inst_compare_inst_number0_10_), .B(_506_), .Y(_508_) );
NAND3X1 NAND3X1_33 ( .A(_507_), .B(_508_), .C(_505_), .Y(_509_) );
INVX1 INVX1_128 ( .A(loop_limit_inst_compare_inst_number0_9_), .Y(_510_) );
INVX1 INVX1_129 ( .A(loop_limit_inst_compare_inst_number0_8_), .Y(_511_) );
AOI22X1 AOI22X1_19 ( .A(_510_), .B(loop_limit_inst_compare_inst_number1_9_), .C(loop_limit_inst_compare_inst_number1_8_), .D(_511_), .Y(_512_) );
INVX1 INVX1_130 ( .A(loop_limit_inst_compare_inst_number1_9_), .Y(_513_) );
NAND2X1 NAND2X1_63 ( .A(loop_limit_inst_compare_inst_number0_9_), .B(_513_), .Y(_514_) );
INVX1 INVX1_131 ( .A(loop_limit_inst_compare_inst_number1_8_), .Y(_515_) );
NAND2X1 NAND2X1_64 ( .A(loop_limit_inst_compare_inst_number0_8_), .B(_515_), .Y(_516_) );
NAND3X1 NAND3X1_34 ( .A(_514_), .B(_516_), .C(_512_), .Y(_517_) );
NOR2X1 NOR2X1_96 ( .A(_517_), .B(_509_), .Y(_518_) );
AND2X2 AND2X2_11 ( .A(_518_), .B(_504_), .Y(_519_) );
XOR2X1 XOR2X1_7 ( .A(loop_limit_inst_compare_inst_number0_7_), .B(loop_limit_inst_compare_inst_number1_7_), .Y(_520_) );
XOR2X1 XOR2X1_8 ( .A(loop_limit_inst_compare_inst_number1_6_), .B(loop_limit_inst_compare_inst_number0_6_), .Y(_521_) );
NOR2X1 NOR2X1_97 ( .A(_520_), .B(_521_), .Y(_522_) );
INVX1 INVX1_132 ( .A(loop_limit_inst_compare_inst_number0_5_), .Y(_523_) );
INVX1 INVX1_133 ( .A(loop_limit_inst_compare_inst_number0_4_), .Y(_524_) );
AOI22X1 AOI22X1_20 ( .A(_523_), .B(loop_limit_inst_compare_inst_number1_5_), .C(loop_limit_inst_compare_inst_number1_4_), .D(_524_), .Y(_525_) );
INVX1 INVX1_134 ( .A(loop_limit_inst_compare_inst_number1_5_), .Y(_526_) );
INVX1 INVX1_135 ( .A(loop_limit_inst_compare_inst_number1_4_), .Y(_527_) );
AOI22X1 AOI22X1_21 ( .A(_526_), .B(loop_limit_inst_compare_inst_number0_5_), .C(_527_), .D(loop_limit_inst_compare_inst_number0_4_), .Y(_528_) );
AND2X2 AND2X2_12 ( .A(_525_), .B(_528_), .Y(_529_) );
NAND2X1 NAND2X1_65 ( .A(_522_), .B(_529_), .Y(_530_) );
NOR2X1 NOR2X1_98 ( .A(loop_limit_inst_compare_inst_number1_3_), .B(loop_limit_inst_compare_inst_number0_3_), .Y(_531_) );
INVX1 INVX1_136 ( .A(_531_), .Y(_532_) );
NAND2X1 NAND2X1_66 ( .A(loop_limit_inst_compare_inst_number1_3_), .B(loop_limit_inst_compare_inst_number0_3_), .Y(_533_) );
XOR2X1 XOR2X1_9 ( .A(loop_limit_inst_compare_inst_number1_2_), .B(loop_limit_inst_compare_inst_number0_2_), .Y(_534_) );
AOI21X1 AOI21X1_57 ( .A(_532_), .B(_533_), .C(_534_), .Y(_535_) );
INVX1 INVX1_137 ( .A(loop_limit_inst_compare_inst_number0_1_), .Y(_536_) );
NAND2X1 NAND2X1_67 ( .A(loop_limit_inst_compare_inst_number1_1_), .B(_536_), .Y(_537_) );
NOR2X1 NOR2X1_99 ( .A(loop_limit_inst_compare_inst_number1_1_), .B(_536_), .Y(_538_) );
INVX1 INVX1_138 ( .A(loop_limit_inst_compare_inst_number0_0_), .Y(_539_) );
NOR2X1 NOR2X1_100 ( .A(loop_limit_inst_compare_inst_number1_0_), .B(_539_), .Y(_540_) );
OAI21X1 OAI21X1_72 ( .A(_538_), .B(_540_), .C(_537_), .Y(_541_) );
NAND2X1 NAND2X1_68 ( .A(_541_), .B(_535_), .Y(_542_) );
INVX1 INVX1_139 ( .A(loop_limit_inst_compare_inst_number1_3_), .Y(_543_) );
NOR2X1 NOR2X1_101 ( .A(loop_limit_inst_compare_inst_number0_3_), .B(_543_), .Y(_544_) );
NAND2X1 NAND2X1_69 ( .A(loop_limit_inst_compare_inst_number0_3_), .B(_543_), .Y(_545_) );
INVX1 INVX1_140 ( .A(loop_limit_inst_compare_inst_number1_2_), .Y(_546_) );
NOR2X1 NOR2X1_102 ( .A(loop_limit_inst_compare_inst_number0_2_), .B(_546_), .Y(_547_) );
AOI21X1 AOI21X1_58 ( .A(_545_), .B(_547_), .C(_544_), .Y(_435_) );
AOI21X1 AOI21X1_59 ( .A(_435_), .B(_542_), .C(_530_), .Y(_436_) );
XNOR2X1 XNOR2X1_14 ( .A(loop_limit_inst_compare_inst_number0_7_), .B(loop_limit_inst_compare_inst_number1_7_), .Y(_437_) );
XNOR2X1 XNOR2X1_15 ( .A(loop_limit_inst_compare_inst_number1_6_), .B(loop_limit_inst_compare_inst_number0_6_), .Y(_438_) );
NAND2X1 NAND2X1_70 ( .A(_437_), .B(_438_), .Y(_439_) );
OAI22X1 OAI22X1_5 ( .A(_526_), .B(loop_limit_inst_compare_inst_number0_5_), .C(_527_), .D(loop_limit_inst_compare_inst_number0_4_), .Y(_440_) );
OAI21X1 OAI21X1_73 ( .A(_523_), .B(loop_limit_inst_compare_inst_number1_5_), .C(_440_), .Y(_441_) );
INVX1 INVX1_141 ( .A(loop_limit_inst_compare_inst_number1_7_), .Y(_442_) );
NOR2X1 NOR2X1_103 ( .A(loop_limit_inst_compare_inst_number0_7_), .B(_442_), .Y(_443_) );
INVX1 INVX1_142 ( .A(loop_limit_inst_compare_inst_number1_6_), .Y(_444_) );
NOR2X1 NOR2X1_104 ( .A(loop_limit_inst_compare_inst_number0_6_), .B(_444_), .Y(_445_) );
AOI21X1 AOI21X1_60 ( .A(_445_), .B(_437_), .C(_443_), .Y(_446_) );
OAI21X1 OAI21X1_74 ( .A(_439_), .B(_441_), .C(_446_), .Y(_447_) );
OAI21X1 OAI21X1_75 ( .A(_436_), .B(_447_), .C(_519_), .Y(_448_) );
INVX1 INVX1_143 ( .A(loop_limit_inst_compare_inst_number1_11_), .Y(_449_) );
NOR2X1 NOR2X1_105 ( .A(loop_limit_inst_compare_inst_number0_11_), .B(_449_), .Y(_450_) );
NOR2X1 NOR2X1_106 ( .A(loop_limit_inst_compare_inst_number0_10_), .B(_506_), .Y(_451_) );
AOI21X1 AOI21X1_61 ( .A(_451_), .B(_505_), .C(_450_), .Y(_452_) );
OAI22X1 OAI22X1_6 ( .A(_513_), .B(loop_limit_inst_compare_inst_number0_9_), .C(_515_), .D(loop_limit_inst_compare_inst_number0_8_), .Y(_453_) );
OAI21X1 OAI21X1_76 ( .A(_510_), .B(loop_limit_inst_compare_inst_number1_9_), .C(_453_), .Y(_454_) );
OAI21X1 OAI21X1_77 ( .A(_509_), .B(_454_), .C(_452_), .Y(_455_) );
NOR2X1 NOR2X1_107 ( .A(loop_limit_inst_compare_inst_number1_13_), .B(_496_), .Y(_456_) );
OR2X2 OR2X2_16 ( .A(_498_), .B(_456_), .Y(_457_) );
AOI21X1 AOI21X1_62 ( .A(_492_), .B(loop_limit_inst_compare_inst_number0_15_), .C(_491_), .Y(_458_) );
OAI21X1 OAI21X1_78 ( .A(_492_), .B(loop_limit_inst_compare_inst_number0_15_), .C(reset_bF_buf5), .Y(_459_) );
NOR2X1 NOR2X1_108 ( .A(_459_), .B(_458_), .Y(_460_) );
OAI21X1 OAI21X1_79 ( .A(_495_), .B(_457_), .C(_460_), .Y(_461_) );
AOI21X1 AOI21X1_63 ( .A(_504_), .B(_455_), .C(_461_), .Y(_462_) );
INVX1 INVX1_144 ( .A(reset_bF_buf4), .Y(_463_) );
NAND2X1 NAND2X1_71 ( .A(loop_limit_inst_compare_inst_compare_var_0_), .B(_463_), .Y(_464_) );
NAND2X1 NAND2X1_72 ( .A(_504_), .B(_518_), .Y(_465_) );
NAND2X1 NAND2X1_73 ( .A(_525_), .B(_528_), .Y(_466_) );
NOR2X1 NOR2X1_109 ( .A(_466_), .B(_439_), .Y(_467_) );
INVX1 INVX1_145 ( .A(_533_), .Y(_468_) );
XNOR2X1 XNOR2X1_16 ( .A(loop_limit_inst_compare_inst_number1_2_), .B(loop_limit_inst_compare_inst_number0_2_), .Y(_469_) );
OAI21X1 OAI21X1_80 ( .A(_531_), .B(_468_), .C(_469_), .Y(_470_) );
XNOR2X1 XNOR2X1_17 ( .A(loop_limit_inst_compare_inst_number1_1_), .B(loop_limit_inst_compare_inst_number0_1_), .Y(_471_) );
XNOR2X1 XNOR2X1_18 ( .A(loop_limit_inst_compare_inst_number1_0_), .B(loop_limit_inst_compare_inst_number0_0_), .Y(_472_) );
NAND2X1 NAND2X1_74 ( .A(_471_), .B(_472_), .Y(_473_) );
NOR2X1 NOR2X1_110 ( .A(_473_), .B(_470_), .Y(_474_) );
NAND2X1 NAND2X1_75 ( .A(_467_), .B(_474_), .Y(_475_) );
OAI21X1 OAI21X1_81 ( .A(_465_), .B(_475_), .C(reset_bF_buf3), .Y(_476_) );
AOI22X1 AOI22X1_22 ( .A(_464_), .B(_476_), .C(_448_), .D(_462_), .Y(_434__0_) );
OR2X2 OR2X2_17 ( .A(reset_bF_buf2), .B(loop_limit_inst_compare_inst_compare_var_1_), .Y(_477_) );
AND2X2 AND2X2_13 ( .A(_476_), .B(_477_), .Y(_434__1_) );
INVX1 INVX1_146 ( .A(loop_limit_inst_compare_inst_compare_var_2_), .Y(_478_) );
INVX1 INVX1_147 ( .A(loop_limit_inst_compare_inst_number1_1_), .Y(_479_) );
NOR2X1 NOR2X1_111 ( .A(loop_limit_inst_compare_inst_number0_1_), .B(_479_), .Y(_480_) );
NAND2X1 NAND2X1_76 ( .A(loop_limit_inst_compare_inst_number0_1_), .B(_479_), .Y(_481_) );
INVX1 INVX1_148 ( .A(loop_limit_inst_compare_inst_number1_0_), .Y(_482_) );
NAND2X1 NAND2X1_77 ( .A(loop_limit_inst_compare_inst_number0_0_), .B(_482_), .Y(_483_) );
AOI21X1 AOI21X1_64 ( .A(_481_), .B(_483_), .C(_480_), .Y(_484_) );
OAI21X1 OAI21X1_82 ( .A(_470_), .B(_484_), .C(_435_), .Y(_485_) );
AOI21X1 AOI21X1_65 ( .A(_467_), .B(_485_), .C(_447_), .Y(_486_) );
OAI21X1 OAI21X1_83 ( .A(_486_), .B(_465_), .C(_462_), .Y(_487_) );
OAI21X1 OAI21X1_84 ( .A(reset_bF_buf1), .B(_478_), .C(_487_), .Y(_434__2_) );
DFFPOSX1 DFFPOSX1_100 ( .CLK(clk_bF_buf8), .D(_434__0_), .Q(loop_limit_inst_compare_inst_compare_var_0_) );
DFFPOSX1 DFFPOSX1_101 ( .CLK(clk_bF_buf7), .D(_434__1_), .Q(loop_limit_inst_compare_inst_compare_var_1_) );
DFFPOSX1 DFFPOSX1_102 ( .CLK(clk_bF_buf6), .D(_434__2_), .Q(loop_limit_inst_compare_inst_compare_var_2_) );
OAI21X1 OAI21X1_85 ( .A(micro_abc_calculation_ints_b_8_), .B(micro_abc_calculation_ints_c_16_), .C(reset_bF_buf0), .Y(_549_) );
AOI21X1 AOI21X1_66 ( .A(micro_abc_calculation_ints_b_8_), .B(micro_abc_calculation_ints_c_16_), .C(_549_), .Y(_548__0_) );
INVX1 INVX1_149 ( .A(micro_abc_calculation_ints_counter_3_), .Y(_550_) );
INVX1 INVX1_150 ( .A(micro_abc_calculation_ints_counter_2_), .Y(_551_) );
NOR2X1 NOR2X1_112 ( .A(_550_), .B(_551_), .Y(_552_) );
INVX2 INVX2_10 ( .A(micro_abc_calculation_ints_counter_0_), .Y(_553_) );
NOR2X1 NOR2X1_113 ( .A(micro_abc_calculation_ints_counter_1_), .B(_553_), .Y(_554_) );
NAND2X1 NAND2X1_78 ( .A(_554_), .B(_552_), .Y(_555_) );
NOR2X1 NOR2X1_114 ( .A(micro_abc_calculation_ints_counter_4_bF_buf4_), .B(_555_), .Y(_556_) );
INVX2 INVX2_11 ( .A(micro_abc_calculation_ints_counter_1_), .Y(_557_) );
NAND2X1 NAND2X1_79 ( .A(_557_), .B(_553_), .Y(_558_) );
INVX2 INVX2_12 ( .A(_558_), .Y(_559_) );
NAND2X1 NAND2X1_80 ( .A(_552_), .B(_559_), .Y(_560_) );
NOR2X1 NOR2X1_115 ( .A(micro_abc_calculation_ints_counter_4_bF_buf3_), .B(_560_), .Y(_561_) );
NOR2X1 NOR2X1_116 ( .A(micro_abc_calculation_ints_counter_2_), .B(_550_), .Y(_562_) );
NAND2X1 NAND2X1_81 ( .A(_554_), .B(_562_), .Y(_563_) );
NOR2X1 NOR2X1_117 ( .A(micro_abc_calculation_ints_counter_4_bF_buf2_), .B(_563_), .Y(_564_) );
INVX1 INVX1_151 ( .A(_564_), .Y(_565_) );
NAND2X1 NAND2X1_82 ( .A(_562_), .B(_559_), .Y(_566_) );
NOR2X1 NOR2X1_118 ( .A(micro_abc_calculation_ints_counter_4_bF_buf1_), .B(_566_), .Y(_567_) );
INVX1 INVX1_152 ( .A(_567_), .Y(_568_) );
NOR2X1 NOR2X1_119 ( .A(_557_), .B(_553_), .Y(_569_) );
NOR2X1 NOR2X1_120 ( .A(micro_abc_calculation_ints_counter_3_), .B(_551_), .Y(_570_) );
NAND2X1 NAND2X1_83 ( .A(_570_), .B(_569_), .Y(_571_) );
NOR2X1 NOR2X1_121 ( .A(micro_abc_calculation_ints_counter_4_bF_buf0_), .B(_571_), .Y(_572_) );
NAND2X1 NAND2X1_84 ( .A(_554_), .B(_570_), .Y(_573_) );
NOR2X1 NOR2X1_122 ( .A(micro_abc_calculation_ints_counter_4_bF_buf4_), .B(_573_), .Y(_574_) );
NAND2X1 NAND2X1_85 ( .A(_570_), .B(_559_), .Y(_575_) );
NOR2X1 NOR2X1_123 ( .A(micro_abc_calculation_ints_counter_4_bF_buf3_), .B(_575_), .Y(_576_) );
INVX1 INVX1_153 ( .A(_576_), .Y(_577_) );
NOR2X1 NOR2X1_124 ( .A(micro_abc_calculation_ints_counter_3_), .B(micro_abc_calculation_ints_counter_2_), .Y(_578_) );
NAND2X1 NAND2X1_86 ( .A(_578_), .B(_569_), .Y(_579_) );
NOR2X1 NOR2X1_125 ( .A(micro_abc_calculation_ints_counter_4_bF_buf2_), .B(_579_), .Y(_580_) );
NOR2X1 NOR2X1_126 ( .A(micro_abc_calculation_ints_k_0_), .B(micro_abc_calculation_ints_x_0_), .Y(_581_) );
AND2X2 AND2X2_14 ( .A(micro_abc_calculation_ints_k_0_), .B(micro_abc_calculation_ints_x_0_), .Y(_582_) );
NOR2X1 NOR2X1_127 ( .A(_581_), .B(_582_), .Y(_583_) );
NAND2X1 NAND2X1_87 ( .A(block3[0]), .B(_583__bF_buf6), .Y(_584_) );
INVX1 INVX1_154 ( .A(_584_), .Y(_585_) );
NOR2X1 NOR2X1_128 ( .A(block3[0]), .B(_583__bF_buf5), .Y(_586_) );
OAI21X1 OAI21X1_86 ( .A(_585_), .B(_586_), .C(_580_), .Y(_587_) );
NOR2X1 NOR2X1_129 ( .A(micro_abc_calculation_ints_counter_0_), .B(_557_), .Y(_588_) );
NAND2X1 NAND2X1_88 ( .A(_578_), .B(_588_), .Y(_589_) );
NOR2X1 NOR2X1_130 ( .A(micro_abc_calculation_ints_counter_4_bF_buf1_), .B(_589_), .Y(_590_) );
INVX8 INVX8_2 ( .A(micro_abc_calculation_ints_counter_4_bF_buf0_), .Y(_591_) );
AND2X2 AND2X2_15 ( .A(_554_), .B(_578_), .Y(_592_) );
NAND2X1 NAND2X1_89 ( .A(_591__bF_buf3), .B(_592_), .Y(_593_) );
INVX1 INVX1_155 ( .A(_593_), .Y(_594_) );
NAND2X1 NAND2X1_90 ( .A(block1[0]), .B(_583__bF_buf4), .Y(_595_) );
INVX1 INVX1_156 ( .A(_595_), .Y(_596_) );
NOR2X1 NOR2X1_131 ( .A(block1[0]), .B(_583__bF_buf3), .Y(_597_) );
OAI21X1 OAI21X1_87 ( .A(_596_), .B(_597_), .C(_594_), .Y(_598_) );
INVX1 INVX1_157 ( .A(micro_abc_calculation_ints_out_logic_final_16_), .Y(_599_) );
AND2X2 AND2X2_16 ( .A(_559_), .B(_578_), .Y(_600_) );
NAND2X1 NAND2X1_91 ( .A(_591__bF_buf2), .B(_600_), .Y(_601_) );
INVX1 INVX1_158 ( .A(_601_), .Y(_602_) );
NAND2X1 NAND2X1_92 ( .A(block0[0]), .B(_583__bF_buf2), .Y(_603_) );
INVX1 INVX1_159 ( .A(block0[0]), .Y(_604_) );
OAI21X1 OAI21X1_88 ( .A(_582_), .B(_581_), .C(_604_), .Y(_605_) );
NAND3X1 NAND3X1_35 ( .A(_603_), .B(_605_), .C(_602_), .Y(_606_) );
OAI21X1 OAI21X1_89 ( .A(_599_), .B(_602_), .C(_606_), .Y(_607_) );
OAI21X1 OAI21X1_90 ( .A(_607_), .B(_594_), .C(_598_), .Y(_608_) );
NOR2X1 NOR2X1_132 ( .A(_590_), .B(_608_), .Y(_609_) );
INVX1 INVX1_160 ( .A(_580_), .Y(_610_) );
INVX1 INVX1_161 ( .A(_590_), .Y(_611_) );
XNOR2X1 XNOR2X1_19 ( .A(_583__bF_buf1), .B(block2[0]), .Y(_612_) );
OAI21X1 OAI21X1_91 ( .A(_611_), .B(_612_), .C(_610_), .Y(_613_) );
OAI21X1 OAI21X1_92 ( .A(_609_), .B(_613_), .C(_587_), .Y(_614_) );
XNOR2X1 XNOR2X1_20 ( .A(_583__bF_buf0), .B(block4[0]), .Y(_615_) );
MUX2X1 MUX2X1_1 ( .A(_614_), .B(_615_), .S(_577_), .Y(_616_) );
NAND2X1 NAND2X1_93 ( .A(_570_), .B(_588_), .Y(_617_) );
NOR2X1 NOR2X1_133 ( .A(micro_abc_calculation_ints_counter_4_bF_buf4_), .B(_617_), .Y(_618_) );
XNOR2X1 XNOR2X1_21 ( .A(_583__bF_buf6), .B(block5[0]), .Y(_619_) );
AOI21X1 AOI21X1_67 ( .A(_574_), .B(_619_), .C(_618_), .Y(_620_) );
OAI21X1 OAI21X1_93 ( .A(_616_), .B(_574_), .C(_620_), .Y(_621_) );
NAND2X1 NAND2X1_94 ( .A(block6[0]), .B(_583__bF_buf5), .Y(_622_) );
INVX1 INVX1_162 ( .A(_622_), .Y(_623_) );
OAI21X1 OAI21X1_94 ( .A(block6[0]), .B(_583__bF_buf4), .C(_618_), .Y(_624_) );
OAI21X1 OAI21X1_95 ( .A(_623_), .B(_624_), .C(_621_), .Y(_625_) );
NOR2X1 NOR2X1_134 ( .A(block7[0]), .B(_583__bF_buf3), .Y(_626_) );
INVX1 INVX1_163 ( .A(block7[0]), .Y(_627_) );
INVX4 INVX4_1 ( .A(_583__bF_buf2), .Y(_628_) );
NOR2X1 NOR2X1_135 ( .A(_627_), .B(_628_), .Y(_629_) );
OAI21X1 OAI21X1_96 ( .A(_629_), .B(_626_), .C(_572_), .Y(_630_) );
OAI21X1 OAI21X1_97 ( .A(_625_), .B(_572_), .C(_630_), .Y(_631_) );
NAND2X1 NAND2X1_95 ( .A(block8[0]), .B(_583__bF_buf1), .Y(_632_) );
OR2X2 OR2X2_18 ( .A(_583__bF_buf0), .B(block8[0]), .Y(_633_) );
AOI21X1 AOI21X1_68 ( .A(_632_), .B(_633_), .C(_568_), .Y(_634_) );
AOI21X1 AOI21X1_69 ( .A(_568_), .B(_631_), .C(_634_), .Y(_635_) );
NAND2X1 NAND2X1_96 ( .A(_588_), .B(_562_), .Y(_636_) );
NOR2X1 NOR2X1_136 ( .A(micro_abc_calculation_ints_counter_4_bF_buf3_), .B(_636_), .Y(_637_) );
INVX1 INVX1_164 ( .A(_637_), .Y(_638_) );
NOR2X1 NOR2X1_137 ( .A(block9[0]), .B(_583__bF_buf6), .Y(_639_) );
INVX1 INVX1_165 ( .A(block9[0]), .Y(_640_) );
OAI21X1 OAI21X1_98 ( .A(_640_), .B(_628_), .C(_564_), .Y(_641_) );
OAI21X1 OAI21X1_99 ( .A(_641_), .B(_639_), .C(_638_), .Y(_642_) );
AOI21X1 AOI21X1_70 ( .A(_565_), .B(_635_), .C(_642_), .Y(_643_) );
NAND2X1 NAND2X1_97 ( .A(_562_), .B(_569_), .Y(_644_) );
AND2X2 AND2X2_17 ( .A(_583__bF_buf5), .B(block10[0]), .Y(_645_) );
NOR2X1 NOR2X1_138 ( .A(block10[0]), .B(_583__bF_buf4), .Y(_646_) );
OAI21X1 OAI21X1_100 ( .A(_645_), .B(_646_), .C(_637_), .Y(_647_) );
OAI21X1 OAI21X1_101 ( .A(micro_abc_calculation_ints_counter_4_bF_buf2_), .B(_644_), .C(_647_), .Y(_648_) );
INVX1 INVX1_166 ( .A(block11[0]), .Y(_649_) );
NOR2X1 NOR2X1_139 ( .A(_649_), .B(_628_), .Y(_650_) );
NOR2X1 NOR2X1_140 ( .A(micro_abc_calculation_ints_counter_4_bF_buf1_), .B(_644_), .Y(_651_) );
OAI21X1 OAI21X1_102 ( .A(block11[0]), .B(_583__bF_buf3), .C(_651_), .Y(_652_) );
OAI22X1 OAI22X1_7 ( .A(_650_), .B(_652_), .C(_643_), .D(_648_), .Y(_653_) );
NAND2X1 NAND2X1_98 ( .A(nonce_2_0), .B(_583__bF_buf2), .Y(_654_) );
INVX1 INVX1_167 ( .A(_654_), .Y(_655_) );
NOR2X1 NOR2X1_141 ( .A(nonce_2_0), .B(_583__bF_buf1), .Y(_656_) );
OAI21X1 OAI21X1_103 ( .A(_655_), .B(_656_), .C(_561_), .Y(_657_) );
OAI21X1 OAI21X1_104 ( .A(_653_), .B(_561_), .C(_657_), .Y(_658_) );
NAND2X1 NAND2X1_99 ( .A(_588_), .B(_552_), .Y(_659_) );
NOR2X1 NOR2X1_142 ( .A(micro_abc_calculation_ints_counter_4_bF_buf0_), .B(_659_), .Y(_660_) );
NOR2X1 NOR2X1_143 ( .A(nonce_2_1), .B(_583__bF_buf0), .Y(_661_) );
NAND2X1 NAND2X1_100 ( .A(nonce_2_1), .B(_583__bF_buf6), .Y(_662_) );
INVX1 INVX1_168 ( .A(_662_), .Y(_663_) );
NOR2X1 NOR2X1_144 ( .A(_661_), .B(_663_), .Y(_664_) );
AOI21X1 AOI21X1_71 ( .A(_556_), .B(_664_), .C(_660_), .Y(_665_) );
OAI21X1 OAI21X1_105 ( .A(_658_), .B(_556_), .C(_665_), .Y(_666_) );
NAND2X1 NAND2X1_101 ( .A(_552_), .B(_569_), .Y(_667_) );
NOR2X1 NOR2X1_145 ( .A(micro_abc_calculation_ints_counter_4_bF_buf4_), .B(_667_), .Y(_668_) );
INVX1 INVX1_169 ( .A(_668_), .Y(_669_) );
AND2X2 AND2X2_18 ( .A(_583__bF_buf5), .B(nonce_2_2), .Y(_670_) );
NOR2X1 NOR2X1_146 ( .A(nonce_2_2), .B(_583__bF_buf4), .Y(_671_) );
OAI21X1 OAI21X1_106 ( .A(_670_), .B(_671_), .C(_660_), .Y(_672_) );
NAND3X1 NAND3X1_36 ( .A(_669_), .B(_672_), .C(_666_), .Y(_673_) );
INVX1 INVX1_170 ( .A(nonce_2_3), .Y(_674_) );
OAI21X1 OAI21X1_107 ( .A(_582_), .B(_581_), .C(_674_), .Y(_675_) );
NOR2X1 NOR2X1_147 ( .A(_674_), .B(_628_), .Y(_676_) );
NOR2X1 NOR2X1_148 ( .A(_667_), .B(_676_), .Y(_677_) );
AOI21X1 AOI21X1_72 ( .A(_675_), .B(_677_), .C(micro_abc_calculation_ints_counter_4_bF_buf3_), .Y(_678_) );
NOR2X1 NOR2X1_149 ( .A(_591__bF_buf1), .B(_659_), .Y(_679_) );
INVX1 INVX1_171 ( .A(_679_), .Y(_680_) );
NOR2X1 NOR2X1_150 ( .A(_591__bF_buf0), .B(_636_), .Y(_681_) );
NOR2X1 NOR2X1_151 ( .A(_591__bF_buf3), .B(_563_), .Y(_682_) );
NOR2X1 NOR2X1_152 ( .A(_591__bF_buf2), .B(_566_), .Y(_683_) );
NOR2X1 NOR2X1_153 ( .A(_591__bF_buf1), .B(_617_), .Y(_684_) );
NOR2X1 NOR2X1_154 ( .A(_591__bF_buf0), .B(_573_), .Y(_685_) );
INVX1 INVX1_172 ( .A(_685_), .Y(_686_) );
NOR2X1 NOR2X1_155 ( .A(_591__bF_buf3), .B(_575_), .Y(_687_) );
OR2X2 OR2X2_19 ( .A(_579_), .B(_591__bF_buf2), .Y(_688_) );
INVX1 INVX1_173 ( .A(_688_), .Y(_689_) );
NOR2X1 NOR2X1_156 ( .A(_591__bF_buf1), .B(_589_), .Y(_690_) );
NAND2X1 NAND2X1_102 ( .A(micro_abc_calculation_ints_imput_W2_logic_16_), .B(_583__bF_buf3), .Y(_691_) );
INVX1 INVX1_174 ( .A(_691_), .Y(_692_) );
NOR2X1 NOR2X1_157 ( .A(micro_abc_calculation_ints_imput_W2_logic_16_), .B(_583__bF_buf2), .Y(_693_) );
OAI21X1 OAI21X1_108 ( .A(_692_), .B(_693_), .C(_690_), .Y(_694_) );
INVX1 INVX1_175 ( .A(micro_abc_calculation_ints_imput_W2_logic_8_), .Y(_695_) );
NAND2X1 NAND2X1_103 ( .A(micro_abc_calculation_ints_counter_4_bF_buf2_), .B(_592_), .Y(_696_) );
INVX1 INVX1_176 ( .A(_696_), .Y(_697_) );
OAI21X1 OAI21X1_109 ( .A(_695_), .B(_628_), .C(_697_), .Y(_698_) );
AOI21X1 AOI21X1_73 ( .A(_695_), .B(_628_), .C(_698_), .Y(_699_) );
INVX1 INVX1_177 ( .A(_690_), .Y(_700_) );
OAI21X1 OAI21X1_110 ( .A(_697_), .B(_599_), .C(_700_), .Y(_701_) );
OAI21X1 OAI21X1_111 ( .A(_699_), .B(_701_), .C(_694_), .Y(_702_) );
NAND2X1 NAND2X1_104 ( .A(micro_abc_calculation_ints_imput_W2_logic_24_), .B(_583__bF_buf1), .Y(_703_) );
INVX1 INVX1_178 ( .A(micro_abc_calculation_ints_imput_W2_logic_24_), .Y(_704_) );
OAI21X1 OAI21X1_112 ( .A(_582_), .B(_581_), .C(_704_), .Y(_705_) );
NAND3X1 NAND3X1_37 ( .A(_703_), .B(_705_), .C(_689_), .Y(_706_) );
OAI21X1 OAI21X1_113 ( .A(_702_), .B(_689_), .C(_706_), .Y(_707_) );
NAND2X1 NAND2X1_105 ( .A(micro_abc_calculation_ints_imput_W2_logic_32_), .B(_583__bF_buf0), .Y(_708_) );
INVX1 INVX1_179 ( .A(_708_), .Y(_709_) );
NOR2X1 NOR2X1_158 ( .A(micro_abc_calculation_ints_imput_W2_logic_32_), .B(_583__bF_buf6), .Y(_710_) );
OAI21X1 OAI21X1_114 ( .A(_709_), .B(_710_), .C(_687_), .Y(_711_) );
OAI21X1 OAI21X1_115 ( .A(_707_), .B(_687_), .C(_711_), .Y(_712_) );
XNOR2X1 XNOR2X1_22 ( .A(_583__bF_buf5), .B(micro_abc_calculation_ints_imput_W2_logic_40_), .Y(_713_) );
MUX2X1 MUX2X1_2 ( .A(_712_), .B(_713_), .S(_686_), .Y(_714_) );
NOR2X1 NOR2X1_159 ( .A(_591__bF_buf0), .B(_571_), .Y(_715_) );
XNOR2X1 XNOR2X1_23 ( .A(_583__bF_buf4), .B(micro_abc_calculation_ints_imput_W2_logic_48_), .Y(_716_) );
AOI21X1 AOI21X1_74 ( .A(_684_), .B(_716_), .C(_715_), .Y(_717_) );
OAI21X1 OAI21X1_116 ( .A(_714_), .B(_684_), .C(_717_), .Y(_718_) );
NAND2X1 NAND2X1_106 ( .A(micro_abc_calculation_ints_imput_W2_logic_56_), .B(_583__bF_buf3), .Y(_719_) );
INVX1 INVX1_180 ( .A(_719_), .Y(_720_) );
OAI21X1 OAI21X1_117 ( .A(micro_abc_calculation_ints_imput_W2_logic_56_), .B(_583__bF_buf2), .C(_715_), .Y(_721_) );
OAI21X1 OAI21X1_118 ( .A(_720_), .B(_721_), .C(_718_), .Y(_722_) );
NAND2X1 NAND2X1_107 ( .A(micro_abc_calculation_ints_imput_W2_logic_64_), .B(_583__bF_buf1), .Y(_723_) );
INVX1 INVX1_181 ( .A(_723_), .Y(_724_) );
NOR2X1 NOR2X1_160 ( .A(micro_abc_calculation_ints_imput_W2_logic_64_), .B(_583__bF_buf0), .Y(_725_) );
OAI21X1 OAI21X1_119 ( .A(_724_), .B(_725_), .C(_683_), .Y(_726_) );
OAI21X1 OAI21X1_120 ( .A(_722_), .B(_683_), .C(_726_), .Y(_727_) );
AND2X2 AND2X2_19 ( .A(_583__bF_buf6), .B(micro_abc_calculation_ints_imput_W2_logic_72_), .Y(_728_) );
OAI21X1 OAI21X1_121 ( .A(micro_abc_calculation_ints_imput_W2_logic_72_), .B(_583__bF_buf5), .C(_682_), .Y(_729_) );
OAI22X1 OAI22X1_8 ( .A(_728_), .B(_729_), .C(_727_), .D(_682_), .Y(_730_) );
NOR2X1 NOR2X1_161 ( .A(_591__bF_buf3), .B(_644_), .Y(_731_) );
XNOR2X1 XNOR2X1_24 ( .A(_583__bF_buf4), .B(micro_abc_calculation_ints_imput_W2_logic_80_), .Y(_732_) );
AOI21X1 AOI21X1_75 ( .A(_681_), .B(_732_), .C(_731_), .Y(_733_) );
OAI21X1 OAI21X1_122 ( .A(_730_), .B(_681_), .C(_733_), .Y(_734_) );
NOR2X1 NOR2X1_162 ( .A(_591__bF_buf2), .B(_560_), .Y(_735_) );
NOR2X1 NOR2X1_163 ( .A(micro_abc_calculation_ints_imput_W2_logic_88_), .B(_583__bF_buf3), .Y(_736_) );
NAND2X1 NAND2X1_108 ( .A(micro_abc_calculation_ints_imput_W2_logic_88_), .B(_583__bF_buf2), .Y(_737_) );
INVX1 INVX1_182 ( .A(_737_), .Y(_738_) );
NOR2X1 NOR2X1_164 ( .A(_736_), .B(_738_), .Y(_739_) );
AOI21X1 AOI21X1_76 ( .A(_731_), .B(_739_), .C(_735_), .Y(_740_) );
AND2X2 AND2X2_20 ( .A(_583__bF_buf1), .B(micro_abc_calculation_ints_imput_W2_logic_96_), .Y(_741_) );
NOR2X1 NOR2X1_165 ( .A(micro_abc_calculation_ints_imput_W2_logic_96_), .B(_583__bF_buf0), .Y(_742_) );
OAI21X1 OAI21X1_123 ( .A(_741_), .B(_742_), .C(_735_), .Y(_743_) );
OAI21X1 OAI21X1_124 ( .A(_591__bF_buf1), .B(_555_), .C(_743_), .Y(_744_) );
AOI21X1 AOI21X1_77 ( .A(_740_), .B(_734_), .C(_744_), .Y(_745_) );
AND2X2 AND2X2_21 ( .A(_583__bF_buf6), .B(micro_abc_calculation_ints_imput_W2_logic_104_), .Y(_746_) );
NOR2X1 NOR2X1_166 ( .A(_591__bF_buf0), .B(_555_), .Y(_747_) );
OAI21X1 OAI21X1_125 ( .A(micro_abc_calculation_ints_imput_W2_logic_104_), .B(_583__bF_buf5), .C(_747_), .Y(_748_) );
NOR2X1 NOR2X1_167 ( .A(_746_), .B(_748_), .Y(_749_) );
OAI21X1 OAI21X1_126 ( .A(_745_), .B(_749_), .C(_680_), .Y(_750_) );
NOR2X1 NOR2X1_168 ( .A(_591__bF_buf3), .B(_667_), .Y(_751_) );
NOR2X1 NOR2X1_169 ( .A(micro_abc_calculation_ints_imput_W2_logic_112_), .B(_583__bF_buf4), .Y(_752_) );
NAND2X1 NAND2X1_109 ( .A(micro_abc_calculation_ints_imput_W2_logic_112_), .B(_583__bF_buf3), .Y(_753_) );
INVX1 INVX1_183 ( .A(_753_), .Y(_754_) );
NOR2X1 NOR2X1_170 ( .A(_752_), .B(_754_), .Y(_755_) );
AOI21X1 AOI21X1_78 ( .A(_679_), .B(_755_), .C(_751_), .Y(_756_) );
INVX1 INVX1_184 ( .A(_600_), .Y(_757_) );
AND2X2 AND2X2_22 ( .A(_583__bF_buf2), .B(micro_abc_calculation_ints_imput_W2_logic_120_), .Y(_758_) );
NOR2X1 NOR2X1_171 ( .A(micro_abc_calculation_ints_imput_W2_logic_120_), .B(_583__bF_buf1), .Y(_759_) );
OAI21X1 OAI21X1_127 ( .A(_758_), .B(_759_), .C(_751_), .Y(_760_) );
OAI21X1 OAI21X1_128 ( .A(_591__bF_buf2), .B(_757_), .C(_760_), .Y(_761_) );
AOI21X1 AOI21X1_79 ( .A(_756_), .B(_750_), .C(_761_), .Y(_762_) );
AND2X2 AND2X2_23 ( .A(_583__bF_buf0), .B(micro_abc_calculation_ints_imput_W2_logic_0_), .Y(_763_) );
OAI21X1 OAI21X1_129 ( .A(micro_abc_calculation_ints_imput_W2_logic_0_), .B(_583__bF_buf6), .C(_600_), .Y(_764_) );
OAI21X1 OAI21X1_130 ( .A(_764_), .B(_763_), .C(micro_abc_calculation_ints_counter_4_bF_buf1_), .Y(_765_) );
OAI21X1 OAI21X1_131 ( .A(_762_), .B(_765_), .C(reset_bF_buf5), .Y(_766_) );
AOI21X1 AOI21X1_80 ( .A(_678_), .B(_673_), .C(_766_), .Y(_548__16_) );
DFFPOSX1 DFFPOSX1_103 ( .CLK(clk_bF_buf5), .D(_548__0_), .Q(micro_abc_calculation_ints_out_logic_final_0_) );
DFFPOSX1 DFFPOSX1_104 ( .CLK(clk_bF_buf4), .D(gnd), .Q(micro_abc_calculation_ints_out_logic_final_8_) );
DFFPOSX1 DFFPOSX1_105 ( .CLK(clk_bF_buf3), .D(_548__16_), .Q(micro_abc_calculation_ints_out_logic_final_16_) );
AND2X2 AND2X2_24 ( .A(micro_abc_calculation_ints_counter_2_), .B(micro_abc_calculation_ints_counter_1_), .Y(_768_) );
AND2X2 AND2X2_25 ( .A(micro_abc_calculation_ints_counter_4_bF_buf0_), .B(micro_abc_calculation_ints_counter_3_), .Y(_769_) );
NAND3X1 NAND3X1_38 ( .A(micro_abc_calculation_ints_counter_0_), .B(_768_), .C(_769_), .Y(_770_) );
NAND2X1 NAND2X1_110 ( .A(micro_counter_inst_ready), .B(reset_bF_buf4), .Y(_771_) );
AOI21X1 AOI21X1_81 ( .A(micro_abc_calculation_ints_counter_0_), .B(_770_), .C(_771_), .Y(_767__0_) );
XNOR2X1 XNOR2X1_25 ( .A(micro_abc_calculation_ints_counter_0_), .B(micro_abc_calculation_ints_counter_1_), .Y(_772_) );
AOI21X1 AOI21X1_82 ( .A(_772_), .B(_770_), .C(_771_), .Y(_767__1_) );
NAND3X1 NAND3X1_39 ( .A(micro_abc_calculation_ints_counter_0_), .B(micro_abc_calculation_ints_counter_2_), .C(micro_abc_calculation_ints_counter_1_), .Y(_773_) );
INVX1 INVX1_185 ( .A(micro_abc_calculation_ints_counter_2_), .Y(_774_) );
NAND2X1 NAND2X1_111 ( .A(micro_abc_calculation_ints_counter_0_), .B(micro_abc_calculation_ints_counter_1_), .Y(_775_) );
NAND2X1 NAND2X1_112 ( .A(_774_), .B(_775_), .Y(_776_) );
NAND2X1 NAND2X1_113 ( .A(_773_), .B(_776_), .Y(_777_) );
AOI21X1 AOI21X1_83 ( .A(_770_), .B(_777_), .C(_771_), .Y(_767__2_) );
INVX2 INVX2_13 ( .A(micro_abc_calculation_ints_counter_3_), .Y(_778_) );
NOR3X1 NOR3X1_4 ( .A(micro_abc_calculation_ints_counter_4_bF_buf4_), .B(_778_), .C(_773_), .Y(_779_) );
AND2X2 AND2X2_26 ( .A(_773_), .B(_778_), .Y(_780_) );
NOR3X1 NOR3X1_5 ( .A(_780_), .B(_771_), .C(_779_), .Y(_767__3_) );
INVX1 INVX1_186 ( .A(micro_abc_calculation_ints_counter_4_bF_buf3_), .Y(_781_) );
OR2X2 OR2X2_20 ( .A(_773_), .B(_778_), .Y(_782_) );
AOI21X1 AOI21X1_84 ( .A(_781_), .B(_782_), .C(_771_), .Y(_767__4_) );
DFFPOSX1 DFFPOSX1_106 ( .CLK(clk_bF_buf2), .D(_767__0_), .Q(micro_abc_calculation_ints_counter_0_) );
DFFPOSX1 DFFPOSX1_107 ( .CLK(clk_bF_buf1), .D(_767__1_), .Q(micro_abc_calculation_ints_counter_1_) );
DFFPOSX1 DFFPOSX1_108 ( .CLK(clk_bF_buf0), .D(_767__2_), .Q(micro_abc_calculation_ints_counter_2_) );
DFFPOSX1 DFFPOSX1_109 ( .CLK(clk_bF_buf11), .D(_767__3_), .Q(micro_abc_calculation_ints_counter_3_) );
DFFPOSX1 DFFPOSX1_110 ( .CLK(clk_bF_buf10), .D(_767__4_), .Q(micro_abc_calculation_ints_counter_4_) );
NAND2X1 NAND2X1_114 ( .A(micro_abc_calculation_ints_counter_4_bF_buf2_), .B(micro_abc_calculation_ints_counter_3_), .Y(_793_) );
NAND3X1 NAND3X1_40 ( .A(micro_abc_calculation_ints_counter_2_), .B(micro_abc_calculation_ints_counter_1_), .C(micro_abc_calculation_ints_counter_0_), .Y(_794_) );
NOR2X1 NOR2X1_172 ( .A(_793_), .B(_794_), .Y(_795_) );
NAND2X1 NAND2X1_115 ( .A(reset_bF_buf3), .B(_795_), .Y(_783_) );
INVX1 INVX1_187 ( .A(micro_abc_calculation_ints_out_logic_final_16_), .Y(_796_) );
INVX1 INVX1_188 ( .A(micro_hash_final_ints_flag), .Y(_797_) );
NAND2X1 NAND2X1_116 ( .A(_797_), .B(_795_), .Y(_798_) );
OAI21X1 OAI21X1_132 ( .A(_798_), .B(hash_array2_2), .C(reset_bF_buf2), .Y(_799_) );
AOI21X1 AOI21X1_85 ( .A(_796_), .B(_798_), .C(_799_), .Y(_786__0_) );
INVX1 INVX1_189 ( .A(reset_bF_buf1), .Y(_800_) );
INVX1 INVX1_190 ( .A(_798_), .Y(_801_) );
OR2X2 OR2X2_21 ( .A(_794_), .B(_793_), .Y(_802_) );
NOR2X1 NOR2X1_173 ( .A(_797_), .B(_802_), .Y(_803_) );
NAND2X1 NAND2X1_117 ( .A(hash_array2_1), .B(_801_), .Y(_787_) );
INVX1 INVX1_191 ( .A(micro_abc_calculation_ints_out_logic_final_8_), .Y(_788_) );
MUX2X1 MUX2X1_3 ( .A(_803_), .B(_802_), .S(_788_), .Y(_789_) );
AOI21X1 AOI21X1_86 ( .A(_789_), .B(_787_), .C(_800_), .Y(_785__0_) );
NAND2X1 NAND2X1_118 ( .A(hash_array2_0), .B(_801_), .Y(_790_) );
INVX1 INVX1_192 ( .A(micro_abc_calculation_ints_out_logic_final_0_), .Y(_791_) );
MUX2X1 MUX2X1_4 ( .A(_803_), .B(_802_), .S(_791_), .Y(_792_) );
AOI21X1 AOI21X1_87 ( .A(_792_), .B(_790_), .C(_800_), .Y(_784__0_) );
DFFPOSX1 DFFPOSX1_111 ( .CLK(clk_bF_buf9), .D(_784__0_), .Q(hash_array2_0) );
DFFPOSX1 DFFPOSX1_112 ( .CLK(clk_bF_buf8), .D(_785__0_), .Q(hash_array2_1) );
DFFPOSX1 DFFPOSX1_113 ( .CLK(clk_bF_buf7), .D(_786__0_), .Q(hash_array2_2) );
DFFPOSX1 DFFPOSX1_114 ( .CLK(clk_bF_buf6), .D(_783_), .Q(micro_hash_final_ints_flag) );
AND2X2 AND2X2_27 ( .A(reset_bF_buf0), .B(micro_abc_calculation_ints_b_8_), .Y(_805__0_) );
OR2X2 OR2X2_22 ( .A(micro_abc_calculation_ints_counter_0_), .B(micro_abc_calculation_ints_counter_3_), .Y(_808_) );
OR2X2 OR2X2_23 ( .A(micro_abc_calculation_ints_counter_2_), .B(micro_abc_calculation_ints_counter_1_), .Y(_809_) );
OAI21X1 OAI21X1_133 ( .A(_808_), .B(_809_), .C(micro_abc_calculation_ints_counter_4_bF_buf1_), .Y(_810_) );
AND2X2 AND2X2_28 ( .A(micro_mod_x_k_inst_b_0_), .B(micro_mod_x_k_inst_a_0_), .Y(_811_) );
OAI21X1 OAI21X1_134 ( .A(micro_mod_x_k_inst_b_0_), .B(micro_mod_x_k_inst_a_0_), .C(reset_bF_buf5), .Y(_812_) );
AOI21X1 AOI21X1_88 ( .A(_811_), .B(_810_), .C(_812_), .Y(_807__0_) );
AND2X2 AND2X2_29 ( .A(reset_bF_buf4), .B(micro_abc_calculation_ints_a_0_), .Y(_804__0_) );
BUFX2 BUFX2_34 ( .A(reset_bF_buf3), .Y(_806__0_) );
DFFPOSX1 DFFPOSX1_115 ( .CLK(clk_bF_buf5), .D(_804__0_), .Q(micro_mod_x_k_inst_a_0_) );
DFFPOSX1 DFFPOSX1_116 ( .CLK(clk_bF_buf4), .D(_807__0_), .Q(micro_abc_calculation_ints_x_0_) );
DFFPOSX1 DFFPOSX1_117 ( .CLK(clk_bF_buf3), .D(_806__0_), .Q(micro_abc_calculation_ints_k_0_) );
DFFPOSX1 DFFPOSX1_118 ( .CLK(clk_bF_buf2), .D(_805__0_), .Q(micro_mod_x_k_inst_b_0_) );
INVX1 INVX1_193 ( .A(hash_array2_1), .Y(_814_) );
NAND2X1 NAND2X1_119 ( .A(micro_counter_inst_ready), .B(_814_), .Y(_813__8_) );
AND2X2 AND2X2_30 ( .A(micro_counter_inst_ready), .B(hash_array2_2), .Y(_813__16_) );
INVX1 INVX1_194 ( .A(hash_array2_0), .Y(_815_) );
NAND2X1 NAND2X1_120 ( .A(micro_counter_inst_ready), .B(_815_), .Y(_813__0_) );
DFFPOSX1 DFFPOSX1_119 ( .CLK(clk_bF_buf1), .D(_813__0_), .Q(micro_abc_calculation_ints_a_0_) );
DFFPOSX1 DFFPOSX1_120 ( .CLK(clk_bF_buf0), .D(_813__8_), .Q(micro_abc_calculation_ints_b_8_) );
DFFPOSX1 DFFPOSX1_121 ( .CLK(clk_bF_buf11), .D(_813__16_), .Q(micro_abc_calculation_ints_c_16_) );
INVX1 INVX1_195 ( .A(micro_abc_calculation_ints_imput_W2_logic_120_), .Y(_817_) );
NAND2X1 NAND2X1_121 ( .A(micro_abc_calculation_ints_counter_1_), .B(micro_abc_calculation_ints_counter_0_), .Y(_818_) );
INVX4 INVX4_2 ( .A(micro_abc_calculation_ints_counter_4_bF_buf0_), .Y(_819_) );
NAND3X1 NAND3X1_41 ( .A(micro_abc_calculation_ints_counter_3_), .B(micro_abc_calculation_ints_counter_2_), .C(_819_), .Y(_820_) );
OAI21X1 OAI21X1_135 ( .A(_820_), .B(_818_), .C(reset_bF_buf2), .Y(_821_) );
NOR2X1 NOR2X1_174 ( .A(_817_), .B(_821_), .Y(_816__120_) );
INVX8 INVX8_3 ( .A(reset_bF_buf1), .Y(_822_) );
INVX2 INVX2_14 ( .A(micro_abc_calculation_ints_counter_1_), .Y(_823_) );
NAND2X1 NAND2X1_122 ( .A(micro_abc_calculation_ints_counter_0_), .B(_823_), .Y(_824_) );
NOR2X1 NOR2X1_175 ( .A(_824_), .B(_820_), .Y(_825_) );
NAND2X1 NAND2X1_123 ( .A(nonce_2_2), .B(_825_), .Y(_826_) );
OAI21X1 OAI21X1_136 ( .A(_820_), .B(_824_), .C(micro_abc_calculation_ints_imput_W2_logic_104_), .Y(_827_) );
AOI21X1 AOI21X1_89 ( .A(_827_), .B(_826_), .C(_822_), .Y(_816__104_) );
INVX2 INVX2_15 ( .A(micro_abc_calculation_ints_counter_0_), .Y(_828_) );
NAND2X1 NAND2X1_124 ( .A(_823_), .B(_828_), .Y(_829_) );
NOR2X1 NOR2X1_176 ( .A(_829_), .B(_820_), .Y(_830_) );
NAND2X1 NAND2X1_125 ( .A(nonce_2_1), .B(_830_), .Y(_831_) );
OAI21X1 OAI21X1_137 ( .A(_820_), .B(_829_), .C(micro_abc_calculation_ints_imput_W2_logic_96_), .Y(_832_) );
AOI21X1 AOI21X1_90 ( .A(_832_), .B(_831_), .C(_822_), .Y(_816__96_) );
INVX1 INVX1_196 ( .A(micro_abc_calculation_ints_counter_2_), .Y(_833_) );
NAND3X1 NAND3X1_42 ( .A(micro_abc_calculation_ints_counter_3_), .B(_819_), .C(_833_), .Y(_834_) );
NOR2X1 NOR2X1_177 ( .A(_818_), .B(_834_), .Y(_835_) );
NAND2X1 NAND2X1_126 ( .A(nonce_2_1), .B(_835_), .Y(_836_) );
OAI21X1 OAI21X1_138 ( .A(_834_), .B(_818_), .C(micro_abc_calculation_ints_imput_W2_logic_88_), .Y(_837_) );
AOI21X1 AOI21X1_91 ( .A(_837_), .B(_836_), .C(_822_), .Y(_816__88_) );
NAND2X1 NAND2X1_127 ( .A(micro_abc_calculation_ints_counter_1_), .B(_828_), .Y(_838_) );
NOR2X1 NOR2X1_178 ( .A(_838_), .B(_834_), .Y(_839_) );
NAND2X1 NAND2X1_128 ( .A(nonce_2_0), .B(_839_), .Y(_840_) );
OAI21X1 OAI21X1_139 ( .A(_834_), .B(_838_), .C(micro_abc_calculation_ints_imput_W2_logic_80_), .Y(_841_) );
AOI21X1 AOI21X1_92 ( .A(_841_), .B(_840_), .C(_822_), .Y(_816__80_) );
NOR2X1 NOR2X1_179 ( .A(_824_), .B(_834_), .Y(_842_) );
NAND2X1 NAND2X1_129 ( .A(block11[0]), .B(_842_), .Y(_843_) );
OAI21X1 OAI21X1_140 ( .A(_834_), .B(_824_), .C(micro_abc_calculation_ints_imput_W2_logic_72_), .Y(_844_) );
AOI21X1 AOI21X1_93 ( .A(_844_), .B(_843_), .C(_822_), .Y(_816__72_) );
NOR2X1 NOR2X1_180 ( .A(_829_), .B(_834_), .Y(_845_) );
XOR2X1 XOR2X1_10 ( .A(block10[0]), .B(nonce_2_3), .Y(_846_) );
NAND2X1 NAND2X1_130 ( .A(_846_), .B(_845_), .Y(_847_) );
OAI21X1 OAI21X1_141 ( .A(_834_), .B(_829_), .C(micro_abc_calculation_ints_imput_W2_logic_64_), .Y(_848_) );
AOI21X1 AOI21X1_94 ( .A(_848_), .B(_847_), .C(_822_), .Y(_816__64_) );
INVX1 INVX1_197 ( .A(micro_abc_calculation_ints_counter_3_), .Y(_849_) );
NAND2X1 NAND2X1_131 ( .A(micro_abc_calculation_ints_counter_2_), .B(_849_), .Y(_850_) );
NAND3X1 NAND3X1_43 ( .A(micro_abc_calculation_ints_counter_1_), .B(micro_abc_calculation_ints_counter_0_), .C(_819_), .Y(_851_) );
NOR2X1 NOR2X1_181 ( .A(_850_), .B(_851_), .Y(_852_) );
XOR2X1 XOR2X1_11 ( .A(nonce_2_2), .B(block9[0]), .Y(_853_) );
NAND2X1 NAND2X1_132 ( .A(_853_), .B(_852_), .Y(_854_) );
OAI21X1 OAI21X1_142 ( .A(_851_), .B(_850_), .C(micro_abc_calculation_ints_imput_W2_logic_56_), .Y(_855_) );
AOI21X1 AOI21X1_95 ( .A(_855_), .B(_854_), .C(_822_), .Y(_816__56_) );
NAND3X1 NAND3X1_44 ( .A(micro_abc_calculation_ints_counter_1_), .B(_819_), .C(_828_), .Y(_856_) );
NOR2X1 NOR2X1_182 ( .A(_850_), .B(_856_), .Y(_857_) );
XOR2X1 XOR2X1_12 ( .A(nonce_2_1), .B(block8[0]), .Y(_858_) );
NAND2X1 NAND2X1_133 ( .A(_858_), .B(_857_), .Y(_859_) );
OAI21X1 OAI21X1_143 ( .A(_856_), .B(_850_), .C(micro_abc_calculation_ints_imput_W2_logic_48_), .Y(_860_) );
AOI21X1 AOI21X1_96 ( .A(_860_), .B(_859_), .C(_822_), .Y(_816__48_) );
NAND3X1 NAND3X1_45 ( .A(micro_abc_calculation_ints_counter_0_), .B(_819_), .C(_823_), .Y(_861_) );
NOR2X1 NOR2X1_183 ( .A(_850_), .B(_861_), .Y(_862_) );
XOR2X1 XOR2X1_13 ( .A(nonce_2_0), .B(block7[0]), .Y(_863_) );
NAND2X1 NAND2X1_134 ( .A(_863_), .B(_862_), .Y(_864_) );
OAI21X1 OAI21X1_144 ( .A(_861_), .B(_850_), .C(micro_abc_calculation_ints_imput_W2_logic_40_), .Y(_865_) );
AOI21X1 AOI21X1_97 ( .A(_865_), .B(_864_), .C(_822_), .Y(_816__40_) );
INVX1 INVX1_198 ( .A(_850_), .Y(_866_) );
NOR2X1 NOR2X1_184 ( .A(micro_abc_calculation_ints_counter_1_), .B(micro_abc_calculation_ints_counter_0_), .Y(_867_) );
NAND2X1 NAND2X1_135 ( .A(_819_), .B(_867_), .Y(_868_) );
INVX1 INVX1_199 ( .A(_868_), .Y(_869_) );
XOR2X1 XOR2X1_14 ( .A(block11[0]), .B(block6[0]), .Y(_870_) );
NAND3X1 NAND3X1_46 ( .A(_866_), .B(_870_), .C(_869_), .Y(_871_) );
OAI21X1 OAI21X1_145 ( .A(_868_), .B(_850_), .C(micro_abc_calculation_ints_imput_W2_logic_32_), .Y(_872_) );
AOI21X1 AOI21X1_98 ( .A(_872_), .B(_871_), .C(_822_), .Y(_816__32_) );
NOR2X1 NOR2X1_185 ( .A(micro_abc_calculation_ints_counter_3_), .B(micro_abc_calculation_ints_counter_2_), .Y(_873_) );
INVX4 INVX4_3 ( .A(_873_), .Y(_874_) );
NOR2X1 NOR2X1_186 ( .A(_874_), .B(_851_), .Y(_875_) );
XOR2X1 XOR2X1_15 ( .A(block10[0]), .B(block5[0]), .Y(_876_) );
NAND2X1 NAND2X1_136 ( .A(_876_), .B(_875_), .Y(_877_) );
OAI21X1 OAI21X1_146 ( .A(_851_), .B(_874_), .C(micro_abc_calculation_ints_imput_W2_logic_24_), .Y(_878_) );
AOI21X1 AOI21X1_99 ( .A(_878_), .B(_877_), .C(_822_), .Y(_816__24_) );
NOR2X1 NOR2X1_187 ( .A(_874_), .B(_856_), .Y(_879_) );
NOR2X1 NOR2X1_188 ( .A(nonce_2_3), .B(block9[0]), .Y(_880_) );
XOR2X1 XOR2X1_16 ( .A(_880_), .B(block4[0]), .Y(_881_) );
INVX1 INVX1_200 ( .A(micro_abc_calculation_ints_imput_W2_logic_16_), .Y(_882_) );
OAI21X1 OAI21X1_147 ( .A(_856_), .B(_874_), .C(_882_), .Y(_883_) );
NAND2X1 NAND2X1_137 ( .A(reset_bF_buf0), .B(_883_), .Y(_884_) );
AOI21X1 AOI21X1_100 ( .A(_879_), .B(_881_), .C(_884_), .Y(_816__16_) );
NOR2X1 NOR2X1_189 ( .A(_874_), .B(_861_), .Y(_885_) );
NOR2X1 NOR2X1_190 ( .A(nonce_2_2), .B(block8[0]), .Y(_886_) );
XOR2X1 XOR2X1_17 ( .A(_886_), .B(block3[0]), .Y(_887_) );
INVX1 INVX1_201 ( .A(micro_abc_calculation_ints_imput_W2_logic_8_), .Y(_888_) );
OAI21X1 OAI21X1_148 ( .A(_861_), .B(_874_), .C(_888_), .Y(_889_) );
NAND2X1 NAND2X1_138 ( .A(reset_bF_buf5), .B(_889_), .Y(_890_) );
AOI21X1 AOI21X1_101 ( .A(_885_), .B(_887_), .C(_890_), .Y(_816__8_) );
INVX1 INVX1_202 ( .A(micro_abc_calculation_ints_imput_W2_logic_0_), .Y(_891_) );
NAND3X1 NAND3X1_47 ( .A(_819_), .B(_867_), .C(_873_), .Y(_892_) );
AND2X2 AND2X2_31 ( .A(_892_), .B(_891_), .Y(_893_) );
OAI21X1 OAI21X1_149 ( .A(nonce_2_1), .B(block7[0]), .C(block2[0]), .Y(_894_) );
INVX1 INVX1_203 ( .A(block2[0]), .Y(_895_) );
NOR2X1 NOR2X1_191 ( .A(nonce_2_1), .B(block7[0]), .Y(_896_) );
NAND2X1 NAND2X1_139 ( .A(_895_), .B(_896_), .Y(_897_) );
AOI21X1 AOI21X1_102 ( .A(_894_), .B(_897_), .C(_892_), .Y(_898_) );
NOR3X1 NOR3X1_6 ( .A(_898_), .B(_822_), .C(_893_), .Y(_816__0_) );
NOR2X1 NOR2X1_192 ( .A(_838_), .B(_820_), .Y(_899_) );
NAND2X1 NAND2X1_140 ( .A(nonce_2_3), .B(_899_), .Y(_900_) );
OAI21X1 OAI21X1_150 ( .A(_820_), .B(_838_), .C(micro_abc_calculation_ints_imput_W2_logic_112_), .Y(_901_) );
AOI21X1 AOI21X1_103 ( .A(_901_), .B(_900_), .C(_822_), .Y(_816__112_) );
DFFPOSX1 DFFPOSX1_122 ( .CLK(clk_bF_buf10), .D(_816__0_), .Q(micro_abc_calculation_ints_imput_W2_logic_0_) );
DFFPOSX1 DFFPOSX1_123 ( .CLK(clk_bF_buf9), .D(_816__8_), .Q(micro_abc_calculation_ints_imput_W2_logic_8_) );
DFFPOSX1 DFFPOSX1_124 ( .CLK(clk_bF_buf8), .D(_816__16_), .Q(micro_abc_calculation_ints_imput_W2_logic_16_) );
DFFPOSX1 DFFPOSX1_125 ( .CLK(clk_bF_buf7), .D(_816__24_), .Q(micro_abc_calculation_ints_imput_W2_logic_24_) );
DFFPOSX1 DFFPOSX1_126 ( .CLK(clk_bF_buf6), .D(_816__32_), .Q(micro_abc_calculation_ints_imput_W2_logic_32_) );
DFFPOSX1 DFFPOSX1_127 ( .CLK(clk_bF_buf5), .D(_816__40_), .Q(micro_abc_calculation_ints_imput_W2_logic_40_) );
DFFPOSX1 DFFPOSX1_128 ( .CLK(clk_bF_buf4), .D(_816__48_), .Q(micro_abc_calculation_ints_imput_W2_logic_48_) );
DFFPOSX1 DFFPOSX1_129 ( .CLK(clk_bF_buf3), .D(_816__56_), .Q(micro_abc_calculation_ints_imput_W2_logic_56_) );
DFFPOSX1 DFFPOSX1_130 ( .CLK(clk_bF_buf2), .D(_816__64_), .Q(micro_abc_calculation_ints_imput_W2_logic_64_) );
DFFPOSX1 DFFPOSX1_131 ( .CLK(clk_bF_buf1), .D(_816__72_), .Q(micro_abc_calculation_ints_imput_W2_logic_72_) );
DFFPOSX1 DFFPOSX1_132 ( .CLK(clk_bF_buf0), .D(_816__80_), .Q(micro_abc_calculation_ints_imput_W2_logic_80_) );
DFFPOSX1 DFFPOSX1_133 ( .CLK(clk_bF_buf11), .D(_816__88_), .Q(micro_abc_calculation_ints_imput_W2_logic_88_) );
DFFPOSX1 DFFPOSX1_134 ( .CLK(clk_bF_buf10), .D(_816__96_), .Q(micro_abc_calculation_ints_imput_W2_logic_96_) );
DFFPOSX1 DFFPOSX1_135 ( .CLK(clk_bF_buf9), .D(_816__104_), .Q(micro_abc_calculation_ints_imput_W2_logic_104_) );
DFFPOSX1 DFFPOSX1_136 ( .CLK(clk_bF_buf8), .D(_816__112_), .Q(micro_abc_calculation_ints_imput_W2_logic_112_) );
DFFPOSX1 DFFPOSX1_137 ( .CLK(clk_bF_buf7), .D(_816__120_), .Q(micro_abc_calculation_ints_imput_W2_logic_120_) );
INVX2 INVX2_16 ( .A(gnd), .Y(_911_) );
INVX1 INVX1_204 ( .A(nonce_nonce_int_3_0_), .Y(_912_) );
INVX1 INVX1_205 ( .A(reset_bF_buf4), .Y(_913_) );
NOR2X1 NOR2X1_193 ( .A(fail), .B(_913_), .Y(_914_) );
INVX2 INVX2_17 ( .A(_914_), .Y(_915_) );
NOR2X1 NOR2X1_194 ( .A(nonce_delay), .B(_915_), .Y(_916_) );
INVX1 INVX1_206 ( .A(_916_), .Y(_917_) );
INVX4 INVX4_4 ( .A(gnd), .Y(_918_) );
NOR2X1 NOR2X1_195 ( .A(gnd), .B(_918_), .Y(_919_) );
INVX1 INVX1_207 ( .A(_919_), .Y(_920_) );
NOR2X1 NOR2X1_196 ( .A(_920_), .B(_917_), .Y(_921_) );
MUX2X1 MUX2X1_5 ( .A(_911_), .B(_912_), .S(_921_), .Y(_910__0_) );
INVX2 INVX2_18 ( .A(nonce_nonce_int_2_0_), .Y(_922_) );
INVX2 INVX2_19 ( .A(gnd), .Y(_923_) );
NOR2X1 NOR2X1_197 ( .A(gnd), .B(_923_), .Y(_924_) );
NAND2X1 NAND2X1_141 ( .A(_924_), .B(_916_), .Y(_925_) );
MUX2X1 MUX2X1_6 ( .A(_922_), .B(_911_), .S(_925_), .Y(_909__0_) );
INVX2 INVX2_20 ( .A(nonce_nonce_int_1_0_), .Y(_926_) );
NAND2X1 NAND2X1_142 ( .A(_923_), .B(_914_), .Y(_927_) );
NOR2X1 NOR2X1_198 ( .A(nonce_delay), .B(_927_), .Y(_928_) );
MUX2X1 MUX2X1_7 ( .A(_911_), .B(_926_), .S(_928_), .Y(_908__0_) );
INVX4 INVX4_5 ( .A(nonce_delay), .Y(_929_) );
NOR2X1 NOR2X1_199 ( .A(gnd), .B(_929_), .Y(_930_) );
INVX1 INVX1_208 ( .A(_930_), .Y(_931_) );
NOR2X1 NOR2X1_200 ( .A(gnd), .B(nonce_nonce_int_0_0_), .Y(_932_) );
NAND2X1 NAND2X1_143 ( .A(gnd), .B(nonce_nonce_int_0_0_), .Y(_933_) );
INVX1 INVX1_209 ( .A(_933_), .Y(_934_) );
NOR2X1 NOR2X1_201 ( .A(_932_), .B(_934_), .Y(_935_) );
NAND2X1 NAND2X1_144 ( .A(nonce_delay), .B(_924_), .Y(_936_) );
INVX1 INVX1_210 ( .A(_936_), .Y(_937_) );
OAI21X1 OAI21X1_151 ( .A(_923_), .B(_918_), .C(nonce_delay), .Y(_938_) );
AOI22X1 AOI22X1_23 ( .A(nonce_2_1), .B(_938_), .C(_937_), .D(_935_), .Y(_939_) );
OAI21X1 OAI21X1_152 ( .A(_926_), .B(_931_), .C(_939_), .Y(_940_) );
AND2X2 AND2X2_32 ( .A(_940_), .B(_914_), .Y(_904__0_) );
NAND2X1 NAND2X1_145 ( .A(nonce_delay), .B(_919_), .Y(_941_) );
NOR2X1 NOR2X1_202 ( .A(gnd), .B(gnd), .Y(_942_) );
INVX1 INVX1_211 ( .A(_942_), .Y(_943_) );
OAI21X1 OAI21X1_153 ( .A(_929_), .B(gnd), .C(gnd), .Y(_944_) );
INVX1 INVX1_212 ( .A(nonce_nonce_int_0_0_), .Y(_945_) );
OAI21X1 OAI21X1_154 ( .A(_929_), .B(_945_), .C(_918_), .Y(_946_) );
AOI21X1 AOI21X1_104 ( .A(_944_), .B(_946_), .C(nonce_2_0), .Y(_947_) );
INVX1 INVX1_213 ( .A(_941_), .Y(_948_) );
INVX2 INVX2_21 ( .A(gnd), .Y(_949_) );
NAND2X1 NAND2X1_146 ( .A(_926_), .B(_949_), .Y(_950_) );
NAND2X1 NAND2X1_147 ( .A(nonce_nonce_int_1_0_), .B(gnd), .Y(_951_) );
AND2X2 AND2X2_33 ( .A(_950_), .B(_951_), .Y(_952_) );
INVX1 INVX1_214 ( .A(_952_), .Y(_953_) );
AOI21X1 AOI21X1_105 ( .A(_948_), .B(_953_), .C(_915_), .Y(_954_) );
OAI21X1 OAI21X1_155 ( .A(_929_), .B(_946_), .C(_954_), .Y(_955_) );
NOR2X1 NOR2X1_203 ( .A(_947_), .B(_955_), .Y(_903__0_) );
NOR2X1 NOR2X1_204 ( .A(gnd), .B(_929_), .Y(_956_) );
INVX1 INVX1_215 ( .A(_946_), .Y(_957_) );
AOI21X1 AOI21X1_106 ( .A(_918_), .B(_914_), .C(nonce_nonce_int_0_0_), .Y(_958_) );
AOI21X1 AOI21X1_107 ( .A(gnd), .B(_929_), .C(_915_), .Y(_959_) );
AOI21X1 AOI21X1_108 ( .A(_957_), .B(_959_), .C(_958_), .Y(_907__0_) );
AND2X2 AND2X2_34 ( .A(_929_), .B(nonce_2_3), .Y(_960_) );
OAI21X1 OAI21X1_156 ( .A(_922_), .B(_949_), .C(nonce_delay), .Y(_961_) );
AOI21X1 AOI21X1_109 ( .A(_922_), .B(_949_), .C(_961_), .Y(_962_) );
OAI21X1 OAI21X1_157 ( .A(_962_), .B(_960_), .C(_924_), .Y(_963_) );
OAI21X1 OAI21X1_158 ( .A(_943_), .B(nonce_delay), .C(_944_), .Y(_964_) );
NAND2X1 NAND2X1_148 ( .A(_918_), .B(_930_), .Y(_965_) );
OAI22X1 OAI22X1_9 ( .A(_941_), .B(_912_), .C(_953_), .D(_965_), .Y(_966_) );
AOI21X1 AOI21X1_110 ( .A(nonce_2_3), .B(_964_), .C(_966_), .Y(_967_) );
AOI21X1 AOI21X1_111 ( .A(_963_), .B(_967_), .C(_915_), .Y(_906__0_) );
NOR2X1 NOR2X1_205 ( .A(nonce_nonce_int_3_0_), .B(gnd), .Y(_968_) );
AND2X2 AND2X2_35 ( .A(nonce_nonce_int_3_0_), .B(gnd), .Y(_969_) );
OAI21X1 OAI21X1_159 ( .A(_969_), .B(_968_), .C(gnd), .Y(_970_) );
OAI21X1 OAI21X1_160 ( .A(_935_), .B(gnd), .C(_970_), .Y(_971_) );
NAND2X1 NAND2X1_149 ( .A(_930_), .B(_971_), .Y(_972_) );
NAND2X1 NAND2X1_150 ( .A(_922_), .B(_956_), .Y(_973_) );
OAI21X1 OAI21X1_161 ( .A(_918_), .B(nonce_2_2), .C(_973_), .Y(_974_) );
OAI21X1 OAI21X1_162 ( .A(nonce_delay), .B(nonce_2_2), .C(_914_), .Y(_975_) );
AOI21X1 AOI21X1_112 ( .A(gnd), .B(_974_), .C(_975_), .Y(_976_) );
AND2X2 AND2X2_36 ( .A(_976_), .B(_972_), .Y(_905__0_) );
OAI21X1 OAI21X1_163 ( .A(_923_), .B(_918_), .C(_914_), .Y(_977_) );
XNOR2X1 XNOR2X1_26 ( .A(_977_), .B(nonce_delay), .Y(_902_) );
DFFPOSX1 DFFPOSX1_138 ( .CLK(clk_bF_buf6), .D(_902_), .Q(nonce_delay) );
DFFPOSX1 DFFPOSX1_139 ( .CLK(clk_bF_buf5), .D(_905__0_), .Q(nonce_2_2) );
DFFPOSX1 DFFPOSX1_140 ( .CLK(clk_bF_buf4), .D(_906__0_), .Q(nonce_2_3) );
DFFPOSX1 DFFPOSX1_141 ( .CLK(clk_bF_buf3), .D(_907__0_), .Q(nonce_nonce_int_0_0_) );
DFFPOSX1 DFFPOSX1_142 ( .CLK(clk_bF_buf2), .D(_903__0_), .Q(nonce_2_0) );
DFFPOSX1 DFFPOSX1_143 ( .CLK(clk_bF_buf1), .D(_904__0_), .Q(nonce_2_1) );
DFFPOSX1 DFFPOSX1_144 ( .CLK(clk_bF_buf0), .D(_908__0_), .Q(nonce_nonce_int_1_0_) );
DFFPOSX1 DFFPOSX1_145 ( .CLK(clk_bF_buf11), .D(_909__0_), .Q(nonce_nonce_int_2_0_) );
DFFPOSX1 DFFPOSX1_146 ( .CLK(clk_bF_buf10), .D(_910__0_), .Q(nonce_nonce_int_3_0_) );
INVX1 INVX1_216 ( .A(compare_hash_0_compare_var_0_), .Y(_987_) );
AND2X2 AND2X2_37 ( .A(compare_hash_1_compare_var_2_), .B(compare_hash_0_compare_var_2_), .Y(_979_) );
NOR2X1 NOR2X1_206 ( .A(compare_hash_1_compare_var_2_), .B(compare_hash_0_compare_var_2_), .Y(_980_) );
OAI22X1 OAI22X1_10 ( .A(compare_hash_1_compare_var_0_), .B(_987_), .C(_979_), .D(_980_), .Y(_981_) );
INVX1 INVX1_217 ( .A(compare_hash_1_compare_var_0_), .Y(_982_) );
INVX1 INVX1_218 ( .A(compare_hash_1_compare_var_1_), .Y(_983_) );
OAI22X1 OAI22X1_11 ( .A(_982_), .B(compare_hash_0_compare_var_0_), .C(_983_), .D(compare_hash_0_compare_var_1_), .Y(_984_) );
INVX1 INVX1_219 ( .A(compare_hash_0_compare_var_1_), .Y(_985_) );
OAI21X1 OAI21X1_164 ( .A(_985_), .B(compare_hash_1_compare_var_1_), .C(reset_bF_buf3), .Y(_986_) );
NOR3X1 NOR3X1_7 ( .A(_984_), .B(_986_), .C(_981_), .Y(_978_) );
DFFPOSX1 DFFPOSX1_147 ( .CLK(clk_bF_buf9), .D(_978_), .Q(validity_validity_reg) );
INVX8 INVX8_4 ( .A(reset_bF_buf2), .Y(_10_) );
INVX1 INVX1_220 ( .A(counter_1_), .Y(_11_) );
NAND3X1 NAND3X1_48 ( .A(counter_0_), .B(invalid_nonce), .C(_11_), .Y(_12_) );
NOR2X1 NOR2X1_207 ( .A(counter_5_), .B(counter_4_), .Y(_13_) );
NOR2X1 NOR2X1_208 ( .A(counter_7_), .B(counter_6_), .Y(_14_) );
NAND2X1 NAND2X1_151 ( .A(_13_), .B(_14_), .Y(_15_) );
INVX1 INVX1_221 ( .A(counter_2_), .Y(_16_) );
NAND2X1 NAND2X1_152 ( .A(counter_3_), .B(_16_), .Y(_17_) );
NOR3X1 NOR3X1_8 ( .A(_12_), .B(_17_), .C(_15_), .Y(_18_) );
INVX1 INVX1_222 ( .A(start), .Y(_19_) );
NOR2X1 NOR2X1_209 ( .A(_135_), .B(_19_), .Y(_20_) );
NAND3X1 NAND3X1_49 ( .A(current_loop_actualize_0_), .B(_20__bF_buf2), .C(_18__bF_buf3), .Y(_21_) );
BUFX2 BUFX2_35 ( .A(gnd), .Y(_548__8_) );
BUFX2 BUFX2_36 ( .A(gnd), .Y(_548__9_) );
BUFX2 BUFX2_37 ( .A(gnd), .Y(_548__10_) );
BUFX2 BUFX2_38 ( .A(gnd), .Y(_548__11_) );
BUFX2 BUFX2_39 ( .A(gnd), .Y(_806__1_) );
BUFX2 BUFX2_40 ( .A(gnd), .Y(_806__2_) );
BUFX2 BUFX2_41 ( .A(gnd), .Y(_806__6_) );
endmodule
